library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"24",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"0a",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"24",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"e0",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"1a",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"24",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"0a",	--29
		x"f9",	--30
		x"31",	--31
		x"a6",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"42",	--44
		x"b0",	--45
		x"f4",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"f8",	--50
		x"b0",	--51
		x"06",	--52
		x"21",	--53
		x"3d",	--54
		x"15",	--55
		x"3e",	--56
		x"b4",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"24",	--61
		x"3d",	--62
		x"26",	--63
		x"3e",	--64
		x"24",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"24",	--69
		x"3d",	--70
		x"2c",	--71
		x"3e",	--72
		x"98",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"24",	--77
		x"3d",	--78
		x"31",	--79
		x"3e",	--80
		x"54",	--81
		x"7f",	--82
		x"70",	--83
		x"b0",	--84
		x"24",	--85
		x"3d",	--86
		x"35",	--87
		x"3e",	--88
		x"94",	--89
		x"7f",	--90
		x"65",	--91
		x"b0",	--92
		x"24",	--93
		x"3d",	--94
		x"3d",	--95
		x"3e",	--96
		x"dc",	--97
		x"7f",	--98
		x"73",	--99
		x"b0",	--100
		x"24",	--101
		x"3d",	--102
		x"4e",	--103
		x"3e",	--104
		x"e0",	--105
		x"7f",	--106
		x"63",	--107
		x"b0",	--108
		x"24",	--109
		x"3d",	--110
		x"62",	--111
		x"3e",	--112
		x"e4",	--113
		x"7f",	--114
		x"62",	--115
		x"b0",	--116
		x"24",	--117
		x"0e",	--118
		x"0f",	--119
		x"b0",	--120
		x"ba",	--121
		x"2c",	--122
		x"3d",	--123
		x"20",	--124
		x"3e",	--125
		x"80",	--126
		x"0f",	--127
		x"3f",	--128
		x"0e",	--129
		x"b0",	--130
		x"c2",	--131
		x"0f",	--132
		x"3f",	--133
		x"0e",	--134
		x"b0",	--135
		x"0a",	--136
		x"2c",	--137
		x"3d",	--138
		x"20",	--139
		x"3e",	--140
		x"88",	--141
		x"0f",	--142
		x"2f",	--143
		x"b0",	--144
		x"c2",	--145
		x"0f",	--146
		x"2f",	--147
		x"b0",	--148
		x"0a",	--149
		x"0e",	--150
		x"2e",	--151
		x"0f",	--152
		x"3f",	--153
		x"0e",	--154
		x"b0",	--155
		x"4a",	--156
		x"3e",	--157
		x"98",	--158
		x"0f",	--159
		x"2f",	--160
		x"b0",	--161
		x"18",	--162
		x"3e",	--163
		x"9c",	--164
		x"0f",	--165
		x"b0",	--166
		x"18",	--167
		x"0e",	--168
		x"0f",	--169
		x"2f",	--170
		x"b0",	--171
		x"80",	--172
		x"0e",	--173
		x"2e",	--174
		x"0f",	--175
		x"3f",	--176
		x"0e",	--177
		x"b0",	--178
		x"8a",	--179
		x"b0",	--180
		x"f0",	--181
		x"3e",	--182
		x"ff",	--183
		x"3f",	--184
		x"9e",	--185
		x"b0",	--186
		x"00",	--187
		x"0d",	--188
		x"3e",	--189
		x"e8",	--190
		x"b0",	--191
		x"44",	--192
		x"0c",	--193
		x"0d",	--194
		x"1e",	--195
		x"0f",	--196
		x"3f",	--197
		x"24",	--198
		x"b0",	--199
		x"12",	--200
		x"0c",	--201
		x"0d",	--202
		x"1e",	--203
		x"0f",	--204
		x"3f",	--205
		x"18",	--206
		x"b0",	--207
		x"12",	--208
		x"0e",	--209
		x"3e",	--210
		x"18",	--211
		x"0f",	--212
		x"3f",	--213
		x"24",	--214
		x"b0",	--215
		x"da",	--216
		x"f2",	--217
		x"80",	--218
		x"19",	--219
		x"32",	--220
		x"0b",	--221
		x"b0",	--222
		x"60",	--223
		x"0f",	--224
		x"fc",	--225
		x"b0",	--226
		x"88",	--227
		x"7f",	--228
		x"15",	--229
		x"7f",	--230
		x"0d",	--231
		x"1b",	--232
		x"30",	--233
		x"6d",	--234
		x"b0",	--235
		x"06",	--236
		x"21",	--237
		x"3f",	--238
		x"30",	--239
		x"0f",	--240
		x"0b",	--241
		x"cb",	--242
		x"00",	--243
		x"0e",	--244
		x"5f",	--245
		x"30",	--246
		x"b0",	--247
		x"58",	--248
		x"0b",	--249
		x"e3",	--250
		x"0b",	--251
		x"e1",	--252
		x"3b",	--253
		x"30",	--254
		x"70",	--255
		x"b0",	--256
		x"06",	--257
		x"21",	--258
		x"da",	--259
		x"3b",	--260
		x"28",	--261
		x"d7",	--262
		x"82",	--263
		x"0c",	--264
		x"0c",	--265
		x"4e",	--266
		x"8e",	--267
		x"0e",	--268
		x"30",	--269
		x"74",	--270
		x"81",	--271
		x"5c",	--272
		x"b0",	--273
		x"06",	--274
		x"21",	--275
		x"1f",	--276
		x"58",	--277
		x"3e",	--278
		x"30",	--279
		x"0e",	--280
		x"0e",	--281
		x"ce",	--282
		x"00",	--283
		x"1b",	--284
		x"c0",	--285
		x"30",	--286
		x"3e",	--287
		x"8f",	--288
		x"00",	--289
		x"8f",	--290
		x"02",	--291
		x"8f",	--292
		x"04",	--293
		x"8f",	--294
		x"06",	--295
		x"8f",	--296
		x"08",	--297
		x"8f",	--298
		x"0a",	--299
		x"30",	--300
		x"8f",	--301
		x"06",	--302
		x"8f",	--303
		x"08",	--304
		x"8f",	--305
		x"0a",	--306
		x"30",	--307
		x"8f",	--308
		x"00",	--309
		x"30",	--310
		x"8f",	--311
		x"02",	--312
		x"30",	--313
		x"8f",	--314
		x"04",	--315
		x"30",	--316
		x"8f",	--317
		x"06",	--318
		x"30",	--319
		x"1d",	--320
		x"06",	--321
		x"0d",	--322
		x"0e",	--323
		x"1d",	--324
		x"08",	--325
		x"8f",	--326
		x"08",	--327
		x"02",	--328
		x"32",	--329
		x"03",	--330
		x"82",	--331
		x"32",	--332
		x"a2",	--333
		x"38",	--334
		x"1c",	--335
		x"3a",	--336
		x"32",	--337
		x"02",	--338
		x"32",	--339
		x"03",	--340
		x"82",	--341
		x"32",	--342
		x"92",	--343
		x"02",	--344
		x"38",	--345
		x"1d",	--346
		x"3a",	--347
		x"32",	--348
		x"0d",	--349
		x"1e",	--350
		x"0a",	--351
		x"02",	--352
		x"32",	--353
		x"03",	--354
		x"82",	--355
		x"32",	--356
		x"92",	--357
		x"04",	--358
		x"38",	--359
		x"1f",	--360
		x"3a",	--361
		x"32",	--362
		x"0f",	--363
		x"30",	--364
		x"30",	--365
		x"0f",	--366
		x"30",	--367
		x"0f",	--368
		x"30",	--369
		x"b2",	--370
		x"00",	--371
		x"92",	--372
		x"b2",	--373
		x"30",	--374
		x"94",	--375
		x"b2",	--376
		x"41",	--377
		x"96",	--378
		x"30",	--379
		x"46",	--380
		x"b0",	--381
		x"06",	--382
		x"92",	--383
		x"90",	--384
		x"b1",	--385
		x"64",	--386
		x"00",	--387
		x"b0",	--388
		x"06",	--389
		x"21",	--390
		x"0f",	--391
		x"30",	--392
		x"b0",	--393
		x"40",	--394
		x"30",	--395
		x"0b",	--396
		x"0a",	--397
		x"0a",	--398
		x"3b",	--399
		x"00",	--400
		x"0d",	--401
		x"0e",	--402
		x"1f",	--403
		x"1e",	--404
		x"b0",	--405
		x"5e",	--406
		x"0d",	--407
		x"0e",	--408
		x"1f",	--409
		x"1c",	--410
		x"b0",	--411
		x"5e",	--412
		x"30",	--413
		x"7d",	--414
		x"b0",	--415
		x"06",	--416
		x"21",	--417
		x"3a",	--418
		x"3b",	--419
		x"30",	--420
		x"82",	--421
		x"1e",	--422
		x"82",	--423
		x"1c",	--424
		x"30",	--425
		x"0b",	--426
		x"0a",	--427
		x"21",	--428
		x"0a",	--429
		x"0b",	--430
		x"b2",	--431
		x"00",	--432
		x"4e",	--433
		x"3a",	--434
		x"03",	--435
		x"53",	--436
		x"3e",	--437
		x"0e",	--438
		x"1f",	--439
		x"02",	--440
		x"b0",	--441
		x"f4",	--442
		x"0a",	--443
		x"0e",	--444
		x"1f",	--445
		x"04",	--446
		x"b0",	--447
		x"f4",	--448
		x"0b",	--449
		x"0f",	--450
		x"0a",	--451
		x"30",	--452
		x"ca",	--453
		x"b0",	--454
		x"06",	--455
		x"31",	--456
		x"06",	--457
		x"0e",	--458
		x"0f",	--459
		x"b0",	--460
		x"7a",	--461
		x"0c",	--462
		x"3d",	--463
		x"c8",	--464
		x"b0",	--465
		x"4a",	--466
		x"0c",	--467
		x"0d",	--468
		x"0e",	--469
		x"3f",	--470
		x"80",	--471
		x"b0",	--472
		x"d6",	--473
		x"0d",	--474
		x"0e",	--475
		x"1f",	--476
		x"1e",	--477
		x"b0",	--478
		x"5e",	--479
		x"0e",	--480
		x"0f",	--481
		x"b0",	--482
		x"7a",	--483
		x"0c",	--484
		x"3d",	--485
		x"c8",	--486
		x"b0",	--487
		x"4a",	--488
		x"0d",	--489
		x"0e",	--490
		x"1f",	--491
		x"1c",	--492
		x"b0",	--493
		x"5e",	--494
		x"0f",	--495
		x"21",	--496
		x"3a",	--497
		x"3b",	--498
		x"30",	--499
		x"0e",	--500
		x"1f",	--501
		x"06",	--502
		x"b0",	--503
		x"f4",	--504
		x"1d",	--505
		x"0e",	--506
		x"1f",	--507
		x"00",	--508
		x"b0",	--509
		x"44",	--510
		x"b6",	--511
		x"0e",	--512
		x"3f",	--513
		x"18",	--514
		x"b0",	--515
		x"00",	--516
		x"82",	--517
		x"00",	--518
		x"aa",	--519
		x"30",	--520
		x"84",	--521
		x"b0",	--522
		x"06",	--523
		x"b1",	--524
		x"9e",	--525
		x"00",	--526
		x"b0",	--527
		x"06",	--528
		x"a1",	--529
		x"00",	--530
		x"30",	--531
		x"af",	--532
		x"b0",	--533
		x"06",	--534
		x"21",	--535
		x"3f",	--536
		x"d6",	--537
		x"0b",	--538
		x"0a",	--539
		x"1f",	--540
		x"22",	--541
		x"b0",	--542
		x"20",	--543
		x"0a",	--544
		x"0b",	--545
		x"1f",	--546
		x"20",	--547
		x"b0",	--548
		x"20",	--549
		x"0b",	--550
		x"0a",	--551
		x"3e",	--552
		x"3f",	--553
		x"1e",	--554
		x"0f",	--555
		x"0f",	--556
		x"0e",	--557
		x"30",	--558
		x"d2",	--559
		x"30",	--560
		x"24",	--561
		x"b0",	--562
		x"d2",	--563
		x"31",	--564
		x"0c",	--565
		x"30",	--566
		x"24",	--567
		x"30",	--568
		x"da",	--569
		x"b0",	--570
		x"06",	--571
		x"21",	--572
		x"3a",	--573
		x"3b",	--574
		x"30",	--575
		x"82",	--576
		x"20",	--577
		x"82",	--578
		x"22",	--579
		x"30",	--580
		x"82",	--581
		x"1e",	--582
		x"82",	--583
		x"1c",	--584
		x"30",	--585
		x"0b",	--586
		x"0a",	--587
		x"09",	--588
		x"08",	--589
		x"21",	--590
		x"0a",	--591
		x"0b",	--592
		x"81",	--593
		x"00",	--594
		x"1f",	--595
		x"1c",	--596
		x"b2",	--597
		x"02",	--598
		x"6f",	--599
		x"92",	--600
		x"0a",	--601
		x"0e",	--602
		x"1f",	--603
		x"02",	--604
		x"b0",	--605
		x"f4",	--606
		x"08",	--607
		x"3a",	--608
		x"03",	--609
		x"1e",	--610
		x"09",	--611
		x"0d",	--612
		x"0e",	--613
		x"1f",	--614
		x"02",	--615
		x"b0",	--616
		x"44",	--617
		x"0f",	--618
		x"21",	--619
		x"38",	--620
		x"39",	--621
		x"3a",	--622
		x"3b",	--623
		x"30",	--624
		x"82",	--625
		x"0a",	--626
		x"49",	--627
		x"82",	--628
		x"0a",	--629
		x"1f",	--630
		x"02",	--631
		x"b0",	--632
		x"6c",	--633
		x"0f",	--634
		x"21",	--635
		x"38",	--636
		x"39",	--637
		x"3a",	--638
		x"3b",	--639
		x"30",	--640
		x"0e",	--641
		x"1f",	--642
		x"04",	--643
		x"b0",	--644
		x"f4",	--645
		x"09",	--646
		x"3a",	--647
		x"05",	--648
		x"da",	--649
		x"0e",	--650
		x"1f",	--651
		x"06",	--652
		x"b0",	--653
		x"f4",	--654
		x"0a",	--655
		x"0e",	--656
		x"1f",	--657
		x"08",	--658
		x"b0",	--659
		x"f4",	--660
		x"0b",	--661
		x"0f",	--662
		x"0a",	--663
		x"30",	--664
		x"df",	--665
		x"b0",	--666
		x"06",	--667
		x"31",	--668
		x"06",	--669
		x"0e",	--670
		x"0f",	--671
		x"b0",	--672
		x"7a",	--673
		x"0c",	--674
		x"3d",	--675
		x"c8",	--676
		x"b0",	--677
		x"4a",	--678
		x"0d",	--679
		x"0e",	--680
		x"1f",	--681
		x"1e",	--682
		x"b0",	--683
		x"5e",	--684
		x"0e",	--685
		x"0f",	--686
		x"b0",	--687
		x"7a",	--688
		x"0c",	--689
		x"3d",	--690
		x"c8",	--691
		x"b0",	--692
		x"4a",	--693
		x"0d",	--694
		x"0e",	--695
		x"1f",	--696
		x"1c",	--697
		x"b0",	--698
		x"5e",	--699
		x"a7",	--700
		x"0f",	--701
		x"b0",	--702
		x"34",	--703
		x"0f",	--704
		x"21",	--705
		x"38",	--706
		x"39",	--707
		x"3a",	--708
		x"3b",	--709
		x"30",	--710
		x"0e",	--711
		x"3f",	--712
		x"34",	--713
		x"b0",	--714
		x"00",	--715
		x"82",	--716
		x"02",	--717
		x"89",	--718
		x"5e",	--719
		x"19",	--720
		x"4e",	--721
		x"0f",	--722
		x"03",	--723
		x"c2",	--724
		x"19",	--725
		x"30",	--726
		x"c2",	--727
		x"19",	--728
		x"30",	--729
		x"1f",	--730
		x"82",	--731
		x"0c",	--732
		x"01",	--733
		x"0f",	--734
		x"82",	--735
		x"0c",	--736
		x"0f",	--737
		x"30",	--738
		x"1e",	--739
		x"0e",	--740
		x"3e",	--741
		x"06",	--742
		x"0f",	--743
		x"0f",	--744
		x"10",	--745
		x"e8",	--746
		x"c2",	--747
		x"19",	--748
		x"3e",	--749
		x"07",	--750
		x"03",	--751
		x"82",	--752
		x"0e",	--753
		x"30",	--754
		x"1e",	--755
		x"82",	--756
		x"0e",	--757
		x"30",	--758
		x"f2",	--759
		x"0e",	--760
		x"19",	--761
		x"f2",	--762
		x"f2",	--763
		x"0a",	--764
		x"19",	--765
		x"ee",	--766
		x"e2",	--767
		x"19",	--768
		x"eb",	--769
		x"f2",	--770
		x"0d",	--771
		x"19",	--772
		x"e7",	--773
		x"f2",	--774
		x"09",	--775
		x"19",	--776
		x"e3",	--777
		x"f2",	--778
		x"03",	--779
		x"19",	--780
		x"df",	--781
		x"f2",	--782
		x"07",	--783
		x"19",	--784
		x"db",	--785
		x"0b",	--786
		x"0a",	--787
		x"21",	--788
		x"0a",	--789
		x"0b",	--790
		x"30",	--791
		x"78",	--792
		x"b0",	--793
		x"06",	--794
		x"21",	--795
		x"3a",	--796
		x"03",	--797
		x"1b",	--798
		x"0e",	--799
		x"1f",	--800
		x"02",	--801
		x"b0",	--802
		x"f4",	--803
		x"0a",	--804
		x"0e",	--805
		x"1f",	--806
		x"04",	--807
		x"b0",	--808
		x"f4",	--809
		x"0b",	--810
		x"0f",	--811
		x"0a",	--812
		x"30",	--813
		x"c0",	--814
		x"b0",	--815
		x"06",	--816
		x"31",	--817
		x"06",	--818
		x"8a",	--819
		x"00",	--820
		x"0f",	--821
		x"21",	--822
		x"3a",	--823
		x"3b",	--824
		x"30",	--825
		x"30",	--826
		x"80",	--827
		x"b0",	--828
		x"06",	--829
		x"b1",	--830
		x"9a",	--831
		x"00",	--832
		x"b0",	--833
		x"06",	--834
		x"a1",	--835
		x"00",	--836
		x"30",	--837
		x"ab",	--838
		x"b0",	--839
		x"06",	--840
		x"21",	--841
		x"3f",	--842
		x"ea",	--843
		x"0b",	--844
		x"21",	--845
		x"0b",	--846
		x"1f",	--847
		x"17",	--848
		x"16",	--849
		x"30",	--850
		x"db",	--851
		x"b0",	--852
		x"06",	--853
		x"21",	--854
		x"0e",	--855
		x"1f",	--856
		x"02",	--857
		x"b0",	--858
		x"f4",	--859
		x"2f",	--860
		x"0f",	--861
		x"30",	--862
		x"c0",	--863
		x"b0",	--864
		x"06",	--865
		x"31",	--866
		x"06",	--867
		x"0f",	--868
		x"21",	--869
		x"3b",	--870
		x"30",	--871
		x"30",	--872
		x"80",	--873
		x"b0",	--874
		x"06",	--875
		x"b1",	--876
		x"9a",	--877
		x"00",	--878
		x"b0",	--879
		x"06",	--880
		x"a1",	--881
		x"00",	--882
		x"30",	--883
		x"cc",	--884
		x"b0",	--885
		x"06",	--886
		x"21",	--887
		x"3f",	--888
		x"eb",	--889
		x"0b",	--890
		x"0a",	--891
		x"8e",	--892
		x"00",	--893
		x"6d",	--894
		x"4d",	--895
		x"5e",	--896
		x"1f",	--897
		x"0a",	--898
		x"0c",	--899
		x"0f",	--900
		x"7b",	--901
		x"0a",	--902
		x"2b",	--903
		x"0c",	--904
		x"0c",	--905
		x"0c",	--906
		x"0c",	--907
		x"8d",	--908
		x"0c",	--909
		x"3c",	--910
		x"d0",	--911
		x"1a",	--912
		x"7d",	--913
		x"4d",	--914
		x"17",	--915
		x"7d",	--916
		x"78",	--917
		x"1a",	--918
		x"4b",	--919
		x"7b",	--920
		x"d0",	--921
		x"0a",	--922
		x"e9",	--923
		x"7b",	--924
		x"0a",	--925
		x"34",	--926
		x"0c",	--927
		x"0b",	--928
		x"0b",	--929
		x"0b",	--930
		x"0c",	--931
		x"8d",	--932
		x"0c",	--933
		x"3c",	--934
		x"d0",	--935
		x"7d",	--936
		x"4d",	--937
		x"e9",	--938
		x"9e",	--939
		x"00",	--940
		x"0f",	--941
		x"3a",	--942
		x"3b",	--943
		x"30",	--944
		x"1a",	--945
		x"de",	--946
		x"4b",	--947
		x"7b",	--948
		x"9f",	--949
		x"7b",	--950
		x"06",	--951
		x"0a",	--952
		x"0c",	--953
		x"0c",	--954
		x"0c",	--955
		x"0c",	--956
		x"8d",	--957
		x"0c",	--958
		x"3c",	--959
		x"a9",	--960
		x"1a",	--961
		x"ce",	--962
		x"4b",	--963
		x"7b",	--964
		x"bf",	--965
		x"7b",	--966
		x"06",	--967
		x"0a",	--968
		x"0c",	--969
		x"0c",	--970
		x"0c",	--971
		x"0c",	--972
		x"8d",	--973
		x"0c",	--974
		x"3c",	--975
		x"c9",	--976
		x"1a",	--977
		x"be",	--978
		x"8d",	--979
		x"0d",	--980
		x"30",	--981
		x"e2",	--982
		x"b0",	--983
		x"06",	--984
		x"21",	--985
		x"0c",	--986
		x"0f",	--987
		x"3a",	--988
		x"3b",	--989
		x"30",	--990
		x"0c",	--991
		x"ca",	--992
		x"0b",	--993
		x"0a",	--994
		x"0b",	--995
		x"0a",	--996
		x"8f",	--997
		x"00",	--998
		x"8f",	--999
		x"02",	--1000
		x"8f",	--1001
		x"04",	--1002
		x"0c",	--1003
		x"0d",	--1004
		x"3e",	--1005
		x"00",	--1006
		x"3f",	--1007
		x"6e",	--1008
		x"b0",	--1009
		x"e0",	--1010
		x"8b",	--1011
		x"02",	--1012
		x"02",	--1013
		x"32",	--1014
		x"03",	--1015
		x"82",	--1016
		x"32",	--1017
		x"b2",	--1018
		x"18",	--1019
		x"38",	--1020
		x"9b",	--1021
		x"3a",	--1022
		x"06",	--1023
		x"32",	--1024
		x"0f",	--1025
		x"3a",	--1026
		x"3b",	--1027
		x"30",	--1028
		x"0b",	--1029
		x"09",	--1030
		x"08",	--1031
		x"8f",	--1032
		x"06",	--1033
		x"bf",	--1034
		x"00",	--1035
		x"08",	--1036
		x"2b",	--1037
		x"1e",	--1038
		x"02",	--1039
		x"0f",	--1040
		x"b0",	--1041
		x"7a",	--1042
		x"0c",	--1043
		x"3d",	--1044
		x"00",	--1045
		x"b0",	--1046
		x"26",	--1047
		x"08",	--1048
		x"09",	--1049
		x"1e",	--1050
		x"06",	--1051
		x"0f",	--1052
		x"b0",	--1053
		x"7a",	--1054
		x"0c",	--1055
		x"0d",	--1056
		x"0e",	--1057
		x"0f",	--1058
		x"b0",	--1059
		x"d6",	--1060
		x"b0",	--1061
		x"b6",	--1062
		x"8b",	--1063
		x"04",	--1064
		x"9b",	--1065
		x"00",	--1066
		x"38",	--1067
		x"39",	--1068
		x"3b",	--1069
		x"30",	--1070
		x"0b",	--1071
		x"0a",	--1072
		x"09",	--1073
		x"0a",	--1074
		x"0b",	--1075
		x"8f",	--1076
		x"06",	--1077
		x"8f",	--1078
		x"08",	--1079
		x"29",	--1080
		x"1e",	--1081
		x"02",	--1082
		x"0f",	--1083
		x"b0",	--1084
		x"7a",	--1085
		x"0c",	--1086
		x"0d",	--1087
		x"0e",	--1088
		x"0f",	--1089
		x"b0",	--1090
		x"26",	--1091
		x"0a",	--1092
		x"0b",	--1093
		x"1e",	--1094
		x"06",	--1095
		x"0f",	--1096
		x"b0",	--1097
		x"7a",	--1098
		x"0c",	--1099
		x"0d",	--1100
		x"0e",	--1101
		x"0f",	--1102
		x"b0",	--1103
		x"d6",	--1104
		x"b0",	--1105
		x"b6",	--1106
		x"89",	--1107
		x"04",	--1108
		x"39",	--1109
		x"3a",	--1110
		x"3b",	--1111
		x"30",	--1112
		x"2f",	--1113
		x"8f",	--1114
		x"04",	--1115
		x"30",	--1116
		x"0b",	--1117
		x"0a",	--1118
		x"92",	--1119
		x"10",	--1120
		x"14",	--1121
		x"3b",	--1122
		x"68",	--1123
		x"0a",	--1124
		x"2b",	--1125
		x"5f",	--1126
		x"fc",	--1127
		x"8f",	--1128
		x"0f",	--1129
		x"30",	--1130
		x"f7",	--1131
		x"b0",	--1132
		x"06",	--1133
		x"31",	--1134
		x"06",	--1135
		x"1a",	--1136
		x"3b",	--1137
		x"06",	--1138
		x"1a",	--1139
		x"10",	--1140
		x"ef",	--1141
		x"0f",	--1142
		x"3a",	--1143
		x"3b",	--1144
		x"30",	--1145
		x"1e",	--1146
		x"10",	--1147
		x"3e",	--1148
		x"20",	--1149
		x"12",	--1150
		x"0f",	--1151
		x"0f",	--1152
		x"0f",	--1153
		x"0f",	--1154
		x"3f",	--1155
		x"64",	--1156
		x"ff",	--1157
		x"68",	--1158
		x"00",	--1159
		x"bf",	--1160
		x"ba",	--1161
		x"02",	--1162
		x"bf",	--1163
		x"04",	--1164
		x"04",	--1165
		x"1e",	--1166
		x"82",	--1167
		x"10",	--1168
		x"30",	--1169
		x"0b",	--1170
		x"1b",	--1171
		x"10",	--1172
		x"3b",	--1173
		x"20",	--1174
		x"12",	--1175
		x"0c",	--1176
		x"0c",	--1177
		x"0c",	--1178
		x"0c",	--1179
		x"3c",	--1180
		x"64",	--1181
		x"cc",	--1182
		x"00",	--1183
		x"8c",	--1184
		x"02",	--1185
		x"8c",	--1186
		x"04",	--1187
		x"1b",	--1188
		x"82",	--1189
		x"10",	--1190
		x"0f",	--1191
		x"3b",	--1192
		x"30",	--1193
		x"3f",	--1194
		x"fc",	--1195
		x"0b",	--1196
		x"31",	--1197
		x"f0",	--1198
		x"1b",	--1199
		x"10",	--1200
		x"1b",	--1201
		x"0f",	--1202
		x"5f",	--1203
		x"64",	--1204
		x"16",	--1205
		x"3d",	--1206
		x"6a",	--1207
		x"0c",	--1208
		x"05",	--1209
		x"3d",	--1210
		x"06",	--1211
		x"cd",	--1212
		x"fa",	--1213
		x"0e",	--1214
		x"1c",	--1215
		x"0c",	--1216
		x"f8",	--1217
		x"30",	--1218
		x"ff",	--1219
		x"b0",	--1220
		x"06",	--1221
		x"21",	--1222
		x"3f",	--1223
		x"31",	--1224
		x"10",	--1225
		x"3b",	--1226
		x"30",	--1227
		x"0c",	--1228
		x"81",	--1229
		x"00",	--1230
		x"6d",	--1231
		x"4d",	--1232
		x"24",	--1233
		x"1e",	--1234
		x"1f",	--1235
		x"06",	--1236
		x"6d",	--1237
		x"4d",	--1238
		x"11",	--1239
		x"1e",	--1240
		x"3f",	--1241
		x"0e",	--1242
		x"7d",	--1243
		x"20",	--1244
		x"f7",	--1245
		x"ce",	--1246
		x"ff",	--1247
		x"0d",	--1248
		x"0d",	--1249
		x"0d",	--1250
		x"8d",	--1251
		x"00",	--1252
		x"1f",	--1253
		x"6d",	--1254
		x"4d",	--1255
		x"ef",	--1256
		x"0e",	--1257
		x"0e",	--1258
		x"0c",	--1259
		x"0c",	--1260
		x"3c",	--1261
		x"64",	--1262
		x"0e",	--1263
		x"9c",	--1264
		x"02",	--1265
		x"31",	--1266
		x"10",	--1267
		x"3b",	--1268
		x"30",	--1269
		x"1f",	--1270
		x"f1",	--1271
		x"b2",	--1272
		x"d2",	--1273
		x"60",	--1274
		x"b2",	--1275
		x"b8",	--1276
		x"72",	--1277
		x"0f",	--1278
		x"30",	--1279
		x"0b",	--1280
		x"0b",	--1281
		x"1f",	--1282
		x"12",	--1283
		x"3f",	--1284
		x"20",	--1285
		x"19",	--1286
		x"0c",	--1287
		x"0c",	--1288
		x"0d",	--1289
		x"0d",	--1290
		x"0d",	--1291
		x"0d",	--1292
		x"0d",	--1293
		x"3d",	--1294
		x"24",	--1295
		x"8d",	--1296
		x"00",	--1297
		x"8d",	--1298
		x"02",	--1299
		x"8d",	--1300
		x"08",	--1301
		x"8d",	--1302
		x"0a",	--1303
		x"8d",	--1304
		x"0c",	--1305
		x"0e",	--1306
		x"1e",	--1307
		x"82",	--1308
		x"12",	--1309
		x"3b",	--1310
		x"30",	--1311
		x"3f",	--1312
		x"fc",	--1313
		x"0f",	--1314
		x"0c",	--1315
		x"0c",	--1316
		x"0c",	--1317
		x"0c",	--1318
		x"0c",	--1319
		x"3c",	--1320
		x"24",	--1321
		x"8c",	--1322
		x"02",	--1323
		x"8c",	--1324
		x"04",	--1325
		x"8c",	--1326
		x"06",	--1327
		x"8c",	--1328
		x"08",	--1329
		x"9c",	--1330
		x"00",	--1331
		x"0f",	--1332
		x"30",	--1333
		x"0f",	--1334
		x"0e",	--1335
		x"0e",	--1336
		x"0e",	--1337
		x"0e",	--1338
		x"0e",	--1339
		x"8e",	--1340
		x"24",	--1341
		x"0f",	--1342
		x"30",	--1343
		x"0f",	--1344
		x"0e",	--1345
		x"0d",	--1346
		x"0c",	--1347
		x"0b",	--1348
		x"0a",	--1349
		x"09",	--1350
		x"08",	--1351
		x"07",	--1352
		x"92",	--1353
		x"12",	--1354
		x"33",	--1355
		x"3a",	--1356
		x"24",	--1357
		x"0b",	--1358
		x"2b",	--1359
		x"08",	--1360
		x"38",	--1361
		x"07",	--1362
		x"37",	--1363
		x"06",	--1364
		x"09",	--1365
		x"0f",	--1366
		x"1f",	--1367
		x"8b",	--1368
		x"00",	--1369
		x"19",	--1370
		x"3a",	--1371
		x"0e",	--1372
		x"3b",	--1373
		x"0e",	--1374
		x"38",	--1375
		x"0e",	--1376
		x"37",	--1377
		x"0e",	--1378
		x"19",	--1379
		x"12",	--1380
		x"19",	--1381
		x"8a",	--1382
		x"00",	--1383
		x"f1",	--1384
		x"2f",	--1385
		x"1f",	--1386
		x"02",	--1387
		x"ea",	--1388
		x"8b",	--1389
		x"00",	--1390
		x"1f",	--1391
		x"0a",	--1392
		x"9b",	--1393
		x"08",	--1394
		x"88",	--1395
		x"00",	--1396
		x"e4",	--1397
		x"2f",	--1398
		x"1f",	--1399
		x"87",	--1400
		x"00",	--1401
		x"2f",	--1402
		x"de",	--1403
		x"8a",	--1404
		x"00",	--1405
		x"db",	--1406
		x"b2",	--1407
		x"fe",	--1408
		x"60",	--1409
		x"37",	--1410
		x"38",	--1411
		x"39",	--1412
		x"3a",	--1413
		x"3b",	--1414
		x"3c",	--1415
		x"3d",	--1416
		x"3e",	--1417
		x"3f",	--1418
		x"00",	--1419
		x"8f",	--1420
		x"00",	--1421
		x"0f",	--1422
		x"30",	--1423
		x"2f",	--1424
		x"2e",	--1425
		x"1f",	--1426
		x"02",	--1427
		x"30",	--1428
		x"5e",	--1429
		x"81",	--1430
		x"3e",	--1431
		x"fc",	--1432
		x"c2",	--1433
		x"84",	--1434
		x"0f",	--1435
		x"30",	--1436
		x"3f",	--1437
		x"0f",	--1438
		x"5f",	--1439
		x"be",	--1440
		x"8f",	--1441
		x"b0",	--1442
		x"2a",	--1443
		x"30",	--1444
		x"0b",	--1445
		x"0b",	--1446
		x"0e",	--1447
		x"0e",	--1448
		x"0e",	--1449
		x"0e",	--1450
		x"0e",	--1451
		x"0f",	--1452
		x"b0",	--1453
		x"3a",	--1454
		x"0f",	--1455
		x"b0",	--1456
		x"3a",	--1457
		x"3b",	--1458
		x"30",	--1459
		x"0b",	--1460
		x"0a",	--1461
		x"0a",	--1462
		x"3b",	--1463
		x"07",	--1464
		x"0e",	--1465
		x"4d",	--1466
		x"7d",	--1467
		x"0f",	--1468
		x"03",	--1469
		x"0e",	--1470
		x"7d",	--1471
		x"fd",	--1472
		x"1e",	--1473
		x"0a",	--1474
		x"3f",	--1475
		x"31",	--1476
		x"b0",	--1477
		x"2a",	--1478
		x"3b",	--1479
		x"3b",	--1480
		x"ef",	--1481
		x"3a",	--1482
		x"3b",	--1483
		x"30",	--1484
		x"3f",	--1485
		x"30",	--1486
		x"f5",	--1487
		x"0b",	--1488
		x"0b",	--1489
		x"0e",	--1490
		x"8e",	--1491
		x"8e",	--1492
		x"0f",	--1493
		x"b0",	--1494
		x"4a",	--1495
		x"0f",	--1496
		x"b0",	--1497
		x"4a",	--1498
		x"3b",	--1499
		x"30",	--1500
		x"0b",	--1501
		x"0a",	--1502
		x"0a",	--1503
		x"0b",	--1504
		x"0d",	--1505
		x"8d",	--1506
		x"8d",	--1507
		x"0f",	--1508
		x"b0",	--1509
		x"4a",	--1510
		x"0f",	--1511
		x"b0",	--1512
		x"4a",	--1513
		x"0c",	--1514
		x"0d",	--1515
		x"8d",	--1516
		x"8c",	--1517
		x"4d",	--1518
		x"0d",	--1519
		x"0f",	--1520
		x"b0",	--1521
		x"4a",	--1522
		x"0f",	--1523
		x"b0",	--1524
		x"4a",	--1525
		x"3a",	--1526
		x"3b",	--1527
		x"30",	--1528
		x"0b",	--1529
		x"0a",	--1530
		x"09",	--1531
		x"0a",	--1532
		x"0e",	--1533
		x"19",	--1534
		x"09",	--1535
		x"39",	--1536
		x"0b",	--1537
		x"0d",	--1538
		x"0d",	--1539
		x"6f",	--1540
		x"8f",	--1541
		x"b0",	--1542
		x"4a",	--1543
		x"0b",	--1544
		x"0e",	--1545
		x"1b",	--1546
		x"3b",	--1547
		x"07",	--1548
		x"05",	--1549
		x"3f",	--1550
		x"20",	--1551
		x"b0",	--1552
		x"2a",	--1553
		x"ef",	--1554
		x"3f",	--1555
		x"3a",	--1556
		x"b0",	--1557
		x"2a",	--1558
		x"ea",	--1559
		x"39",	--1560
		x"3a",	--1561
		x"3b",	--1562
		x"30",	--1563
		x"0b",	--1564
		x"0a",	--1565
		x"09",	--1566
		x"0a",	--1567
		x"0e",	--1568
		x"17",	--1569
		x"09",	--1570
		x"39",	--1571
		x"0b",	--1572
		x"6f",	--1573
		x"8f",	--1574
		x"b0",	--1575
		x"3a",	--1576
		x"0b",	--1577
		x"0e",	--1578
		x"1b",	--1579
		x"3b",	--1580
		x"07",	--1581
		x"f6",	--1582
		x"3f",	--1583
		x"20",	--1584
		x"b0",	--1585
		x"2a",	--1586
		x"6f",	--1587
		x"8f",	--1588
		x"b0",	--1589
		x"3a",	--1590
		x"0b",	--1591
		x"f2",	--1592
		x"39",	--1593
		x"3a",	--1594
		x"3b",	--1595
		x"30",	--1596
		x"0b",	--1597
		x"0a",	--1598
		x"09",	--1599
		x"31",	--1600
		x"ec",	--1601
		x"0b",	--1602
		x"0f",	--1603
		x"34",	--1604
		x"3b",	--1605
		x"0a",	--1606
		x"38",	--1607
		x"09",	--1608
		x"0a",	--1609
		x"0a",	--1610
		x"3e",	--1611
		x"0a",	--1612
		x"0f",	--1613
		x"b0",	--1614
		x"98",	--1615
		x"7f",	--1616
		x"30",	--1617
		x"ca",	--1618
		x"00",	--1619
		x"19",	--1620
		x"3e",	--1621
		x"0a",	--1622
		x"0f",	--1623
		x"b0",	--1624
		x"66",	--1625
		x"0b",	--1626
		x"3f",	--1627
		x"0a",	--1628
		x"eb",	--1629
		x"0a",	--1630
		x"1a",	--1631
		x"09",	--1632
		x"3e",	--1633
		x"0a",	--1634
		x"0f",	--1635
		x"b0",	--1636
		x"98",	--1637
		x"7f",	--1638
		x"30",	--1639
		x"c9",	--1640
		x"00",	--1641
		x"3a",	--1642
		x"0f",	--1643
		x"0f",	--1644
		x"6f",	--1645
		x"8f",	--1646
		x"b0",	--1647
		x"2a",	--1648
		x"0a",	--1649
		x"f7",	--1650
		x"31",	--1651
		x"14",	--1652
		x"39",	--1653
		x"3a",	--1654
		x"3b",	--1655
		x"30",	--1656
		x"3f",	--1657
		x"2d",	--1658
		x"b0",	--1659
		x"2a",	--1660
		x"3b",	--1661
		x"1b",	--1662
		x"c5",	--1663
		x"1a",	--1664
		x"09",	--1665
		x"dd",	--1666
		x"0b",	--1667
		x"0a",	--1668
		x"09",	--1669
		x"0b",	--1670
		x"3b",	--1671
		x"39",	--1672
		x"6f",	--1673
		x"4f",	--1674
		x"0b",	--1675
		x"1a",	--1676
		x"8f",	--1677
		x"b0",	--1678
		x"2a",	--1679
		x"0a",	--1680
		x"09",	--1681
		x"19",	--1682
		x"5f",	--1683
		x"01",	--1684
		x"4f",	--1685
		x"10",	--1686
		x"7f",	--1687
		x"25",	--1688
		x"f3",	--1689
		x"0a",	--1690
		x"1a",	--1691
		x"5f",	--1692
		x"01",	--1693
		x"7f",	--1694
		x"db",	--1695
		x"7f",	--1696
		x"54",	--1697
		x"ee",	--1698
		x"4f",	--1699
		x"0f",	--1700
		x"10",	--1701
		x"16",	--1702
		x"39",	--1703
		x"3a",	--1704
		x"3b",	--1705
		x"30",	--1706
		x"09",	--1707
		x"29",	--1708
		x"1e",	--1709
		x"02",	--1710
		x"2f",	--1711
		x"b0",	--1712
		x"f2",	--1713
		x"0b",	--1714
		x"dd",	--1715
		x"09",	--1716
		x"29",	--1717
		x"2f",	--1718
		x"b0",	--1719
		x"a0",	--1720
		x"0b",	--1721
		x"d6",	--1722
		x"0f",	--1723
		x"2b",	--1724
		x"29",	--1725
		x"6f",	--1726
		x"4f",	--1727
		x"d0",	--1728
		x"19",	--1729
		x"8f",	--1730
		x"b0",	--1731
		x"2a",	--1732
		x"7f",	--1733
		x"4f",	--1734
		x"fa",	--1735
		x"c8",	--1736
		x"09",	--1737
		x"29",	--1738
		x"1e",	--1739
		x"02",	--1740
		x"2f",	--1741
		x"b0",	--1742
		x"38",	--1743
		x"0b",	--1744
		x"bf",	--1745
		x"09",	--1746
		x"29",	--1747
		x"2e",	--1748
		x"0f",	--1749
		x"8f",	--1750
		x"8f",	--1751
		x"8f",	--1752
		x"8f",	--1753
		x"b0",	--1754
		x"ba",	--1755
		x"0b",	--1756
		x"b3",	--1757
		x"09",	--1758
		x"29",	--1759
		x"2f",	--1760
		x"b0",	--1761
		x"7a",	--1762
		x"0b",	--1763
		x"ac",	--1764
		x"09",	--1765
		x"29",	--1766
		x"2f",	--1767
		x"b0",	--1768
		x"2a",	--1769
		x"0b",	--1770
		x"a5",	--1771
		x"09",	--1772
		x"29",	--1773
		x"2f",	--1774
		x"b0",	--1775
		x"4a",	--1776
		x"0b",	--1777
		x"9e",	--1778
		x"09",	--1779
		x"29",	--1780
		x"2f",	--1781
		x"b0",	--1782
		x"68",	--1783
		x"0b",	--1784
		x"97",	--1785
		x"3f",	--1786
		x"25",	--1787
		x"b0",	--1788
		x"2a",	--1789
		x"92",	--1790
		x"0f",	--1791
		x"0e",	--1792
		x"1f",	--1793
		x"14",	--1794
		x"df",	--1795
		x"85",	--1796
		x"e4",	--1797
		x"1f",	--1798
		x"14",	--1799
		x"3f",	--1800
		x"3f",	--1801
		x"13",	--1802
		x"92",	--1803
		x"14",	--1804
		x"1e",	--1805
		x"14",	--1806
		x"1f",	--1807
		x"16",	--1808
		x"0e",	--1809
		x"02",	--1810
		x"92",	--1811
		x"16",	--1812
		x"f2",	--1813
		x"10",	--1814
		x"81",	--1815
		x"3e",	--1816
		x"3f",	--1817
		x"b1",	--1818
		x"f0",	--1819
		x"00",	--1820
		x"00",	--1821
		x"82",	--1822
		x"14",	--1823
		x"ec",	--1824
		x"0c",	--1825
		x"0d",	--1826
		x"3e",	--1827
		x"00",	--1828
		x"3f",	--1829
		x"6e",	--1830
		x"b0",	--1831
		x"a0",	--1832
		x"3e",	--1833
		x"82",	--1834
		x"82",	--1835
		x"f2",	--1836
		x"11",	--1837
		x"80",	--1838
		x"30",	--1839
		x"1e",	--1840
		x"14",	--1841
		x"1f",	--1842
		x"16",	--1843
		x"0e",	--1844
		x"05",	--1845
		x"1f",	--1846
		x"14",	--1847
		x"1f",	--1848
		x"16",	--1849
		x"30",	--1850
		x"1d",	--1851
		x"14",	--1852
		x"1e",	--1853
		x"16",	--1854
		x"3f",	--1855
		x"40",	--1856
		x"0f",	--1857
		x"0f",	--1858
		x"30",	--1859
		x"1f",	--1860
		x"16",	--1861
		x"5f",	--1862
		x"e4",	--1863
		x"1d",	--1864
		x"16",	--1865
		x"1e",	--1866
		x"14",	--1867
		x"0d",	--1868
		x"0b",	--1869
		x"1e",	--1870
		x"16",	--1871
		x"3e",	--1872
		x"3f",	--1873
		x"03",	--1874
		x"82",	--1875
		x"16",	--1876
		x"30",	--1877
		x"92",	--1878
		x"16",	--1879
		x"30",	--1880
		x"4f",	--1881
		x"30",	--1882
		x"0b",	--1883
		x"0a",	--1884
		x"0a",	--1885
		x"0b",	--1886
		x"0c",	--1887
		x"3d",	--1888
		x"00",	--1889
		x"b0",	--1890
		x"9a",	--1891
		x"0f",	--1892
		x"07",	--1893
		x"0e",	--1894
		x"0f",	--1895
		x"b0",	--1896
		x"ea",	--1897
		x"3a",	--1898
		x"3b",	--1899
		x"30",	--1900
		x"0c",	--1901
		x"3d",	--1902
		x"00",	--1903
		x"0e",	--1904
		x"0f",	--1905
		x"b0",	--1906
		x"d6",	--1907
		x"b0",	--1908
		x"ea",	--1909
		x"0e",	--1910
		x"3f",	--1911
		x"00",	--1912
		x"3a",	--1913
		x"3b",	--1914
		x"30",	--1915
		x"0b",	--1916
		x"0a",	--1917
		x"09",	--1918
		x"08",	--1919
		x"07",	--1920
		x"06",	--1921
		x"05",	--1922
		x"04",	--1923
		x"31",	--1924
		x"fa",	--1925
		x"08",	--1926
		x"6b",	--1927
		x"6b",	--1928
		x"67",	--1929
		x"6c",	--1930
		x"6c",	--1931
		x"e9",	--1932
		x"6b",	--1933
		x"02",	--1934
		x"30",	--1935
		x"78",	--1936
		x"6c",	--1937
		x"e3",	--1938
		x"6c",	--1939
		x"bb",	--1940
		x"6b",	--1941
		x"df",	--1942
		x"91",	--1943
		x"02",	--1944
		x"00",	--1945
		x"1b",	--1946
		x"02",	--1947
		x"14",	--1948
		x"04",	--1949
		x"15",	--1950
		x"06",	--1951
		x"16",	--1952
		x"04",	--1953
		x"17",	--1954
		x"06",	--1955
		x"2c",	--1956
		x"0c",	--1957
		x"09",	--1958
		x"0c",	--1959
		x"bf",	--1960
		x"39",	--1961
		x"20",	--1962
		x"50",	--1963
		x"1c",	--1964
		x"d7",	--1965
		x"81",	--1966
		x"02",	--1967
		x"81",	--1968
		x"04",	--1969
		x"4c",	--1970
		x"7c",	--1971
		x"1f",	--1972
		x"0b",	--1973
		x"0a",	--1974
		x"0b",	--1975
		x"12",	--1976
		x"0b",	--1977
		x"0a",	--1978
		x"7c",	--1979
		x"fb",	--1980
		x"81",	--1981
		x"02",	--1982
		x"81",	--1983
		x"04",	--1984
		x"1c",	--1985
		x"0d",	--1986
		x"79",	--1987
		x"1f",	--1988
		x"04",	--1989
		x"0c",	--1990
		x"0d",	--1991
		x"79",	--1992
		x"fc",	--1993
		x"3c",	--1994
		x"3d",	--1995
		x"0c",	--1996
		x"0d",	--1997
		x"1a",	--1998
		x"0b",	--1999
		x"0c",	--2000
		x"02",	--2001
		x"0d",	--2002
		x"e5",	--2003
		x"16",	--2004
		x"02",	--2005
		x"17",	--2006
		x"04",	--2007
		x"06",	--2008
		x"07",	--2009
		x"5f",	--2010
		x"01",	--2011
		x"5f",	--2012
		x"01",	--2013
		x"28",	--2014
		x"c8",	--2015
		x"01",	--2016
		x"a8",	--2017
		x"02",	--2018
		x"0e",	--2019
		x"0f",	--2020
		x"0e",	--2021
		x"0f",	--2022
		x"88",	--2023
		x"04",	--2024
		x"88",	--2025
		x"06",	--2026
		x"f8",	--2027
		x"03",	--2028
		x"00",	--2029
		x"0f",	--2030
		x"4d",	--2031
		x"0f",	--2032
		x"31",	--2033
		x"06",	--2034
		x"34",	--2035
		x"35",	--2036
		x"36",	--2037
		x"37",	--2038
		x"38",	--2039
		x"39",	--2040
		x"3a",	--2041
		x"3b",	--2042
		x"30",	--2043
		x"2b",	--2044
		x"67",	--2045
		x"81",	--2046
		x"00",	--2047
		x"04",	--2048
		x"05",	--2049
		x"5f",	--2050
		x"01",	--2051
		x"5f",	--2052
		x"01",	--2053
		x"d8",	--2054
		x"4f",	--2055
		x"68",	--2056
		x"0e",	--2057
		x"0f",	--2058
		x"0e",	--2059
		x"0f",	--2060
		x"0f",	--2061
		x"69",	--2062
		x"c8",	--2063
		x"01",	--2064
		x"a8",	--2065
		x"02",	--2066
		x"88",	--2067
		x"04",	--2068
		x"88",	--2069
		x"06",	--2070
		x"0c",	--2071
		x"0d",	--2072
		x"3c",	--2073
		x"3d",	--2074
		x"3d",	--2075
		x"ff",	--2076
		x"05",	--2077
		x"3d",	--2078
		x"00",	--2079
		x"17",	--2080
		x"3c",	--2081
		x"15",	--2082
		x"1b",	--2083
		x"02",	--2084
		x"3b",	--2085
		x"0e",	--2086
		x"0f",	--2087
		x"0a",	--2088
		x"3b",	--2089
		x"0c",	--2090
		x"0d",	--2091
		x"3c",	--2092
		x"3d",	--2093
		x"3d",	--2094
		x"ff",	--2095
		x"f5",	--2096
		x"3c",	--2097
		x"88",	--2098
		x"04",	--2099
		x"88",	--2100
		x"06",	--2101
		x"88",	--2102
		x"02",	--2103
		x"f8",	--2104
		x"03",	--2105
		x"00",	--2106
		x"0f",	--2107
		x"b3",	--2108
		x"0c",	--2109
		x"0d",	--2110
		x"1c",	--2111
		x"0d",	--2112
		x"12",	--2113
		x"0f",	--2114
		x"0e",	--2115
		x"0a",	--2116
		x"0b",	--2117
		x"0a",	--2118
		x"0b",	--2119
		x"88",	--2120
		x"04",	--2121
		x"88",	--2122
		x"06",	--2123
		x"98",	--2124
		x"02",	--2125
		x"0f",	--2126
		x"a1",	--2127
		x"6b",	--2128
		x"9f",	--2129
		x"ad",	--2130
		x"00",	--2131
		x"9d",	--2132
		x"02",	--2133
		x"02",	--2134
		x"9d",	--2135
		x"04",	--2136
		x"04",	--2137
		x"9d",	--2138
		x"06",	--2139
		x"06",	--2140
		x"5e",	--2141
		x"01",	--2142
		x"5e",	--2143
		x"01",	--2144
		x"cd",	--2145
		x"01",	--2146
		x"0f",	--2147
		x"8c",	--2148
		x"06",	--2149
		x"07",	--2150
		x"9a",	--2151
		x"39",	--2152
		x"19",	--2153
		x"39",	--2154
		x"20",	--2155
		x"8f",	--2156
		x"3e",	--2157
		x"3c",	--2158
		x"b6",	--2159
		x"c1",	--2160
		x"0e",	--2161
		x"0f",	--2162
		x"0e",	--2163
		x"0f",	--2164
		x"97",	--2165
		x"0f",	--2166
		x"79",	--2167
		x"d8",	--2168
		x"01",	--2169
		x"a8",	--2170
		x"02",	--2171
		x"3e",	--2172
		x"3f",	--2173
		x"1e",	--2174
		x"0f",	--2175
		x"88",	--2176
		x"04",	--2177
		x"88",	--2178
		x"06",	--2179
		x"92",	--2180
		x"0c",	--2181
		x"7b",	--2182
		x"81",	--2183
		x"00",	--2184
		x"81",	--2185
		x"02",	--2186
		x"81",	--2187
		x"04",	--2188
		x"4d",	--2189
		x"7d",	--2190
		x"1f",	--2191
		x"0c",	--2192
		x"4b",	--2193
		x"0c",	--2194
		x"0d",	--2195
		x"12",	--2196
		x"0d",	--2197
		x"0c",	--2198
		x"7b",	--2199
		x"fb",	--2200
		x"81",	--2201
		x"02",	--2202
		x"81",	--2203
		x"04",	--2204
		x"1c",	--2205
		x"0d",	--2206
		x"79",	--2207
		x"1f",	--2208
		x"04",	--2209
		x"0c",	--2210
		x"0d",	--2211
		x"79",	--2212
		x"fc",	--2213
		x"3c",	--2214
		x"3d",	--2215
		x"0c",	--2216
		x"0d",	--2217
		x"1a",	--2218
		x"0b",	--2219
		x"0c",	--2220
		x"04",	--2221
		x"0d",	--2222
		x"02",	--2223
		x"0a",	--2224
		x"0b",	--2225
		x"14",	--2226
		x"02",	--2227
		x"15",	--2228
		x"04",	--2229
		x"04",	--2230
		x"05",	--2231
		x"49",	--2232
		x"0a",	--2233
		x"0b",	--2234
		x"18",	--2235
		x"6c",	--2236
		x"33",	--2237
		x"df",	--2238
		x"01",	--2239
		x"01",	--2240
		x"2f",	--2241
		x"3f",	--2242
		x"d0",	--2243
		x"2c",	--2244
		x"31",	--2245
		x"e0",	--2246
		x"81",	--2247
		x"04",	--2248
		x"81",	--2249
		x"06",	--2250
		x"81",	--2251
		x"00",	--2252
		x"81",	--2253
		x"02",	--2254
		x"0e",	--2255
		x"3e",	--2256
		x"18",	--2257
		x"0f",	--2258
		x"2f",	--2259
		x"b0",	--2260
		x"ac",	--2261
		x"0e",	--2262
		x"3e",	--2263
		x"10",	--2264
		x"0f",	--2265
		x"b0",	--2266
		x"ac",	--2267
		x"0d",	--2268
		x"3d",	--2269
		x"0e",	--2270
		x"3e",	--2271
		x"10",	--2272
		x"0f",	--2273
		x"3f",	--2274
		x"18",	--2275
		x"b0",	--2276
		x"f8",	--2277
		x"b0",	--2278
		x"ce",	--2279
		x"31",	--2280
		x"20",	--2281
		x"30",	--2282
		x"31",	--2283
		x"e0",	--2284
		x"81",	--2285
		x"04",	--2286
		x"81",	--2287
		x"06",	--2288
		x"81",	--2289
		x"00",	--2290
		x"81",	--2291
		x"02",	--2292
		x"0e",	--2293
		x"3e",	--2294
		x"18",	--2295
		x"0f",	--2296
		x"2f",	--2297
		x"b0",	--2298
		x"ac",	--2299
		x"0e",	--2300
		x"3e",	--2301
		x"10",	--2302
		x"0f",	--2303
		x"b0",	--2304
		x"ac",	--2305
		x"d1",	--2306
		x"11",	--2307
		x"0d",	--2308
		x"3d",	--2309
		x"0e",	--2310
		x"3e",	--2311
		x"10",	--2312
		x"0f",	--2313
		x"3f",	--2314
		x"18",	--2315
		x"b0",	--2316
		x"f8",	--2317
		x"b0",	--2318
		x"ce",	--2319
		x"31",	--2320
		x"20",	--2321
		x"30",	--2322
		x"0b",	--2323
		x"0a",	--2324
		x"09",	--2325
		x"08",	--2326
		x"07",	--2327
		x"06",	--2328
		x"05",	--2329
		x"04",	--2330
		x"31",	--2331
		x"dc",	--2332
		x"81",	--2333
		x"04",	--2334
		x"81",	--2335
		x"06",	--2336
		x"81",	--2337
		x"00",	--2338
		x"81",	--2339
		x"02",	--2340
		x"0e",	--2341
		x"3e",	--2342
		x"18",	--2343
		x"0f",	--2344
		x"2f",	--2345
		x"b0",	--2346
		x"ac",	--2347
		x"0e",	--2348
		x"3e",	--2349
		x"10",	--2350
		x"0f",	--2351
		x"b0",	--2352
		x"ac",	--2353
		x"5f",	--2354
		x"18",	--2355
		x"6f",	--2356
		x"b6",	--2357
		x"5e",	--2358
		x"10",	--2359
		x"6e",	--2360
		x"d9",	--2361
		x"6f",	--2362
		x"ae",	--2363
		x"6e",	--2364
		x"e2",	--2365
		x"6f",	--2366
		x"ac",	--2367
		x"6e",	--2368
		x"d1",	--2369
		x"14",	--2370
		x"1c",	--2371
		x"15",	--2372
		x"1e",	--2373
		x"18",	--2374
		x"14",	--2375
		x"19",	--2376
		x"16",	--2377
		x"3c",	--2378
		x"20",	--2379
		x"0e",	--2380
		x"0f",	--2381
		x"06",	--2382
		x"07",	--2383
		x"81",	--2384
		x"20",	--2385
		x"81",	--2386
		x"22",	--2387
		x"0a",	--2388
		x"0b",	--2389
		x"81",	--2390
		x"20",	--2391
		x"08",	--2392
		x"08",	--2393
		x"09",	--2394
		x"12",	--2395
		x"05",	--2396
		x"04",	--2397
		x"b1",	--2398
		x"20",	--2399
		x"19",	--2400
		x"14",	--2401
		x"0d",	--2402
		x"0a",	--2403
		x"0b",	--2404
		x"0e",	--2405
		x"0f",	--2406
		x"1c",	--2407
		x"0d",	--2408
		x"0b",	--2409
		x"03",	--2410
		x"0b",	--2411
		x"0c",	--2412
		x"0d",	--2413
		x"0e",	--2414
		x"0f",	--2415
		x"06",	--2416
		x"07",	--2417
		x"09",	--2418
		x"e5",	--2419
		x"16",	--2420
		x"07",	--2421
		x"e2",	--2422
		x"0a",	--2423
		x"f5",	--2424
		x"f2",	--2425
		x"81",	--2426
		x"20",	--2427
		x"81",	--2428
		x"22",	--2429
		x"0c",	--2430
		x"1a",	--2431
		x"1a",	--2432
		x"1a",	--2433
		x"12",	--2434
		x"06",	--2435
		x"26",	--2436
		x"81",	--2437
		x"0a",	--2438
		x"5d",	--2439
		x"d1",	--2440
		x"11",	--2441
		x"19",	--2442
		x"83",	--2443
		x"c1",	--2444
		x"09",	--2445
		x"0c",	--2446
		x"3c",	--2447
		x"3f",	--2448
		x"00",	--2449
		x"18",	--2450
		x"1d",	--2451
		x"0a",	--2452
		x"3d",	--2453
		x"1a",	--2454
		x"20",	--2455
		x"1b",	--2456
		x"22",	--2457
		x"0c",	--2458
		x"0e",	--2459
		x"0f",	--2460
		x"0b",	--2461
		x"2a",	--2462
		x"0a",	--2463
		x"0b",	--2464
		x"3d",	--2465
		x"3f",	--2466
		x"00",	--2467
		x"f5",	--2468
		x"81",	--2469
		x"20",	--2470
		x"81",	--2471
		x"22",	--2472
		x"81",	--2473
		x"0a",	--2474
		x"0c",	--2475
		x"0d",	--2476
		x"3c",	--2477
		x"7f",	--2478
		x"0d",	--2479
		x"3c",	--2480
		x"40",	--2481
		x"44",	--2482
		x"81",	--2483
		x"0c",	--2484
		x"81",	--2485
		x"0e",	--2486
		x"f1",	--2487
		x"03",	--2488
		x"08",	--2489
		x"0f",	--2490
		x"3f",	--2491
		x"b0",	--2492
		x"ce",	--2493
		x"31",	--2494
		x"24",	--2495
		x"34",	--2496
		x"35",	--2497
		x"36",	--2498
		x"37",	--2499
		x"38",	--2500
		x"39",	--2501
		x"3a",	--2502
		x"3b",	--2503
		x"30",	--2504
		x"1e",	--2505
		x"0f",	--2506
		x"d3",	--2507
		x"3a",	--2508
		x"03",	--2509
		x"08",	--2510
		x"1e",	--2511
		x"10",	--2512
		x"1c",	--2513
		x"20",	--2514
		x"1d",	--2515
		x"22",	--2516
		x"12",	--2517
		x"0d",	--2518
		x"0c",	--2519
		x"06",	--2520
		x"07",	--2521
		x"06",	--2522
		x"37",	--2523
		x"00",	--2524
		x"81",	--2525
		x"20",	--2526
		x"81",	--2527
		x"22",	--2528
		x"12",	--2529
		x"0f",	--2530
		x"0e",	--2531
		x"1a",	--2532
		x"0f",	--2533
		x"e7",	--2534
		x"81",	--2535
		x"0a",	--2536
		x"a6",	--2537
		x"6e",	--2538
		x"36",	--2539
		x"5f",	--2540
		x"d1",	--2541
		x"11",	--2542
		x"19",	--2543
		x"20",	--2544
		x"c1",	--2545
		x"19",	--2546
		x"0f",	--2547
		x"3f",	--2548
		x"18",	--2549
		x"c5",	--2550
		x"0d",	--2551
		x"ba",	--2552
		x"0c",	--2553
		x"0d",	--2554
		x"3c",	--2555
		x"80",	--2556
		x"0d",	--2557
		x"0c",	--2558
		x"b3",	--2559
		x"0d",	--2560
		x"b1",	--2561
		x"81",	--2562
		x"20",	--2563
		x"03",	--2564
		x"81",	--2565
		x"22",	--2566
		x"ab",	--2567
		x"3e",	--2568
		x"40",	--2569
		x"0f",	--2570
		x"3e",	--2571
		x"80",	--2572
		x"3f",	--2573
		x"a4",	--2574
		x"4d",	--2575
		x"7b",	--2576
		x"4f",	--2577
		x"de",	--2578
		x"5f",	--2579
		x"d1",	--2580
		x"11",	--2581
		x"19",	--2582
		x"06",	--2583
		x"c1",	--2584
		x"11",	--2585
		x"0f",	--2586
		x"3f",	--2587
		x"10",	--2588
		x"9e",	--2589
		x"4f",	--2590
		x"f8",	--2591
		x"6f",	--2592
		x"f1",	--2593
		x"3f",	--2594
		x"d0",	--2595
		x"97",	--2596
		x"0b",	--2597
		x"0a",	--2598
		x"09",	--2599
		x"08",	--2600
		x"07",	--2601
		x"31",	--2602
		x"e8",	--2603
		x"81",	--2604
		x"04",	--2605
		x"81",	--2606
		x"06",	--2607
		x"81",	--2608
		x"00",	--2609
		x"81",	--2610
		x"02",	--2611
		x"0e",	--2612
		x"3e",	--2613
		x"10",	--2614
		x"0f",	--2615
		x"2f",	--2616
		x"b0",	--2617
		x"ac",	--2618
		x"0e",	--2619
		x"3e",	--2620
		x"0f",	--2621
		x"b0",	--2622
		x"ac",	--2623
		x"5f",	--2624
		x"10",	--2625
		x"6f",	--2626
		x"5d",	--2627
		x"5e",	--2628
		x"08",	--2629
		x"6e",	--2630
		x"82",	--2631
		x"d1",	--2632
		x"09",	--2633
		x"11",	--2634
		x"6f",	--2635
		x"58",	--2636
		x"6f",	--2637
		x"56",	--2638
		x"6e",	--2639
		x"6f",	--2640
		x"6e",	--2641
		x"4c",	--2642
		x"1d",	--2643
		x"12",	--2644
		x"1d",	--2645
		x"0a",	--2646
		x"81",	--2647
		x"12",	--2648
		x"1e",	--2649
		x"14",	--2650
		x"1f",	--2651
		x"16",	--2652
		x"18",	--2653
		x"0c",	--2654
		x"19",	--2655
		x"0e",	--2656
		x"0f",	--2657
		x"1e",	--2658
		x"0e",	--2659
		x"0f",	--2660
		x"3d",	--2661
		x"81",	--2662
		x"12",	--2663
		x"37",	--2664
		x"1f",	--2665
		x"0c",	--2666
		x"3d",	--2667
		x"00",	--2668
		x"0a",	--2669
		x"0b",	--2670
		x"0b",	--2671
		x"0a",	--2672
		x"0b",	--2673
		x"0e",	--2674
		x"0f",	--2675
		x"12",	--2676
		x"0d",	--2677
		x"0c",	--2678
		x"0e",	--2679
		x"0f",	--2680
		x"37",	--2681
		x"0b",	--2682
		x"0f",	--2683
		x"f7",	--2684
		x"f2",	--2685
		x"0e",	--2686
		x"f4",	--2687
		x"ef",	--2688
		x"09",	--2689
		x"e5",	--2690
		x"0e",	--2691
		x"e3",	--2692
		x"dd",	--2693
		x"0c",	--2694
		x"0d",	--2695
		x"3c",	--2696
		x"7f",	--2697
		x"0d",	--2698
		x"3c",	--2699
		x"40",	--2700
		x"1c",	--2701
		x"81",	--2702
		x"14",	--2703
		x"81",	--2704
		x"16",	--2705
		x"0f",	--2706
		x"3f",	--2707
		x"10",	--2708
		x"b0",	--2709
		x"ce",	--2710
		x"31",	--2711
		x"18",	--2712
		x"37",	--2713
		x"38",	--2714
		x"39",	--2715
		x"3a",	--2716
		x"3b",	--2717
		x"30",	--2718
		x"e1",	--2719
		x"10",	--2720
		x"0f",	--2721
		x"3f",	--2722
		x"10",	--2723
		x"f0",	--2724
		x"4f",	--2725
		x"fa",	--2726
		x"3f",	--2727
		x"d0",	--2728
		x"eb",	--2729
		x"0d",	--2730
		x"e2",	--2731
		x"0c",	--2732
		x"0d",	--2733
		x"3c",	--2734
		x"80",	--2735
		x"0d",	--2736
		x"0c",	--2737
		x"db",	--2738
		x"0d",	--2739
		x"d9",	--2740
		x"0e",	--2741
		x"02",	--2742
		x"0f",	--2743
		x"d5",	--2744
		x"3a",	--2745
		x"40",	--2746
		x"0b",	--2747
		x"3a",	--2748
		x"80",	--2749
		x"3b",	--2750
		x"ce",	--2751
		x"81",	--2752
		x"14",	--2753
		x"81",	--2754
		x"16",	--2755
		x"81",	--2756
		x"12",	--2757
		x"0f",	--2758
		x"3f",	--2759
		x"10",	--2760
		x"cb",	--2761
		x"0f",	--2762
		x"3f",	--2763
		x"c8",	--2764
		x"31",	--2765
		x"e8",	--2766
		x"81",	--2767
		x"04",	--2768
		x"81",	--2769
		x"06",	--2770
		x"81",	--2771
		x"00",	--2772
		x"81",	--2773
		x"02",	--2774
		x"0e",	--2775
		x"3e",	--2776
		x"10",	--2777
		x"0f",	--2778
		x"2f",	--2779
		x"b0",	--2780
		x"ac",	--2781
		x"0e",	--2782
		x"3e",	--2783
		x"0f",	--2784
		x"b0",	--2785
		x"ac",	--2786
		x"e1",	--2787
		x"10",	--2788
		x"0d",	--2789
		x"e1",	--2790
		x"08",	--2791
		x"0a",	--2792
		x"0e",	--2793
		x"3e",	--2794
		x"0f",	--2795
		x"3f",	--2796
		x"10",	--2797
		x"b0",	--2798
		x"d0",	--2799
		x"31",	--2800
		x"18",	--2801
		x"30",	--2802
		x"3f",	--2803
		x"fb",	--2804
		x"31",	--2805
		x"f4",	--2806
		x"81",	--2807
		x"00",	--2808
		x"81",	--2809
		x"02",	--2810
		x"0e",	--2811
		x"2e",	--2812
		x"0f",	--2813
		x"b0",	--2814
		x"ac",	--2815
		x"5f",	--2816
		x"04",	--2817
		x"6f",	--2818
		x"28",	--2819
		x"27",	--2820
		x"6f",	--2821
		x"07",	--2822
		x"1d",	--2823
		x"06",	--2824
		x"0d",	--2825
		x"21",	--2826
		x"3d",	--2827
		x"1f",	--2828
		x"09",	--2829
		x"c1",	--2830
		x"05",	--2831
		x"26",	--2832
		x"3e",	--2833
		x"3f",	--2834
		x"ff",	--2835
		x"31",	--2836
		x"0c",	--2837
		x"30",	--2838
		x"1e",	--2839
		x"08",	--2840
		x"1f",	--2841
		x"0a",	--2842
		x"3c",	--2843
		x"1e",	--2844
		x"4c",	--2845
		x"4d",	--2846
		x"7d",	--2847
		x"1f",	--2848
		x"0f",	--2849
		x"c1",	--2850
		x"05",	--2851
		x"ef",	--2852
		x"3e",	--2853
		x"3f",	--2854
		x"1e",	--2855
		x"0f",	--2856
		x"31",	--2857
		x"0c",	--2858
		x"30",	--2859
		x"0e",	--2860
		x"0f",	--2861
		x"31",	--2862
		x"0c",	--2863
		x"30",	--2864
		x"12",	--2865
		x"0f",	--2866
		x"0e",	--2867
		x"7d",	--2868
		x"fb",	--2869
		x"eb",	--2870
		x"0e",	--2871
		x"3f",	--2872
		x"00",	--2873
		x"31",	--2874
		x"0c",	--2875
		x"30",	--2876
		x"0b",	--2877
		x"0a",	--2878
		x"09",	--2879
		x"08",	--2880
		x"31",	--2881
		x"0a",	--2882
		x"0b",	--2883
		x"c1",	--2884
		x"01",	--2885
		x"0e",	--2886
		x"0d",	--2887
		x"0b",	--2888
		x"0b",	--2889
		x"e1",	--2890
		x"00",	--2891
		x"0f",	--2892
		x"b0",	--2893
		x"ce",	--2894
		x"31",	--2895
		x"38",	--2896
		x"39",	--2897
		x"3a",	--2898
		x"3b",	--2899
		x"30",	--2900
		x"f1",	--2901
		x"03",	--2902
		x"00",	--2903
		x"b1",	--2904
		x"1e",	--2905
		x"02",	--2906
		x"81",	--2907
		x"04",	--2908
		x"81",	--2909
		x"06",	--2910
		x"0e",	--2911
		x"0f",	--2912
		x"b0",	--2913
		x"5c",	--2914
		x"3f",	--2915
		x"0f",	--2916
		x"18",	--2917
		x"e5",	--2918
		x"81",	--2919
		x"04",	--2920
		x"81",	--2921
		x"06",	--2922
		x"4e",	--2923
		x"7e",	--2924
		x"1f",	--2925
		x"06",	--2926
		x"3e",	--2927
		x"1e",	--2928
		x"0e",	--2929
		x"81",	--2930
		x"02",	--2931
		x"d7",	--2932
		x"91",	--2933
		x"04",	--2934
		x"04",	--2935
		x"91",	--2936
		x"06",	--2937
		x"06",	--2938
		x"7e",	--2939
		x"f8",	--2940
		x"f1",	--2941
		x"0e",	--2942
		x"3e",	--2943
		x"1e",	--2944
		x"1c",	--2945
		x"0d",	--2946
		x"48",	--2947
		x"78",	--2948
		x"1f",	--2949
		x"04",	--2950
		x"0c",	--2951
		x"0d",	--2952
		x"78",	--2953
		x"fc",	--2954
		x"3c",	--2955
		x"3d",	--2956
		x"0c",	--2957
		x"0d",	--2958
		x"18",	--2959
		x"09",	--2960
		x"0c",	--2961
		x"04",	--2962
		x"0d",	--2963
		x"02",	--2964
		x"08",	--2965
		x"09",	--2966
		x"7e",	--2967
		x"1f",	--2968
		x"0e",	--2969
		x"0d",	--2970
		x"0e",	--2971
		x"0d",	--2972
		x"0e",	--2973
		x"81",	--2974
		x"04",	--2975
		x"81",	--2976
		x"06",	--2977
		x"3e",	--2978
		x"1e",	--2979
		x"0e",	--2980
		x"81",	--2981
		x"02",	--2982
		x"a4",	--2983
		x"12",	--2984
		x"0b",	--2985
		x"0a",	--2986
		x"7e",	--2987
		x"fb",	--2988
		x"ec",	--2989
		x"0b",	--2990
		x"0a",	--2991
		x"09",	--2992
		x"1f",	--2993
		x"17",	--2994
		x"3e",	--2995
		x"00",	--2996
		x"2c",	--2997
		x"3a",	--2998
		x"18",	--2999
		x"0b",	--3000
		x"39",	--3001
		x"0c",	--3002
		x"0d",	--3003
		x"4f",	--3004
		x"4f",	--3005
		x"17",	--3006
		x"3c",	--3007
		x"d8",	--3008
		x"6e",	--3009
		x"0f",	--3010
		x"0a",	--3011
		x"0b",	--3012
		x"0f",	--3013
		x"39",	--3014
		x"3a",	--3015
		x"3b",	--3016
		x"30",	--3017
		x"3f",	--3018
		x"00",	--3019
		x"0f",	--3020
		x"3a",	--3021
		x"0b",	--3022
		x"39",	--3023
		x"18",	--3024
		x"0c",	--3025
		x"0d",	--3026
		x"4f",	--3027
		x"4f",	--3028
		x"e9",	--3029
		x"12",	--3030
		x"0d",	--3031
		x"0c",	--3032
		x"7f",	--3033
		x"fb",	--3034
		x"e3",	--3035
		x"3a",	--3036
		x"10",	--3037
		x"0b",	--3038
		x"39",	--3039
		x"10",	--3040
		x"ef",	--3041
		x"3a",	--3042
		x"20",	--3043
		x"0b",	--3044
		x"09",	--3045
		x"ea",	--3046
		x"0b",	--3047
		x"0a",	--3048
		x"09",	--3049
		x"08",	--3050
		x"07",	--3051
		x"0d",	--3052
		x"1e",	--3053
		x"04",	--3054
		x"1f",	--3055
		x"06",	--3056
		x"5a",	--3057
		x"01",	--3058
		x"6c",	--3059
		x"6c",	--3060
		x"70",	--3061
		x"6c",	--3062
		x"6a",	--3063
		x"6c",	--3064
		x"36",	--3065
		x"0e",	--3066
		x"32",	--3067
		x"1b",	--3068
		x"02",	--3069
		x"3b",	--3070
		x"82",	--3071
		x"6d",	--3072
		x"3b",	--3073
		x"80",	--3074
		x"5e",	--3075
		x"0c",	--3076
		x"0d",	--3077
		x"3c",	--3078
		x"7f",	--3079
		x"0d",	--3080
		x"3c",	--3081
		x"40",	--3082
		x"40",	--3083
		x"3e",	--3084
		x"3f",	--3085
		x"0f",	--3086
		x"0f",	--3087
		x"4a",	--3088
		x"0d",	--3089
		x"3d",	--3090
		x"7f",	--3091
		x"12",	--3092
		x"0f",	--3093
		x"0e",	--3094
		x"12",	--3095
		x"0f",	--3096
		x"0e",	--3097
		x"12",	--3098
		x"0f",	--3099
		x"0e",	--3100
		x"12",	--3101
		x"0f",	--3102
		x"0e",	--3103
		x"12",	--3104
		x"0f",	--3105
		x"0e",	--3106
		x"12",	--3107
		x"0f",	--3108
		x"0e",	--3109
		x"12",	--3110
		x"0f",	--3111
		x"0e",	--3112
		x"3e",	--3113
		x"3f",	--3114
		x"7f",	--3115
		x"4d",	--3116
		x"05",	--3117
		x"0f",	--3118
		x"cc",	--3119
		x"4d",	--3120
		x"0e",	--3121
		x"0f",	--3122
		x"4d",	--3123
		x"0d",	--3124
		x"0d",	--3125
		x"0d",	--3126
		x"0d",	--3127
		x"0d",	--3128
		x"0d",	--3129
		x"0d",	--3130
		x"0c",	--3131
		x"3c",	--3132
		x"7f",	--3133
		x"0c",	--3134
		x"4f",	--3135
		x"0f",	--3136
		x"0f",	--3137
		x"0f",	--3138
		x"0d",	--3139
		x"0d",	--3140
		x"0f",	--3141
		x"37",	--3142
		x"38",	--3143
		x"39",	--3144
		x"3a",	--3145
		x"3b",	--3146
		x"30",	--3147
		x"0d",	--3148
		x"be",	--3149
		x"0c",	--3150
		x"0d",	--3151
		x"3c",	--3152
		x"80",	--3153
		x"0d",	--3154
		x"0c",	--3155
		x"02",	--3156
		x"0d",	--3157
		x"b8",	--3158
		x"3e",	--3159
		x"40",	--3160
		x"0f",	--3161
		x"b4",	--3162
		x"12",	--3163
		x"0f",	--3164
		x"0e",	--3165
		x"0d",	--3166
		x"3d",	--3167
		x"80",	--3168
		x"b2",	--3169
		x"7d",	--3170
		x"0e",	--3171
		x"0f",	--3172
		x"cd",	--3173
		x"0e",	--3174
		x"3f",	--3175
		x"10",	--3176
		x"3e",	--3177
		x"3f",	--3178
		x"7f",	--3179
		x"7d",	--3180
		x"c5",	--3181
		x"37",	--3182
		x"82",	--3183
		x"07",	--3184
		x"37",	--3185
		x"1a",	--3186
		x"4f",	--3187
		x"0c",	--3188
		x"0d",	--3189
		x"4b",	--3190
		x"7b",	--3191
		x"1f",	--3192
		x"05",	--3193
		x"12",	--3194
		x"0d",	--3195
		x"0c",	--3196
		x"7b",	--3197
		x"fb",	--3198
		x"18",	--3199
		x"09",	--3200
		x"77",	--3201
		x"1f",	--3202
		x"04",	--3203
		x"08",	--3204
		x"09",	--3205
		x"77",	--3206
		x"fc",	--3207
		x"38",	--3208
		x"39",	--3209
		x"08",	--3210
		x"09",	--3211
		x"1e",	--3212
		x"0f",	--3213
		x"08",	--3214
		x"04",	--3215
		x"09",	--3216
		x"02",	--3217
		x"0e",	--3218
		x"0f",	--3219
		x"08",	--3220
		x"09",	--3221
		x"08",	--3222
		x"09",	--3223
		x"0e",	--3224
		x"0f",	--3225
		x"3e",	--3226
		x"7f",	--3227
		x"0f",	--3228
		x"3e",	--3229
		x"40",	--3230
		x"26",	--3231
		x"38",	--3232
		x"3f",	--3233
		x"09",	--3234
		x"0e",	--3235
		x"0f",	--3236
		x"12",	--3237
		x"0f",	--3238
		x"0e",	--3239
		x"12",	--3240
		x"0f",	--3241
		x"0e",	--3242
		x"12",	--3243
		x"0f",	--3244
		x"0e",	--3245
		x"12",	--3246
		x"0f",	--3247
		x"0e",	--3248
		x"12",	--3249
		x"0f",	--3250
		x"0e",	--3251
		x"12",	--3252
		x"0f",	--3253
		x"0e",	--3254
		x"12",	--3255
		x"0f",	--3256
		x"0e",	--3257
		x"3e",	--3258
		x"3f",	--3259
		x"7f",	--3260
		x"5d",	--3261
		x"39",	--3262
		x"00",	--3263
		x"72",	--3264
		x"4d",	--3265
		x"70",	--3266
		x"08",	--3267
		x"09",	--3268
		x"da",	--3269
		x"0f",	--3270
		x"d8",	--3271
		x"0e",	--3272
		x"0f",	--3273
		x"3e",	--3274
		x"80",	--3275
		x"0f",	--3276
		x"0e",	--3277
		x"04",	--3278
		x"38",	--3279
		x"40",	--3280
		x"09",	--3281
		x"d0",	--3282
		x"0f",	--3283
		x"ce",	--3284
		x"f9",	--3285
		x"0b",	--3286
		x"0a",	--3287
		x"2a",	--3288
		x"5b",	--3289
		x"02",	--3290
		x"3b",	--3291
		x"7f",	--3292
		x"1d",	--3293
		x"02",	--3294
		x"12",	--3295
		x"0d",	--3296
		x"12",	--3297
		x"0d",	--3298
		x"12",	--3299
		x"0d",	--3300
		x"12",	--3301
		x"0d",	--3302
		x"12",	--3303
		x"0d",	--3304
		x"12",	--3305
		x"0d",	--3306
		x"12",	--3307
		x"0d",	--3308
		x"4d",	--3309
		x"5f",	--3310
		x"03",	--3311
		x"3f",	--3312
		x"80",	--3313
		x"0f",	--3314
		x"0f",	--3315
		x"ce",	--3316
		x"01",	--3317
		x"0d",	--3318
		x"2d",	--3319
		x"0a",	--3320
		x"51",	--3321
		x"be",	--3322
		x"82",	--3323
		x"02",	--3324
		x"0c",	--3325
		x"0d",	--3326
		x"0c",	--3327
		x"0d",	--3328
		x"0c",	--3329
		x"0d",	--3330
		x"0c",	--3331
		x"0d",	--3332
		x"0c",	--3333
		x"0d",	--3334
		x"0c",	--3335
		x"0d",	--3336
		x"0c",	--3337
		x"0d",	--3338
		x"0c",	--3339
		x"0d",	--3340
		x"fe",	--3341
		x"03",	--3342
		x"00",	--3343
		x"3d",	--3344
		x"00",	--3345
		x"0b",	--3346
		x"3f",	--3347
		x"81",	--3348
		x"0c",	--3349
		x"0d",	--3350
		x"0a",	--3351
		x"3f",	--3352
		x"3d",	--3353
		x"00",	--3354
		x"f9",	--3355
		x"8e",	--3356
		x"02",	--3357
		x"8e",	--3358
		x"04",	--3359
		x"8e",	--3360
		x"06",	--3361
		x"3a",	--3362
		x"3b",	--3363
		x"30",	--3364
		x"3d",	--3365
		x"ff",	--3366
		x"2a",	--3367
		x"3d",	--3368
		x"81",	--3369
		x"8e",	--3370
		x"02",	--3371
		x"fe",	--3372
		x"03",	--3373
		x"00",	--3374
		x"0c",	--3375
		x"0d",	--3376
		x"0c",	--3377
		x"0d",	--3378
		x"0c",	--3379
		x"0d",	--3380
		x"0c",	--3381
		x"0d",	--3382
		x"0c",	--3383
		x"0d",	--3384
		x"0c",	--3385
		x"0d",	--3386
		x"0c",	--3387
		x"0d",	--3388
		x"0c",	--3389
		x"0d",	--3390
		x"0a",	--3391
		x"0b",	--3392
		x"0a",	--3393
		x"3b",	--3394
		x"00",	--3395
		x"8e",	--3396
		x"04",	--3397
		x"8e",	--3398
		x"06",	--3399
		x"3a",	--3400
		x"3b",	--3401
		x"30",	--3402
		x"0b",	--3403
		x"ad",	--3404
		x"ee",	--3405
		x"00",	--3406
		x"3a",	--3407
		x"3b",	--3408
		x"30",	--3409
		x"0a",	--3410
		x"0c",	--3411
		x"0c",	--3412
		x"0d",	--3413
		x"0c",	--3414
		x"3d",	--3415
		x"10",	--3416
		x"0c",	--3417
		x"02",	--3418
		x"0d",	--3419
		x"08",	--3420
		x"de",	--3421
		x"00",	--3422
		x"e4",	--3423
		x"0b",	--3424
		x"f2",	--3425
		x"ee",	--3426
		x"00",	--3427
		x"e3",	--3428
		x"ce",	--3429
		x"00",	--3430
		x"dc",	--3431
		x"0b",	--3432
		x"6d",	--3433
		x"6d",	--3434
		x"12",	--3435
		x"6c",	--3436
		x"6c",	--3437
		x"0f",	--3438
		x"6d",	--3439
		x"41",	--3440
		x"6c",	--3441
		x"11",	--3442
		x"6d",	--3443
		x"0d",	--3444
		x"6c",	--3445
		x"14",	--3446
		x"5d",	--3447
		x"01",	--3448
		x"5d",	--3449
		x"01",	--3450
		x"14",	--3451
		x"4d",	--3452
		x"09",	--3453
		x"1e",	--3454
		x"0f",	--3455
		x"3b",	--3456
		x"30",	--3457
		x"6c",	--3458
		x"28",	--3459
		x"ce",	--3460
		x"01",	--3461
		x"f7",	--3462
		x"3e",	--3463
		x"0f",	--3464
		x"3b",	--3465
		x"30",	--3466
		x"cf",	--3467
		x"01",	--3468
		x"f0",	--3469
		x"3e",	--3470
		x"f8",	--3471
		x"1b",	--3472
		x"02",	--3473
		x"1c",	--3474
		x"02",	--3475
		x"0c",	--3476
		x"e6",	--3477
		x"0b",	--3478
		x"16",	--3479
		x"1b",	--3480
		x"04",	--3481
		x"1f",	--3482
		x"06",	--3483
		x"1c",	--3484
		x"04",	--3485
		x"1e",	--3486
		x"06",	--3487
		x"0e",	--3488
		x"da",	--3489
		x"0f",	--3490
		x"02",	--3491
		x"0c",	--3492
		x"d6",	--3493
		x"0f",	--3494
		x"06",	--3495
		x"0e",	--3496
		x"02",	--3497
		x"0b",	--3498
		x"02",	--3499
		x"0e",	--3500
		x"d1",	--3501
		x"4d",	--3502
		x"ce",	--3503
		x"3e",	--3504
		x"d6",	--3505
		x"6c",	--3506
		x"d7",	--3507
		x"5e",	--3508
		x"01",	--3509
		x"5f",	--3510
		x"01",	--3511
		x"0e",	--3512
		x"c5",	--3513
		x"1e",	--3514
		x"1a",	--3515
		x"1e",	--3516
		x"0b",	--3517
		x"1d",	--3518
		x"18",	--3519
		x"cd",	--3520
		x"00",	--3521
		x"1d",	--3522
		x"82",	--3523
		x"18",	--3524
		x"3e",	--3525
		x"82",	--3526
		x"1a",	--3527
		x"30",	--3528
		x"3f",	--3529
		x"30",	--3530
		x"0b",	--3531
		x"0a",	--3532
		x"21",	--3533
		x"81",	--3534
		x"00",	--3535
		x"1a",	--3536
		x"18",	--3537
		x"1b",	--3538
		x"1a",	--3539
		x"0d",	--3540
		x"0e",	--3541
		x"3f",	--3542
		x"74",	--3543
		x"b0",	--3544
		x"c8",	--3545
		x"0f",	--3546
		x"05",	--3547
		x"0e",	--3548
		x"0e",	--3549
		x"ce",	--3550
		x"ff",	--3551
		x"04",	--3552
		x"1e",	--3553
		x"18",	--3554
		x"ce",	--3555
		x"00",	--3556
		x"21",	--3557
		x"3a",	--3558
		x"3b",	--3559
		x"30",	--3560
		x"92",	--3561
		x"02",	--3562
		x"18",	--3563
		x"b2",	--3564
		x"ff",	--3565
		x"1a",	--3566
		x"0e",	--3567
		x"3e",	--3568
		x"06",	--3569
		x"1f",	--3570
		x"04",	--3571
		x"b0",	--3572
		x"96",	--3573
		x"30",	--3574
		x"92",	--3575
		x"02",	--3576
		x"18",	--3577
		x"92",	--3578
		x"04",	--3579
		x"1a",	--3580
		x"0e",	--3581
		x"3e",	--3582
		x"1f",	--3583
		x"06",	--3584
		x"b0",	--3585
		x"96",	--3586
		x"30",	--3587
		x"0c",	--3588
		x"82",	--3589
		x"18",	--3590
		x"b2",	--3591
		x"ff",	--3592
		x"1a",	--3593
		x"0e",	--3594
		x"0f",	--3595
		x"b0",	--3596
		x"96",	--3597
		x"30",	--3598
		x"82",	--3599
		x"18",	--3600
		x"82",	--3601
		x"1a",	--3602
		x"0e",	--3603
		x"0f",	--3604
		x"b0",	--3605
		x"96",	--3606
		x"30",	--3607
		x"0b",	--3608
		x"0a",	--3609
		x"09",	--3610
		x"08",	--3611
		x"07",	--3612
		x"06",	--3613
		x"05",	--3614
		x"04",	--3615
		x"31",	--3616
		x"08",	--3617
		x"81",	--3618
		x"04",	--3619
		x"09",	--3620
		x"1f",	--3621
		x"1a",	--3622
		x"1d",	--3623
		x"1c",	--3624
		x"4c",	--3625
		x"04",	--3626
		x"84",	--3627
		x"45",	--3628
		x"4e",	--3629
		x"7e",	--3630
		x"40",	--3631
		x"11",	--3632
		x"f1",	--3633
		x"30",	--3634
		x"00",	--3635
		x"0e",	--3636
		x"8e",	--3637
		x"5e",	--3638
		x"03",	--3639
		x"7e",	--3640
		x"58",	--3641
		x"02",	--3642
		x"7e",	--3643
		x"78",	--3644
		x"c1",	--3645
		x"01",	--3646
		x"0c",	--3647
		x"2c",	--3648
		x"0f",	--3649
		x"7e",	--3650
		x"20",	--3651
		x"04",	--3652
		x"f1",	--3653
		x"30",	--3654
		x"00",	--3655
		x"04",	--3656
		x"4c",	--3657
		x"05",	--3658
		x"c1",	--3659
		x"00",	--3660
		x"0c",	--3661
		x"1c",	--3662
		x"01",	--3663
		x"0c",	--3664
		x"0a",	--3665
		x"8c",	--3666
		x"8c",	--3667
		x"8c",	--3668
		x"8c",	--3669
		x"0b",	--3670
		x"06",	--3671
		x"0c",	--3672
		x"8c",	--3673
		x"8c",	--3674
		x"8c",	--3675
		x"8c",	--3676
		x"07",	--3677
		x"0a",	--3678
		x"0b",	--3679
		x"0e",	--3680
		x"8e",	--3681
		x"c1",	--3682
		x"02",	--3683
		x"6e",	--3684
		x"02",	--3685
		x"07",	--3686
		x"01",	--3687
		x"37",	--3688
		x"4f",	--3689
		x"7f",	--3690
		x"10",	--3691
		x"3c",	--3692
		x"1d",	--3693
		x"04",	--3694
		x"3d",	--3695
		x"1d",	--3696
		x"cd",	--3697
		x"00",	--3698
		x"fc",	--3699
		x"1d",	--3700
		x"04",	--3701
		x"09",	--3702
		x"02",	--3703
		x"09",	--3704
		x"01",	--3705
		x"09",	--3706
		x"e1",	--3707
		x"02",	--3708
		x"05",	--3709
		x"09",	--3710
		x"02",	--3711
		x"09",	--3712
		x"01",	--3713
		x"09",	--3714
		x"05",	--3715
		x"07",	--3716
		x"01",	--3717
		x"05",	--3718
		x"4f",	--3719
		x"0d",	--3720
		x"f1",	--3721
		x"20",	--3722
		x"06",	--3723
		x"06",	--3724
		x"0b",	--3725
		x"0e",	--3726
		x"0f",	--3727
		x"0f",	--3728
		x"6f",	--3729
		x"8f",	--3730
		x"16",	--3731
		x"88",	--3732
		x"01",	--3733
		x"06",	--3734
		x"06",	--3735
		x"f6",	--3736
		x"0b",	--3737
		x"f1",	--3738
		x"30",	--3739
		x"06",	--3740
		x"05",	--3741
		x"05",	--3742
		x"5f",	--3743
		x"06",	--3744
		x"8f",	--3745
		x"88",	--3746
		x"1b",	--3747
		x"0f",	--3748
		x"0f",	--3749
		x"0f",	--3750
		x"f7",	--3751
		x"0a",	--3752
		x"06",	--3753
		x"0b",	--3754
		x"07",	--3755
		x"1b",	--3756
		x"0f",	--3757
		x"0f",	--3758
		x"6f",	--3759
		x"8f",	--3760
		x"16",	--3761
		x"88",	--3762
		x"06",	--3763
		x"f7",	--3764
		x"e1",	--3765
		x"02",	--3766
		x"02",	--3767
		x"4a",	--3768
		x"08",	--3769
		x"1a",	--3770
		x"04",	--3771
		x"0a",	--3772
		x"0d",	--3773
		x"3f",	--3774
		x"30",	--3775
		x"88",	--3776
		x"7a",	--3777
		x"4a",	--3778
		x"fa",	--3779
		x"44",	--3780
		x"0b",	--3781
		x"f3",	--3782
		x"37",	--3783
		x"8f",	--3784
		x"88",	--3785
		x"1b",	--3786
		x"0f",	--3787
		x"0f",	--3788
		x"6f",	--3789
		x"4f",	--3790
		x"07",	--3791
		x"07",	--3792
		x"f5",	--3793
		x"04",	--3794
		x"3f",	--3795
		x"20",	--3796
		x"88",	--3797
		x"1b",	--3798
		x"0b",	--3799
		x"fa",	--3800
		x"0f",	--3801
		x"31",	--3802
		x"34",	--3803
		x"35",	--3804
		x"36",	--3805
		x"37",	--3806
		x"38",	--3807
		x"39",	--3808
		x"3a",	--3809
		x"3b",	--3810
		x"30",	--3811
		x"0b",	--3812
		x"0a",	--3813
		x"09",	--3814
		x"08",	--3815
		x"07",	--3816
		x"06",	--3817
		x"05",	--3818
		x"04",	--3819
		x"31",	--3820
		x"b6",	--3821
		x"81",	--3822
		x"3a",	--3823
		x"06",	--3824
		x"05",	--3825
		x"81",	--3826
		x"3e",	--3827
		x"c1",	--3828
		x"2f",	--3829
		x"c1",	--3830
		x"2b",	--3831
		x"c1",	--3832
		x"2e",	--3833
		x"c1",	--3834
		x"2a",	--3835
		x"81",	--3836
		x"30",	--3837
		x"81",	--3838
		x"26",	--3839
		x"07",	--3840
		x"81",	--3841
		x"2c",	--3842
		x"0e",	--3843
		x"3e",	--3844
		x"1c",	--3845
		x"81",	--3846
		x"1c",	--3847
		x"30",	--3848
		x"42",	--3849
		x"0f",	--3850
		x"1f",	--3851
		x"81",	--3852
		x"40",	--3853
		x"07",	--3854
		x"1e",	--3855
		x"7e",	--3856
		x"25",	--3857
		x"13",	--3858
		x"81",	--3859
		x"00",	--3860
		x"81",	--3861
		x"02",	--3862
		x"81",	--3863
		x"3e",	--3864
		x"c1",	--3865
		x"2f",	--3866
		x"c1",	--3867
		x"2b",	--3868
		x"c1",	--3869
		x"2e",	--3870
		x"c1",	--3871
		x"2a",	--3872
		x"81",	--3873
		x"30",	--3874
		x"30",	--3875
		x"38",	--3876
		x"05",	--3877
		x"8e",	--3878
		x"0f",	--3879
		x"91",	--3880
		x"3c",	--3881
		x"91",	--3882
		x"2c",	--3883
		x"30",	--3884
		x"1e",	--3885
		x"7e",	--3886
		x"63",	--3887
		x"c5",	--3888
		x"7e",	--3889
		x"64",	--3890
		x"27",	--3891
		x"7e",	--3892
		x"30",	--3893
		x"94",	--3894
		x"7e",	--3895
		x"31",	--3896
		x"1a",	--3897
		x"7e",	--3898
		x"2a",	--3899
		x"77",	--3900
		x"7e",	--3901
		x"2b",	--3902
		x"0a",	--3903
		x"7e",	--3904
		x"23",	--3905
		x"42",	--3906
		x"7e",	--3907
		x"25",	--3908
		x"e0",	--3909
		x"7e",	--3910
		x"20",	--3911
		x"32",	--3912
		x"56",	--3913
		x"7e",	--3914
		x"2d",	--3915
		x"49",	--3916
		x"7e",	--3917
		x"2e",	--3918
		x"5b",	--3919
		x"7e",	--3920
		x"2b",	--3921
		x"28",	--3922
		x"47",	--3923
		x"7e",	--3924
		x"3a",	--3925
		x"8c",	--3926
		x"7e",	--3927
		x"58",	--3928
		x"21",	--3929
		x"e9",	--3930
		x"7e",	--3931
		x"6f",	--3932
		x"24",	--3933
		x"7e",	--3934
		x"70",	--3935
		x"0a",	--3936
		x"7e",	--3937
		x"69",	--3938
		x"e3",	--3939
		x"7e",	--3940
		x"6c",	--3941
		x"22",	--3942
		x"7e",	--3943
		x"64",	--3944
		x"11",	--3945
		x"dc",	--3946
		x"7e",	--3947
		x"73",	--3948
		x"98",	--3949
		x"7e",	--3950
		x"74",	--3951
		x"04",	--3952
		x"7e",	--3953
		x"70",	--3954
		x"07",	--3955
		x"b8",	--3956
		x"7e",	--3957
		x"75",	--3958
		x"d1",	--3959
		x"7e",	--3960
		x"78",	--3961
		x"d2",	--3962
		x"19",	--3963
		x"3e",	--3964
		x"18",	--3965
		x"2c",	--3966
		x"08",	--3967
		x"30",	--3968
		x"0c",	--3969
		x"b1",	--3970
		x"28",	--3971
		x"cb",	--3972
		x"f1",	--3973
		x"00",	--3974
		x"30",	--3975
		x"3c",	--3976
		x"69",	--3977
		x"59",	--3978
		x"6e",	--3979
		x"04",	--3980
		x"7e",	--3981
		x"fe",	--3982
		x"6e",	--3983
		x"01",	--3984
		x"5e",	--3985
		x"c1",	--3986
		x"00",	--3987
		x"30",	--3988
		x"3c",	--3989
		x"f1",	--3990
		x"10",	--3991
		x"00",	--3992
		x"30",	--3993
		x"3c",	--3994
		x"f1",	--3995
		x"2b",	--3996
		x"02",	--3997
		x"30",	--3998
		x"3c",	--3999
		x"f1",	--4000
		x"2b",	--4001
		x"02",	--4002
		x"02",	--4003
		x"30",	--4004
		x"3c",	--4005
		x"f1",	--4006
		x"20",	--4007
		x"02",	--4008
		x"30",	--4009
		x"3c",	--4010
		x"c1",	--4011
		x"2a",	--4012
		x"02",	--4013
		x"30",	--4014
		x"22",	--4015
		x"d1",	--4016
		x"2e",	--4017
		x"30",	--4018
		x"3c",	--4019
		x"0e",	--4020
		x"2e",	--4021
		x"2a",	--4022
		x"0a",	--4023
		x"03",	--4024
		x"81",	--4025
		x"26",	--4026
		x"0d",	--4027
		x"c1",	--4028
		x"2e",	--4029
		x"02",	--4030
		x"30",	--4031
		x"32",	--4032
		x"f1",	--4033
		x"10",	--4034
		x"00",	--4035
		x"3a",	--4036
		x"81",	--4037
		x"26",	--4038
		x"91",	--4039
		x"26",	--4040
		x"05",	--4041
		x"27",	--4042
		x"81",	--4043
		x"26",	--4044
		x"15",	--4045
		x"c1",	--4046
		x"2e",	--4047
		x"12",	--4048
		x"69",	--4049
		x"79",	--4050
		x"10",	--4051
		x"5e",	--4052
		x"01",	--4053
		x"4e",	--4054
		x"4e",	--4055
		x"0e",	--4056
		x"0e",	--4057
		x"4e",	--4058
		x"6a",	--4059
		x"7a",	--4060
		x"7f",	--4061
		x"4a",	--4062
		x"c1",	--4063
		x"00",	--4064
		x"30",	--4065
		x"3c",	--4066
		x"1a",	--4067
		x"26",	--4068
		x"0a",	--4069
		x"0c",	--4070
		x"0c",	--4071
		x"0c",	--4072
		x"0a",	--4073
		x"81",	--4074
		x"26",	--4075
		x"b1",	--4076
		x"d0",	--4077
		x"26",	--4078
		x"8e",	--4079
		x"81",	--4080
		x"26",	--4081
		x"d1",	--4082
		x"2a",	--4083
		x"30",	--4084
		x"3c",	--4085
		x"07",	--4086
		x"27",	--4087
		x"6e",	--4088
		x"c1",	--4089
		x"2e",	--4090
		x"03",	--4091
		x"c1",	--4092
		x"2a",	--4093
		x"26",	--4094
		x"c1",	--4095
		x"04",	--4096
		x"c1",	--4097
		x"05",	--4098
		x"0e",	--4099
		x"2e",	--4100
		x"03",	--4101
		x"07",	--4102
		x"27",	--4103
		x"2e",	--4104
		x"c1",	--4105
		x"2e",	--4106
		x"07",	--4107
		x"e1",	--4108
		x"01",	--4109
		x"1f",	--4110
		x"26",	--4111
		x"c1",	--4112
		x"03",	--4113
		x"06",	--4114
		x"c1",	--4115
		x"2a",	--4116
		x"03",	--4117
		x"91",	--4118
		x"26",	--4119
		x"30",	--4120
		x"0e",	--4121
		x"02",	--4122
		x"3e",	--4123
		x"d8",	--4124
		x"11",	--4125
		x"04",	--4126
		x"11",	--4127
		x"04",	--4128
		x"1d",	--4129
		x"34",	--4130
		x"1f",	--4131
		x"3e",	--4132
		x"b0",	--4133
		x"30",	--4134
		x"21",	--4135
		x"81",	--4136
		x"2c",	--4137
		x"05",	--4138
		x"30",	--4139
		x"1e",	--4140
		x"07",	--4141
		x"27",	--4142
		x"29",	--4143
		x"81",	--4144
		x"1e",	--4145
		x"5e",	--4146
		x"09",	--4147
		x"01",	--4148
		x"4e",	--4149
		x"4e",	--4150
		x"4e",	--4151
		x"4e",	--4152
		x"6a",	--4153
		x"7a",	--4154
		x"f7",	--4155
		x"4a",	--4156
		x"c1",	--4157
		x"00",	--4158
		x"05",	--4159
		x"b1",	--4160
		x"10",	--4161
		x"28",	--4162
		x"53",	--4163
		x"d1",	--4164
		x"01",	--4165
		x"06",	--4166
		x"e1",	--4167
		x"00",	--4168
		x"b1",	--4169
		x"0a",	--4170
		x"28",	--4171
		x"03",	--4172
		x"b1",	--4173
		x"10",	--4174
		x"28",	--4175
		x"6b",	--4176
		x"6b",	--4177
		x"24",	--4178
		x"0c",	--4179
		x"3c",	--4180
		x"28",	--4181
		x"17",	--4182
		x"02",	--4183
		x"16",	--4184
		x"04",	--4185
		x"1b",	--4186
		x"06",	--4187
		x"81",	--4188
		x"1e",	--4189
		x"81",	--4190
		x"20",	--4191
		x"81",	--4192
		x"22",	--4193
		x"81",	--4194
		x"24",	--4195
		x"d1",	--4196
		x"2b",	--4197
		x"08",	--4198
		x"06",	--4199
		x"07",	--4200
		x"04",	--4201
		x"06",	--4202
		x"02",	--4203
		x"0b",	--4204
		x"02",	--4205
		x"c1",	--4206
		x"2b",	--4207
		x"0b",	--4208
		x"0b",	--4209
		x"0b",	--4210
		x"c1",	--4211
		x"2f",	--4212
		x"05",	--4213
		x"20",	--4214
		x"5b",	--4215
		x"07",	--4216
		x"0d",	--4217
		x"27",	--4218
		x"28",	--4219
		x"1b",	--4220
		x"02",	--4221
		x"81",	--4222
		x"1e",	--4223
		x"81",	--4224
		x"20",	--4225
		x"d1",	--4226
		x"2b",	--4227
		x"08",	--4228
		x"09",	--4229
		x"06",	--4230
		x"27",	--4231
		x"2b",	--4232
		x"81",	--4233
		x"1e",	--4234
		x"d1",	--4235
		x"2b",	--4236
		x"0b",	--4237
		x"02",	--4238
		x"c1",	--4239
		x"2b",	--4240
		x"0b",	--4241
		x"0b",	--4242
		x"0b",	--4243
		x"c1",	--4244
		x"2f",	--4245
		x"05",	--4246
		x"f1",	--4247
		x"00",	--4248
		x"12",	--4249
		x"c1",	--4250
		x"2b",	--4251
		x"0f",	--4252
		x"68",	--4253
		x"b1",	--4254
		x"10",	--4255
		x"28",	--4256
		x"03",	--4257
		x"78",	--4258
		x"40",	--4259
		x"05",	--4260
		x"b1",	--4261
		x"28",	--4262
		x"04",	--4263
		x"78",	--4264
		x"20",	--4265
		x"c1",	--4266
		x"00",	--4267
		x"68",	--4268
		x"68",	--4269
		x"30",	--4270
		x"c1",	--4271
		x"2f",	--4272
		x"2d",	--4273
		x"f1",	--4274
		x"2d",	--4275
		x"02",	--4276
		x"68",	--4277
		x"11",	--4278
		x"b1",	--4279
		x"1e",	--4280
		x"b1",	--4281
		x"20",	--4282
		x"b1",	--4283
		x"22",	--4284
		x"b1",	--4285
		x"24",	--4286
		x"91",	--4287
		x"1e",	--4288
		x"81",	--4289
		x"20",	--4290
		x"81",	--4291
		x"22",	--4292
		x"81",	--4293
		x"24",	--4294
		x"17",	--4295
		x"58",	--4296
		x"0f",	--4297
		x"1a",	--4298
		x"1e",	--4299
		x"1b",	--4300
		x"20",	--4301
		x"3a",	--4302
		x"3b",	--4303
		x"0e",	--4304
		x"0f",	--4305
		x"1e",	--4306
		x"0f",	--4307
		x"81",	--4308
		x"1e",	--4309
		x"81",	--4310
		x"20",	--4311
		x"06",	--4312
		x"1a",	--4313
		x"1e",	--4314
		x"3a",	--4315
		x"1a",	--4316
		x"81",	--4317
		x"1e",	--4318
		x"c1",	--4319
		x"1b",	--4320
		x"68",	--4321
		x"6a",	--4322
		x"16",	--4323
		x"1e",	--4324
		x"91",	--4325
		x"20",	--4326
		x"3c",	--4327
		x"18",	--4328
		x"22",	--4329
		x"14",	--4330
		x"24",	--4331
		x"07",	--4332
		x"37",	--4333
		x"1a",	--4334
		x"09",	--4335
		x"91",	--4336
		x"28",	--4337
		x"32",	--4338
		x"1b",	--4339
		x"28",	--4340
		x"8b",	--4341
		x"8b",	--4342
		x"8b",	--4343
		x"8b",	--4344
		x"81",	--4345
		x"34",	--4346
		x"81",	--4347
		x"36",	--4348
		x"81",	--4349
		x"38",	--4350
		x"11",	--4351
		x"3a",	--4352
		x"11",	--4353
		x"3a",	--4354
		x"11",	--4355
		x"3a",	--4356
		x"11",	--4357
		x"3a",	--4358
		x"0c",	--4359
		x"1d",	--4360
		x"44",	--4361
		x"0e",	--4362
		x"0f",	--4363
		x"b0",	--4364
		x"d2",	--4365
		x"31",	--4366
		x"0b",	--4367
		x"3c",	--4368
		x"0a",	--4369
		x"05",	--4370
		x"7b",	--4371
		x"30",	--4372
		x"c7",	--4373
		x"00",	--4374
		x"0c",	--4375
		x"4b",	--4376
		x"d1",	--4377
		x"01",	--4378
		x"03",	--4379
		x"7a",	--4380
		x"37",	--4381
		x"02",	--4382
		x"7a",	--4383
		x"57",	--4384
		x"4a",	--4385
		x"c7",	--4386
		x"00",	--4387
		x"06",	--4388
		x"36",	--4389
		x"11",	--4390
		x"3a",	--4391
		x"11",	--4392
		x"3a",	--4393
		x"11",	--4394
		x"3a",	--4395
		x"11",	--4396
		x"3a",	--4397
		x"0c",	--4398
		x"1d",	--4399
		x"44",	--4400
		x"0e",	--4401
		x"0f",	--4402
		x"b0",	--4403
		x"ac",	--4404
		x"31",	--4405
		x"09",	--4406
		x"81",	--4407
		x"3c",	--4408
		x"08",	--4409
		x"04",	--4410
		x"37",	--4411
		x"0c",	--4412
		x"b2",	--4413
		x"0d",	--4414
		x"b0",	--4415
		x"0e",	--4416
		x"ae",	--4417
		x"0f",	--4418
		x"ac",	--4419
		x"81",	--4420
		x"1e",	--4421
		x"81",	--4422
		x"20",	--4423
		x"81",	--4424
		x"22",	--4425
		x"81",	--4426
		x"24",	--4427
		x"6c",	--4428
		x"58",	--4429
		x"3e",	--4430
		x"14",	--4431
		x"1e",	--4432
		x"17",	--4433
		x"20",	--4434
		x"08",	--4435
		x"38",	--4436
		x"1a",	--4437
		x"19",	--4438
		x"28",	--4439
		x"89",	--4440
		x"89",	--4441
		x"89",	--4442
		x"89",	--4443
		x"1c",	--4444
		x"28",	--4445
		x"0d",	--4446
		x"0e",	--4447
		x"0f",	--4448
		x"b0",	--4449
		x"d6",	--4450
		x"0b",	--4451
		x"3e",	--4452
		x"0a",	--4453
		x"05",	--4454
		x"7b",	--4455
		x"30",	--4456
		x"c8",	--4457
		x"00",	--4458
		x"0c",	--4459
		x"4b",	--4460
		x"d1",	--4461
		x"01",	--4462
		x"03",	--4463
		x"7a",	--4464
		x"37",	--4465
		x"02",	--4466
		x"7a",	--4467
		x"57",	--4468
		x"4a",	--4469
		x"c8",	--4470
		x"00",	--4471
		x"06",	--4472
		x"36",	--4473
		x"1c",	--4474
		x"28",	--4475
		x"0d",	--4476
		x"0e",	--4477
		x"0f",	--4478
		x"b0",	--4479
		x"a0",	--4480
		x"04",	--4481
		x"07",	--4482
		x"38",	--4483
		x"0e",	--4484
		x"d0",	--4485
		x"0f",	--4486
		x"ce",	--4487
		x"81",	--4488
		x"1e",	--4489
		x"81",	--4490
		x"20",	--4491
		x"2c",	--4492
		x"17",	--4493
		x"1e",	--4494
		x"08",	--4495
		x"38",	--4496
		x"1a",	--4497
		x"1e",	--4498
		x"28",	--4499
		x"0f",	--4500
		x"b0",	--4501
		x"46",	--4502
		x"0d",	--4503
		x"3f",	--4504
		x"0a",	--4505
		x"05",	--4506
		x"7d",	--4507
		x"30",	--4508
		x"c8",	--4509
		x"00",	--4510
		x"0c",	--4511
		x"4d",	--4512
		x"d1",	--4513
		x"01",	--4514
		x"03",	--4515
		x"7c",	--4516
		x"37",	--4517
		x"02",	--4518
		x"7c",	--4519
		x"57",	--4520
		x"4c",	--4521
		x"c8",	--4522
		x"00",	--4523
		x"06",	--4524
		x"36",	--4525
		x"1e",	--4526
		x"28",	--4527
		x"0f",	--4528
		x"b0",	--4529
		x"2c",	--4530
		x"07",	--4531
		x"38",	--4532
		x"0f",	--4533
		x"db",	--4534
		x"81",	--4535
		x"1e",	--4536
		x"b1",	--4537
		x"0a",	--4538
		x"28",	--4539
		x"02",	--4540
		x"c1",	--4541
		x"02",	--4542
		x"c1",	--4543
		x"2e",	--4544
		x"2a",	--4545
		x"0f",	--4546
		x"3f",	--4547
		x"1c",	--4548
		x"81",	--4549
		x"42",	--4550
		x"1a",	--4551
		x"1c",	--4552
		x"8a",	--4553
		x"8a",	--4554
		x"8a",	--4555
		x"8a",	--4556
		x"81",	--4557
		x"44",	--4558
		x"81",	--4559
		x"46",	--4560
		x"0a",	--4561
		x"8a",	--4562
		x"8a",	--4563
		x"8a",	--4564
		x"8a",	--4565
		x"81",	--4566
		x"48",	--4567
		x"1c",	--4568
		x"42",	--4569
		x"1d",	--4570
		x"44",	--4571
		x"1c",	--4572
		x"46",	--4573
		x"1d",	--4574
		x"48",	--4575
		x"2c",	--4576
		x"1c",	--4577
		x"26",	--4578
		x"0e",	--4579
		x"e1",	--4580
		x"01",	--4581
		x"5e",	--4582
		x"26",	--4583
		x"4e",	--4584
		x"c1",	--4585
		x"03",	--4586
		x"06",	--4587
		x"c1",	--4588
		x"2a",	--4589
		x"03",	--4590
		x"91",	--4591
		x"26",	--4592
		x"30",	--4593
		x"11",	--4594
		x"04",	--4595
		x"11",	--4596
		x"04",	--4597
		x"1d",	--4598
		x"34",	--4599
		x"0e",	--4600
		x"1e",	--4601
		x"1f",	--4602
		x"3e",	--4603
		x"b0",	--4604
		x"30",	--4605
		x"21",	--4606
		x"81",	--4607
		x"2c",	--4608
		x"0d",	--4609
		x"7f",	--4610
		x"8f",	--4611
		x"91",	--4612
		x"3c",	--4613
		x"0e",	--4614
		x"0e",	--4615
		x"19",	--4616
		x"40",	--4617
		x"f7",	--4618
		x"81",	--4619
		x"3e",	--4620
		x"81",	--4621
		x"2c",	--4622
		x"07",	--4623
		x"0e",	--4624
		x"91",	--4625
		x"26",	--4626
		x"30",	--4627
		x"d1",	--4628
		x"2e",	--4629
		x"c1",	--4630
		x"2a",	--4631
		x"03",	--4632
		x"05",	--4633
		x"d1",	--4634
		x"2a",	--4635
		x"81",	--4636
		x"26",	--4637
		x"17",	--4638
		x"16",	--4639
		x"40",	--4640
		x"6e",	--4641
		x"4e",	--4642
		x"02",	--4643
		x"30",	--4644
		x"14",	--4645
		x"1f",	--4646
		x"2c",	--4647
		x"31",	--4648
		x"4a",	--4649
		x"34",	--4650
		x"35",	--4651
		x"36",	--4652
		x"37",	--4653
		x"38",	--4654
		x"39",	--4655
		x"3a",	--4656
		x"3b",	--4657
		x"30",	--4658
		x"0d",	--4659
		x"0f",	--4660
		x"04",	--4661
		x"3d",	--4662
		x"03",	--4663
		x"3f",	--4664
		x"1f",	--4665
		x"0e",	--4666
		x"03",	--4667
		x"5d",	--4668
		x"3e",	--4669
		x"1e",	--4670
		x"0d",	--4671
		x"b0",	--4672
		x"2c",	--4673
		x"3d",	--4674
		x"6d",	--4675
		x"02",	--4676
		x"3e",	--4677
		x"1e",	--4678
		x"5d",	--4679
		x"02",	--4680
		x"3f",	--4681
		x"1f",	--4682
		x"30",	--4683
		x"b0",	--4684
		x"66",	--4685
		x"0f",	--4686
		x"30",	--4687
		x"0b",	--4688
		x"0a",	--4689
		x"09",	--4690
		x"79",	--4691
		x"20",	--4692
		x"0a",	--4693
		x"0b",	--4694
		x"0c",	--4695
		x"0d",	--4696
		x"0e",	--4697
		x"0f",	--4698
		x"0c",	--4699
		x"0d",	--4700
		x"0d",	--4701
		x"06",	--4702
		x"02",	--4703
		x"0c",	--4704
		x"03",	--4705
		x"0c",	--4706
		x"0d",	--4707
		x"1e",	--4708
		x"19",	--4709
		x"f2",	--4710
		x"39",	--4711
		x"3a",	--4712
		x"3b",	--4713
		x"30",	--4714
		x"b0",	--4715
		x"a0",	--4716
		x"0e",	--4717
		x"0f",	--4718
		x"30",	--4719
		x"0b",	--4720
		x"0b",	--4721
		x"0f",	--4722
		x"06",	--4723
		x"3b",	--4724
		x"03",	--4725
		x"3e",	--4726
		x"3f",	--4727
		x"1e",	--4728
		x"0f",	--4729
		x"0d",	--4730
		x"05",	--4731
		x"5b",	--4732
		x"3c",	--4733
		x"3d",	--4734
		x"1c",	--4735
		x"0d",	--4736
		x"b0",	--4737
		x"a0",	--4738
		x"6b",	--4739
		x"04",	--4740
		x"3c",	--4741
		x"3d",	--4742
		x"1c",	--4743
		x"0d",	--4744
		x"5b",	--4745
		x"04",	--4746
		x"3e",	--4747
		x"3f",	--4748
		x"1e",	--4749
		x"0f",	--4750
		x"3b",	--4751
		x"30",	--4752
		x"b0",	--4753
		x"e0",	--4754
		x"0e",	--4755
		x"0f",	--4756
		x"30",	--4757
		x"7c",	--4758
		x"10",	--4759
		x"0d",	--4760
		x"0e",	--4761
		x"0f",	--4762
		x"0e",	--4763
		x"0e",	--4764
		x"02",	--4765
		x"0e",	--4766
		x"1f",	--4767
		x"1c",	--4768
		x"f8",	--4769
		x"30",	--4770
		x"b0",	--4771
		x"2c",	--4772
		x"0f",	--4773
		x"30",	--4774
		x"07",	--4775
		x"06",	--4776
		x"05",	--4777
		x"04",	--4778
		x"30",	--4779
		x"40",	--4780
		x"04",	--4781
		x"05",	--4782
		x"06",	--4783
		x"07",	--4784
		x"08",	--4785
		x"09",	--4786
		x"0a",	--4787
		x"0b",	--4788
		x"0c",	--4789
		x"0d",	--4790
		x"0e",	--4791
		x"0f",	--4792
		x"08",	--4793
		x"09",	--4794
		x"0a",	--4795
		x"0b",	--4796
		x"0b",	--4797
		x"0e",	--4798
		x"08",	--4799
		x"0a",	--4800
		x"0b",	--4801
		x"05",	--4802
		x"09",	--4803
		x"08",	--4804
		x"02",	--4805
		x"08",	--4806
		x"05",	--4807
		x"08",	--4808
		x"09",	--4809
		x"0a",	--4810
		x"0b",	--4811
		x"1c",	--4812
		x"91",	--4813
		x"00",	--4814
		x"e5",	--4815
		x"21",	--4816
		x"34",	--4817
		x"35",	--4818
		x"36",	--4819
		x"37",	--4820
		x"30",	--4821
		x"0b",	--4822
		x"0a",	--4823
		x"09",	--4824
		x"08",	--4825
		x"18",	--4826
		x"0a",	--4827
		x"19",	--4828
		x"0c",	--4829
		x"1a",	--4830
		x"0e",	--4831
		x"1b",	--4832
		x"10",	--4833
		x"b0",	--4834
		x"4e",	--4835
		x"38",	--4836
		x"39",	--4837
		x"3a",	--4838
		x"3b",	--4839
		x"30",	--4840
		x"0b",	--4841
		x"0a",	--4842
		x"09",	--4843
		x"08",	--4844
		x"18",	--4845
		x"0a",	--4846
		x"19",	--4847
		x"0c",	--4848
		x"1a",	--4849
		x"0e",	--4850
		x"1b",	--4851
		x"10",	--4852
		x"b0",	--4853
		x"4e",	--4854
		x"0c",	--4855
		x"0d",	--4856
		x"0e",	--4857
		x"0f",	--4858
		x"38",	--4859
		x"39",	--4860
		x"3a",	--4861
		x"3b",	--4862
		x"30",	--4863
		x"0b",	--4864
		x"0a",	--4865
		x"09",	--4866
		x"08",	--4867
		x"07",	--4868
		x"18",	--4869
		x"0c",	--4870
		x"19",	--4871
		x"0e",	--4872
		x"1a",	--4873
		x"10",	--4874
		x"1b",	--4875
		x"12",	--4876
		x"b0",	--4877
		x"4e",	--4878
		x"17",	--4879
		x"14",	--4880
		x"87",	--4881
		x"00",	--4882
		x"87",	--4883
		x"02",	--4884
		x"87",	--4885
		x"04",	--4886
		x"87",	--4887
		x"06",	--4888
		x"37",	--4889
		x"38",	--4890
		x"39",	--4891
		x"3a",	--4892
		x"3b",	--4893
		x"30",	--4894
		x"00",	--4895
		x"32",	--4896
		x"f0",	--4897
		x"fd",	--4898
		x"57",	--4899
		x"69",	--4900
		x"69",	--4901
		x"67",	--4902
		x"66",	--4903
		x"72",	--4904
		x"61",	--4905
		x"6e",	--4906
		x"77",	--4907
		x"2e",	--4908
		x"69",	--4909
		x"20",	--4910
		x"69",	--4911
		x"65",	--4912
		x"0a",	--4913
		x"57",	--4914
		x"20",	--4915
		x"68",	--4916
		x"75",	--4917
		x"64",	--4918
		x"6e",	--4919
		x"74",	--4920
		x"73",	--4921
		x"65",	--4922
		x"74",	--4923
		x"61",	--4924
		x"0d",	--4925
		x"00",	--4926
		x"74",	--4927
		x"70",	--4928
		x"0a",	--4929
		x"65",	--4930
		x"72",	--4931
		x"72",	--4932
		x"20",	--4933
		x"69",	--4934
		x"73",	--4935
		x"6e",	--4936
		x"20",	--4937
		x"72",	--4938
		x"75",	--4939
		x"65",	--4940
		x"74",	--4941
		x"0a",	--4942
		x"63",	--4943
		x"72",	--4944
		x"65",	--4945
		x"74",	--4946
		x"75",	--4947
		x"61",	--4948
		x"65",	--4949
		x"0d",	--4950
		x"00",	--4951
		x"25",	--4952
		x"20",	--4953
		x"45",	--4954
		x"54",	--4955
		x"52",	--4956
		x"47",	--4957
		x"54",	--4958
		x"3c",	--4959
		x"49",	--4960
		x"45",	--4961
		x"55",	--4962
		x"3e",	--4963
		x"0a",	--4964
		x"25",	--4965
		x"20",	--4966
		x"64",	--4967
		x"0a",	--4968
		x"25",	--4969
		x"64",	--4970
		x"25",	--4971
		x"64",	--4972
		x"25",	--4973
		x"0d",	--4974
		x"00",	--4975
		x"64",	--4976
		x"25",	--4977
		x"0d",	--4978
		x"00",	--4979
		x"d6",	--4980
		x"fe",	--4981
		x"04",	--4982
		x"0c",	--4983
		x"14",	--4984
		x"1c",	--4985
		x"ee",	--4986
		x"f6",	--4987
		x"0d",	--4988
		x"3d",	--4989
		x"3d",	--4990
		x"3d",	--4991
		x"20",	--4992
		x"61",	--4993
		x"63",	--4994
		x"6c",	--4995
		x"4d",	--4996
		x"55",	--4997
		x"3d",	--4998
		x"3d",	--4999
		x"3d",	--5000
		x"0d",	--5001
		x"00",	--5002
		x"6e",	--5003
		x"65",	--5004
		x"61",	--5005
		x"74",	--5006
		x"76",	--5007
		x"20",	--5008
		x"6f",	--5009
		x"65",	--5010
		x"77",	--5011
		x"69",	--5012
		x"65",	--5013
		x"72",	--5014
		x"61",	--5015
		x"00",	--5016
		x"77",	--5017
		x"00",	--5018
		x"6e",	--5019
		x"6f",	--5020
		x"65",	--5021
		x"00",	--5022
		x"70",	--5023
		x"65",	--5024
		x"20",	--5025
		x"6f",	--5026
		x"74",	--5027
		x"6f",	--5028
		x"6c",	--5029
		x"72",	--5030
		x"73",	--5031
		x"65",	--5032
		x"64",	--5033
		x"63",	--5034
		x"6e",	--5035
		x"69",	--5036
		x"75",	--5037
		x"61",	--5038
		x"69",	--5039
		x"6e",	--5040
		x"62",	--5041
		x"6f",	--5042
		x"6c",	--5043
		x"61",	--5044
		x"65",	--5045
		x"00",	--5046
		x"0a",	--5047
		x"08",	--5048
		x"08",	--5049
		x"25",	--5050
		x"00",	--5051
		x"77",	--5052
		x"69",	--5053
		x"65",	--5054
		x"0d",	--5055
		x"65",	--5056
		x"72",	--5057
		x"72",	--5058
		x"20",	--5059
		x"69",	--5060
		x"73",	--5061
		x"6e",	--5062
		x"20",	--5063
		x"72",	--5064
		x"75",	--5065
		x"65",	--5066
		x"74",	--5067
		x"0a",	--5068
		x"63",	--5069
		x"72",	--5070
		x"65",	--5071
		x"74",	--5072
		x"75",	--5073
		x"61",	--5074
		x"65",	--5075
		x"0d",	--5076
		x"00",	--5077
		x"25",	--5078
		x"20",	--5079
		x"45",	--5080
		x"49",	--5081
		x"54",	--5082
		x"52",	--5083
		x"56",	--5084
		x"4c",	--5085
		x"45",	--5086
		x"0a",	--5087
		x"72",	--5088
		x"25",	--5089
		x"20",	--5090
		x"3d",	--5091
		x"64",	--5092
		x"0a",	--5093
		x"09",	--5094
		x"73",	--5095
		x"52",	--5096
		x"47",	--5097
		x"53",	--5098
		x"45",	--5099
		x"0d",	--5100
		x"00",	--5101
		x"65",	--5102
		x"64",	--5103
		x"0d",	--5104
		x"25",	--5105
		x"20",	--5106
		x"73",	--5107
		x"6e",	--5108
		x"74",	--5109
		x"61",	--5110
		x"6e",	--5111
		x"6d",	--5112
		x"65",	--5113
		x"0d",	--5114
		x"00",	--5115
		x"63",	--5116
		x"25",	--5117
		x"0d",	--5118
		x"00",	--5119
		x"63",	--5120
		x"20",	--5121
		x"6f",	--5122
		x"73",	--5123
		x"63",	--5124
		x"20",	--5125
		x"6f",	--5126
		x"6d",	--5127
		x"6e",	--5128
		x"0d",	--5129
		x"00",	--5130
		x"f4",	--5131
		x"22",	--5132
		x"22",	--5133
		x"22",	--5134
		x"22",	--5135
		x"22",	--5136
		x"22",	--5137
		x"22",	--5138
		x"22",	--5139
		x"22",	--5140
		x"22",	--5141
		x"22",	--5142
		x"22",	--5143
		x"22",	--5144
		x"22",	--5145
		x"22",	--5146
		x"22",	--5147
		x"22",	--5148
		x"22",	--5149
		x"22",	--5150
		x"22",	--5151
		x"22",	--5152
		x"22",	--5153
		x"22",	--5154
		x"22",	--5155
		x"22",	--5156
		x"22",	--5157
		x"22",	--5158
		x"22",	--5159
		x"e6",	--5160
		x"22",	--5161
		x"22",	--5162
		x"22",	--5163
		x"22",	--5164
		x"22",	--5165
		x"22",	--5166
		x"22",	--5167
		x"22",	--5168
		x"22",	--5169
		x"22",	--5170
		x"22",	--5171
		x"22",	--5172
		x"22",	--5173
		x"22",	--5174
		x"22",	--5175
		x"22",	--5176
		x"22",	--5177
		x"22",	--5178
		x"22",	--5179
		x"22",	--5180
		x"22",	--5181
		x"22",	--5182
		x"22",	--5183
		x"22",	--5184
		x"22",	--5185
		x"22",	--5186
		x"22",	--5187
		x"22",	--5188
		x"22",	--5189
		x"22",	--5190
		x"22",	--5191
		x"d8",	--5192
		x"ca",	--5193
		x"bc",	--5194
		x"22",	--5195
		x"22",	--5196
		x"22",	--5197
		x"22",	--5198
		x"22",	--5199
		x"22",	--5200
		x"22",	--5201
		x"a4",	--5202
		x"22",	--5203
		x"92",	--5204
		x"22",	--5205
		x"22",	--5206
		x"22",	--5207
		x"22",	--5208
		x"76",	--5209
		x"22",	--5210
		x"22",	--5211
		x"22",	--5212
		x"68",	--5213
		x"56",	--5214
		x"30",	--5215
		x"32",	--5216
		x"34",	--5217
		x"36",	--5218
		x"38",	--5219
		x"61",	--5220
		x"63",	--5221
		x"65",	--5222
		x"00",	--5223
		x"00",	--5224
		x"00",	--5225
		x"00",	--5226
		x"00",	--5227
		x"00",	--5228
		x"02",	--5229
		x"03",	--5230
		x"03",	--5231
		x"04",	--5232
		x"04",	--5233
		x"04",	--5234
		x"04",	--5235
		x"05",	--5236
		x"05",	--5237
		x"05",	--5238
		x"05",	--5239
		x"05",	--5240
		x"05",	--5241
		x"05",	--5242
		x"05",	--5243
		x"06",	--5244
		x"06",	--5245
		x"06",	--5246
		x"06",	--5247
		x"06",	--5248
		x"06",	--5249
		x"06",	--5250
		x"06",	--5251
		x"06",	--5252
		x"06",	--5253
		x"06",	--5254
		x"06",	--5255
		x"06",	--5256
		x"06",	--5257
		x"06",	--5258
		x"06",	--5259
		x"07",	--5260
		x"07",	--5261
		x"07",	--5262
		x"07",	--5263
		x"07",	--5264
		x"07",	--5265
		x"07",	--5266
		x"07",	--5267
		x"07",	--5268
		x"07",	--5269
		x"07",	--5270
		x"07",	--5271
		x"07",	--5272
		x"07",	--5273
		x"07",	--5274
		x"07",	--5275
		x"07",	--5276
		x"07",	--5277
		x"07",	--5278
		x"07",	--5279
		x"07",	--5280
		x"07",	--5281
		x"07",	--5282
		x"07",	--5283
		x"07",	--5284
		x"07",	--5285
		x"07",	--5286
		x"07",	--5287
		x"07",	--5288
		x"07",	--5289
		x"07",	--5290
		x"07",	--5291
		x"08",	--5292
		x"08",	--5293
		x"08",	--5294
		x"08",	--5295
		x"08",	--5296
		x"08",	--5297
		x"08",	--5298
		x"08",	--5299
		x"08",	--5300
		x"08",	--5301
		x"08",	--5302
		x"08",	--5303
		x"08",	--5304
		x"08",	--5305
		x"08",	--5306
		x"08",	--5307
		x"08",	--5308
		x"08",	--5309
		x"08",	--5310
		x"08",	--5311
		x"08",	--5312
		x"08",	--5313
		x"08",	--5314
		x"08",	--5315
		x"08",	--5316
		x"08",	--5317
		x"08",	--5318
		x"08",	--5319
		x"08",	--5320
		x"08",	--5321
		x"08",	--5322
		x"08",	--5323
		x"08",	--5324
		x"08",	--5325
		x"08",	--5326
		x"08",	--5327
		x"08",	--5328
		x"08",	--5329
		x"08",	--5330
		x"08",	--5331
		x"08",	--5332
		x"08",	--5333
		x"08",	--5334
		x"08",	--5335
		x"08",	--5336
		x"08",	--5337
		x"08",	--5338
		x"08",	--5339
		x"08",	--5340
		x"08",	--5341
		x"08",	--5342
		x"08",	--5343
		x"08",	--5344
		x"08",	--5345
		x"08",	--5346
		x"08",	--5347
		x"08",	--5348
		x"08",	--5349
		x"08",	--5350
		x"08",	--5351
		x"08",	--5352
		x"08",	--5353
		x"08",	--5354
		x"08",	--5355
		x"28",	--5356
		x"75",	--5357
		x"6c",	--5358
		x"00",	--5359
		x"ff",	--5360
		x"ff",	--5361
		x"68",	--5362
		x"6c",	--5363
		x"00",	--5364
		x"ff",	--5365
		x"ff",	--5366
		x"ff",	--5367
		x"ff",	--5368
		x"ff",	--5369
		x"ff",	--5370
		x"ff",	--5371
		x"ff",	--5372
		x"ff",	--5373
		x"ff",	--5374
		x"ff",	--5375
		x"ff",	--5376
		x"ff",	--5377
		x"ff",	--5378
		x"ff",	--5379
		x"ff",	--5380
		x"ff",	--5381
		x"ff",	--5382
		x"ff",	--5383
		x"ff",	--5384
		x"ff",	--5385
		x"ff",	--5386
		x"ff",	--5387
		x"ff",	--5388
		x"ff",	--5389
		x"ff",	--5390
		x"ff",	--5391
		x"ff",	--5392
		x"ff",	--5393
		x"ff",	--5394
		x"ff",	--5395
		x"ff",	--5396
		x"ff",	--5397
		x"ff",	--5398
		x"ff",	--5399
		x"ff",	--5400
		x"ff",	--5401
		x"ff",	--5402
		x"ff",	--5403
		x"ff",	--5404
		x"ff",	--5405
		x"ff",	--5406
		x"ff",	--5407
		x"ff",	--5408
		x"ff",	--5409
		x"ff",	--5410
		x"ff",	--5411
		x"ff",	--5412
		x"ff",	--5413
		x"ff",	--5414
		x"ff",	--5415
		x"ff",	--5416
		x"ff",	--5417
		x"ff",	--5418
		x"ff",	--5419
		x"ff",	--5420
		x"ff",	--5421
		x"ff",	--5422
		x"ff",	--5423
		x"ff",	--5424
		x"ff",	--5425
		x"ff",	--5426
		x"ff",	--5427
		x"ff",	--5428
		x"ff",	--5429
		x"ff",	--5430
		x"ff",	--5431
		x"ff",	--5432
		x"ff",	--5433
		x"ff",	--5434
		x"ff",	--5435
		x"ff",	--5436
		x"ff",	--5437
		x"ff",	--5438
		x"ff",	--5439
		x"ff",	--5440
		x"ff",	--5441
		x"ff",	--5442
		x"ff",	--5443
		x"ff",	--5444
		x"ff",	--5445
		x"ff",	--5446
		x"ff",	--5447
		x"ff",	--5448
		x"ff",	--5449
		x"ff",	--5450
		x"ff",	--5451
		x"ff",	--5452
		x"ff",	--5453
		x"ff",	--5454
		x"ff",	--5455
		x"ff",	--5456
		x"ff",	--5457
		x"ff",	--5458
		x"ff",	--5459
		x"ff",	--5460
		x"ff",	--5461
		x"ff",	--5462
		x"ff",	--5463
		x"ff",	--5464
		x"ff",	--5465
		x"ff",	--5466
		x"ff",	--5467
		x"ff",	--5468
		x"ff",	--5469
		x"ff",	--5470
		x"ff",	--5471
		x"ff",	--5472
		x"ff",	--5473
		x"ff",	--5474
		x"ff",	--5475
		x"ff",	--5476
		x"ff",	--5477
		x"ff",	--5478
		x"ff",	--5479
		x"ff",	--5480
		x"ff",	--5481
		x"ff",	--5482
		x"ff",	--5483
		x"ff",	--5484
		x"ff",	--5485
		x"ff",	--5486
		x"ff",	--5487
		x"ff",	--5488
		x"ff",	--5489
		x"ff",	--5490
		x"ff",	--5491
		x"ff",	--5492
		x"ff",	--5493
		x"ff",	--5494
		x"ff",	--5495
		x"ff",	--5496
		x"ff",	--5497
		x"ff",	--5498
		x"ff",	--5499
		x"ff",	--5500
		x"ff",	--5501
		x"ff",	--5502
		x"ff",	--5503
		x"ff",	--5504
		x"ff",	--5505
		x"ff",	--5506
		x"ff",	--5507
		x"ff",	--5508
		x"ff",	--5509
		x"ff",	--5510
		x"ff",	--5511
		x"ff",	--5512
		x"ff",	--5513
		x"ff",	--5514
		x"ff",	--5515
		x"ff",	--5516
		x"ff",	--5517
		x"ff",	--5518
		x"ff",	--5519
		x"ff",	--5520
		x"ff",	--5521
		x"ff",	--5522
		x"ff",	--5523
		x"ff",	--5524
		x"ff",	--5525
		x"ff",	--5526
		x"ff",	--5527
		x"ff",	--5528
		x"ff",	--5529
		x"ff",	--5530
		x"ff",	--5531
		x"ff",	--5532
		x"ff",	--5533
		x"ff",	--5534
		x"ff",	--5535
		x"ff",	--5536
		x"ff",	--5537
		x"ff",	--5538
		x"ff",	--5539
		x"ff",	--5540
		x"ff",	--5541
		x"ff",	--5542
		x"ff",	--5543
		x"ff",	--5544
		x"ff",	--5545
		x"ff",	--5546
		x"ff",	--5547
		x"ff",	--5548
		x"ff",	--5549
		x"ff",	--5550
		x"ff",	--5551
		x"ff",	--5552
		x"ff",	--5553
		x"ff",	--5554
		x"ff",	--5555
		x"ff",	--5556
		x"ff",	--5557
		x"ff",	--5558
		x"ff",	--5559
		x"ff",	--5560
		x"ff",	--5561
		x"ff",	--5562
		x"ff",	--5563
		x"ff",	--5564
		x"ff",	--5565
		x"ff",	--5566
		x"ff",	--5567
		x"ff",	--5568
		x"ff",	--5569
		x"ff",	--5570
		x"ff",	--5571
		x"ff",	--5572
		x"ff",	--5573
		x"ff",	--5574
		x"ff",	--5575
		x"ff",	--5576
		x"ff",	--5577
		x"ff",	--5578
		x"ff",	--5579
		x"ff",	--5580
		x"ff",	--5581
		x"ff",	--5582
		x"ff",	--5583
		x"ff",	--5584
		x"ff",	--5585
		x"ff",	--5586
		x"ff",	--5587
		x"ff",	--5588
		x"ff",	--5589
		x"ff",	--5590
		x"ff",	--5591
		x"ff",	--5592
		x"ff",	--5593
		x"ff",	--5594
		x"ff",	--5595
		x"ff",	--5596
		x"ff",	--5597
		x"ff",	--5598
		x"ff",	--5599
		x"ff",	--5600
		x"ff",	--5601
		x"ff",	--5602
		x"ff",	--5603
		x"ff",	--5604
		x"ff",	--5605
		x"ff",	--5606
		x"ff",	--5607
		x"ff",	--5608
		x"ff",	--5609
		x"ff",	--5610
		x"ff",	--5611
		x"ff",	--5612
		x"ff",	--5613
		x"ff",	--5614
		x"ff",	--5615
		x"ff",	--5616
		x"ff",	--5617
		x"ff",	--5618
		x"ff",	--5619
		x"ff",	--5620
		x"ff",	--5621
		x"ff",	--5622
		x"ff",	--5623
		x"ff",	--5624
		x"ff",	--5625
		x"ff",	--5626
		x"ff",	--5627
		x"ff",	--5628
		x"ff",	--5629
		x"ff",	--5630
		x"ff",	--5631
		x"ff",	--5632
		x"ff",	--5633
		x"ff",	--5634
		x"ff",	--5635
		x"ff",	--5636
		x"ff",	--5637
		x"ff",	--5638
		x"ff",	--5639
		x"ff",	--5640
		x"ff",	--5641
		x"ff",	--5642
		x"ff",	--5643
		x"ff",	--5644
		x"ff",	--5645
		x"ff",	--5646
		x"ff",	--5647
		x"ff",	--5648
		x"ff",	--5649
		x"ff",	--5650
		x"ff",	--5651
		x"ff",	--5652
		x"ff",	--5653
		x"ff",	--5654
		x"ff",	--5655
		x"ff",	--5656
		x"ff",	--5657
		x"ff",	--5658
		x"ff",	--5659
		x"ff",	--5660
		x"ff",	--5661
		x"ff",	--5662
		x"ff",	--5663
		x"ff",	--5664
		x"ff",	--5665
		x"ff",	--5666
		x"ff",	--5667
		x"ff",	--5668
		x"ff",	--5669
		x"ff",	--5670
		x"ff",	--5671
		x"ff",	--5672
		x"ff",	--5673
		x"ff",	--5674
		x"ff",	--5675
		x"ff",	--5676
		x"ff",	--5677
		x"ff",	--5678
		x"ff",	--5679
		x"ff",	--5680
		x"ff",	--5681
		x"ff",	--5682
		x"ff",	--5683
		x"ff",	--5684
		x"ff",	--5685
		x"ff",	--5686
		x"ff",	--5687
		x"ff",	--5688
		x"ff",	--5689
		x"ff",	--5690
		x"ff",	--5691
		x"ff",	--5692
		x"ff",	--5693
		x"ff",	--5694
		x"ff",	--5695
		x"ff",	--5696
		x"ff",	--5697
		x"ff",	--5698
		x"ff",	--5699
		x"ff",	--5700
		x"ff",	--5701
		x"ff",	--5702
		x"ff",	--5703
		x"ff",	--5704
		x"ff",	--5705
		x"ff",	--5706
		x"ff",	--5707
		x"ff",	--5708
		x"ff",	--5709
		x"ff",	--5710
		x"ff",	--5711
		x"ff",	--5712
		x"ff",	--5713
		x"ff",	--5714
		x"ff",	--5715
		x"ff",	--5716
		x"ff",	--5717
		x"ff",	--5718
		x"ff",	--5719
		x"ff",	--5720
		x"ff",	--5721
		x"ff",	--5722
		x"ff",	--5723
		x"ff",	--5724
		x"ff",	--5725
		x"ff",	--5726
		x"ff",	--5727
		x"ff",	--5728
		x"ff",	--5729
		x"ff",	--5730
		x"ff",	--5731
		x"ff",	--5732
		x"ff",	--5733
		x"ff",	--5734
		x"ff",	--5735
		x"ff",	--5736
		x"ff",	--5737
		x"ff",	--5738
		x"ff",	--5739
		x"ff",	--5740
		x"ff",	--5741
		x"ff",	--5742
		x"ff",	--5743
		x"ff",	--5744
		x"ff",	--5745
		x"ff",	--5746
		x"ff",	--5747
		x"ff",	--5748
		x"ff",	--5749
		x"ff",	--5750
		x"ff",	--5751
		x"ff",	--5752
		x"ff",	--5753
		x"ff",	--5754
		x"ff",	--5755
		x"ff",	--5756
		x"ff",	--5757
		x"ff",	--5758
		x"ff",	--5759
		x"ff",	--5760
		x"ff",	--5761
		x"ff",	--5762
		x"ff",	--5763
		x"ff",	--5764
		x"ff",	--5765
		x"ff",	--5766
		x"ff",	--5767
		x"ff",	--5768
		x"ff",	--5769
		x"ff",	--5770
		x"ff",	--5771
		x"ff",	--5772
		x"ff",	--5773
		x"ff",	--5774
		x"ff",	--5775
		x"ff",	--5776
		x"ff",	--5777
		x"ff",	--5778
		x"ff",	--5779
		x"ff",	--5780
		x"ff",	--5781
		x"ff",	--5782
		x"ff",	--5783
		x"ff",	--5784
		x"ff",	--5785
		x"ff",	--5786
		x"ff",	--5787
		x"ff",	--5788
		x"ff",	--5789
		x"ff",	--5790
		x"ff",	--5791
		x"ff",	--5792
		x"ff",	--5793
		x"ff",	--5794
		x"ff",	--5795
		x"ff",	--5796
		x"ff",	--5797
		x"ff",	--5798
		x"ff",	--5799
		x"ff",	--5800
		x"ff",	--5801
		x"ff",	--5802
		x"ff",	--5803
		x"ff",	--5804
		x"ff",	--5805
		x"ff",	--5806
		x"ff",	--5807
		x"ff",	--5808
		x"ff",	--5809
		x"ff",	--5810
		x"ff",	--5811
		x"ff",	--5812
		x"ff",	--5813
		x"ff",	--5814
		x"ff",	--5815
		x"ff",	--5816
		x"ff",	--5817
		x"ff",	--5818
		x"ff",	--5819
		x"ff",	--5820
		x"ff",	--5821
		x"ff",	--5822
		x"ff",	--5823
		x"ff",	--5824
		x"ff",	--5825
		x"ff",	--5826
		x"ff",	--5827
		x"ff",	--5828
		x"ff",	--5829
		x"ff",	--5830
		x"ff",	--5831
		x"ff",	--5832
		x"ff",	--5833
		x"ff",	--5834
		x"ff",	--5835
		x"ff",	--5836
		x"ff",	--5837
		x"ff",	--5838
		x"ff",	--5839
		x"ff",	--5840
		x"ff",	--5841
		x"ff",	--5842
		x"ff",	--5843
		x"ff",	--5844
		x"ff",	--5845
		x"ff",	--5846
		x"ff",	--5847
		x"ff",	--5848
		x"ff",	--5849
		x"ff",	--5850
		x"ff",	--5851
		x"ff",	--5852
		x"ff",	--5853
		x"ff",	--5854
		x"ff",	--5855
		x"ff",	--5856
		x"ff",	--5857
		x"ff",	--5858
		x"ff",	--5859
		x"ff",	--5860
		x"ff",	--5861
		x"ff",	--5862
		x"ff",	--5863
		x"ff",	--5864
		x"ff",	--5865
		x"ff",	--5866
		x"ff",	--5867
		x"ff",	--5868
		x"ff",	--5869
		x"ff",	--5870
		x"ff",	--5871
		x"ff",	--5872
		x"ff",	--5873
		x"ff",	--5874
		x"ff",	--5875
		x"ff",	--5876
		x"ff",	--5877
		x"ff",	--5878
		x"ff",	--5879
		x"ff",	--5880
		x"ff",	--5881
		x"ff",	--5882
		x"ff",	--5883
		x"ff",	--5884
		x"ff",	--5885
		x"ff",	--5886
		x"ff",	--5887
		x"ff",	--5888
		x"ff",	--5889
		x"ff",	--5890
		x"ff",	--5891
		x"ff",	--5892
		x"ff",	--5893
		x"ff",	--5894
		x"ff",	--5895
		x"ff",	--5896
		x"ff",	--5897
		x"ff",	--5898
		x"ff",	--5899
		x"ff",	--5900
		x"ff",	--5901
		x"ff",	--5902
		x"ff",	--5903
		x"ff",	--5904
		x"ff",	--5905
		x"ff",	--5906
		x"ff",	--5907
		x"ff",	--5908
		x"ff",	--5909
		x"ff",	--5910
		x"ff",	--5911
		x"ff",	--5912
		x"ff",	--5913
		x"ff",	--5914
		x"ff",	--5915
		x"ff",	--5916
		x"ff",	--5917
		x"ff",	--5918
		x"ff",	--5919
		x"ff",	--5920
		x"ff",	--5921
		x"ff",	--5922
		x"ff",	--5923
		x"ff",	--5924
		x"ff",	--5925
		x"ff",	--5926
		x"ff",	--5927
		x"ff",	--5928
		x"ff",	--5929
		x"ff",	--5930
		x"ff",	--5931
		x"ff",	--5932
		x"ff",	--5933
		x"ff",	--5934
		x"ff",	--5935
		x"ff",	--5936
		x"ff",	--5937
		x"ff",	--5938
		x"ff",	--5939
		x"ff",	--5940
		x"ff",	--5941
		x"ff",	--5942
		x"ff",	--5943
		x"ff",	--5944
		x"ff",	--5945
		x"ff",	--5946
		x"ff",	--5947
		x"ff",	--5948
		x"ff",	--5949
		x"ff",	--5950
		x"ff",	--5951
		x"ff",	--5952
		x"ff",	--5953
		x"ff",	--5954
		x"ff",	--5955
		x"ff",	--5956
		x"ff",	--5957
		x"ff",	--5958
		x"ff",	--5959
		x"ff",	--5960
		x"ff",	--5961
		x"ff",	--5962
		x"ff",	--5963
		x"ff",	--5964
		x"ff",	--5965
		x"ff",	--5966
		x"ff",	--5967
		x"ff",	--5968
		x"ff",	--5969
		x"ff",	--5970
		x"ff",	--5971
		x"ff",	--5972
		x"ff",	--5973
		x"ff",	--5974
		x"ff",	--5975
		x"ff",	--5976
		x"ff",	--5977
		x"ff",	--5978
		x"ff",	--5979
		x"ff",	--5980
		x"ff",	--5981
		x"ff",	--5982
		x"ff",	--5983
		x"ff",	--5984
		x"ff",	--5985
		x"ff",	--5986
		x"ff",	--5987
		x"ff",	--5988
		x"ff",	--5989
		x"ff",	--5990
		x"ff",	--5991
		x"ff",	--5992
		x"ff",	--5993
		x"ff",	--5994
		x"ff",	--5995
		x"ff",	--5996
		x"ff",	--5997
		x"ff",	--5998
		x"ff",	--5999
		x"ff",	--6000
		x"ff",	--6001
		x"ff",	--6002
		x"ff",	--6003
		x"ff",	--6004
		x"ff",	--6005
		x"ff",	--6006
		x"ff",	--6007
		x"ff",	--6008
		x"ff",	--6009
		x"ff",	--6010
		x"ff",	--6011
		x"ff",	--6012
		x"ff",	--6013
		x"ff",	--6014
		x"ff",	--6015
		x"ff",	--6016
		x"ff",	--6017
		x"ff",	--6018
		x"ff",	--6019
		x"ff",	--6020
		x"ff",	--6021
		x"ff",	--6022
		x"ff",	--6023
		x"ff",	--6024
		x"ff",	--6025
		x"ff",	--6026
		x"ff",	--6027
		x"ff",	--6028
		x"ff",	--6029
		x"ff",	--6030
		x"ff",	--6031
		x"ff",	--6032
		x"ff",	--6033
		x"ff",	--6034
		x"ff",	--6035
		x"ff",	--6036
		x"ff",	--6037
		x"ff",	--6038
		x"ff",	--6039
		x"ff",	--6040
		x"ff",	--6041
		x"ff",	--6042
		x"ff",	--6043
		x"ff",	--6044
		x"ff",	--6045
		x"ff",	--6046
		x"ff",	--6047
		x"ff",	--6048
		x"ff",	--6049
		x"ff",	--6050
		x"ff",	--6051
		x"ff",	--6052
		x"ff",	--6053
		x"ff",	--6054
		x"ff",	--6055
		x"ff",	--6056
		x"ff",	--6057
		x"ff",	--6058
		x"ff",	--6059
		x"ff",	--6060
		x"ff",	--6061
		x"ff",	--6062
		x"ff",	--6063
		x"ff",	--6064
		x"ff",	--6065
		x"ff",	--6066
		x"ff",	--6067
		x"ff",	--6068
		x"ff",	--6069
		x"ff",	--6070
		x"ff",	--6071
		x"ff",	--6072
		x"ff",	--6073
		x"ff",	--6074
		x"ff",	--6075
		x"ff",	--6076
		x"ff",	--6077
		x"ff",	--6078
		x"ff",	--6079
		x"ff",	--6080
		x"ff",	--6081
		x"ff",	--6082
		x"ff",	--6083
		x"ff",	--6084
		x"ff",	--6085
		x"ff",	--6086
		x"ff",	--6087
		x"ff",	--6088
		x"ff",	--6089
		x"ff",	--6090
		x"ff",	--6091
		x"ff",	--6092
		x"ff",	--6093
		x"ff",	--6094
		x"ff",	--6095
		x"ff",	--6096
		x"ff",	--6097
		x"ff",	--6098
		x"ff",	--6099
		x"ff",	--6100
		x"ff",	--6101
		x"ff",	--6102
		x"ff",	--6103
		x"ff",	--6104
		x"ff",	--6105
		x"ff",	--6106
		x"ff",	--6107
		x"ff",	--6108
		x"ff",	--6109
		x"ff",	--6110
		x"ff",	--6111
		x"ff",	--6112
		x"ff",	--6113
		x"ff",	--6114
		x"ff",	--6115
		x"ff",	--6116
		x"ff",	--6117
		x"ff",	--6118
		x"ff",	--6119
		x"ff",	--6120
		x"ff",	--6121
		x"ff",	--6122
		x"ff",	--6123
		x"ff",	--6124
		x"ff",	--6125
		x"ff",	--6126
		x"ff",	--6127
		x"ff",	--6128
		x"ff",	--6129
		x"ff",	--6130
		x"ff",	--6131
		x"ff",	--6132
		x"ff",	--6133
		x"ff",	--6134
		x"ff",	--6135
		x"ff",	--6136
		x"ff",	--6137
		x"ff",	--6138
		x"ff",	--6139
		x"ff",	--6140
		x"ff",	--6141
		x"ff",	--6142
		x"ff",	--6143
		x"ff",	--6144
		x"ff",	--6145
		x"ff",	--6146
		x"ff",	--6147
		x"ff",	--6148
		x"ff",	--6149
		x"ff",	--6150
		x"ff",	--6151
		x"ff",	--6152
		x"ff",	--6153
		x"ff",	--6154
		x"ff",	--6155
		x"ff",	--6156
		x"ff",	--6157
		x"ff",	--6158
		x"ff",	--6159
		x"ff",	--6160
		x"ff",	--6161
		x"ff",	--6162
		x"ff",	--6163
		x"ff",	--6164
		x"ff",	--6165
		x"ff",	--6166
		x"ff",	--6167
		x"ff",	--6168
		x"ff",	--6169
		x"ff",	--6170
		x"ff",	--6171
		x"ff",	--6172
		x"ff",	--6173
		x"ff",	--6174
		x"ff",	--6175
		x"ff",	--6176
		x"ff",	--6177
		x"ff",	--6178
		x"ff",	--6179
		x"ff",	--6180
		x"ff",	--6181
		x"ff",	--6182
		x"ff",	--6183
		x"ff",	--6184
		x"ff",	--6185
		x"ff",	--6186
		x"ff",	--6187
		x"ff",	--6188
		x"ff",	--6189
		x"ff",	--6190
		x"ff",	--6191
		x"ff",	--6192
		x"ff",	--6193
		x"ff",	--6194
		x"ff",	--6195
		x"ff",	--6196
		x"ff",	--6197
		x"ff",	--6198
		x"ff",	--6199
		x"ff",	--6200
		x"ff",	--6201
		x"ff",	--6202
		x"ff",	--6203
		x"ff",	--6204
		x"ff",	--6205
		x"ff",	--6206
		x"ff",	--6207
		x"ff",	--6208
		x"ff",	--6209
		x"ff",	--6210
		x"ff",	--6211
		x"ff",	--6212
		x"ff",	--6213
		x"ff",	--6214
		x"ff",	--6215
		x"ff",	--6216
		x"ff",	--6217
		x"ff",	--6218
		x"ff",	--6219
		x"ff",	--6220
		x"ff",	--6221
		x"ff",	--6222
		x"ff",	--6223
		x"ff",	--6224
		x"ff",	--6225
		x"ff",	--6226
		x"ff",	--6227
		x"ff",	--6228
		x"ff",	--6229
		x"ff",	--6230
		x"ff",	--6231
		x"ff",	--6232
		x"ff",	--6233
		x"ff",	--6234
		x"ff",	--6235
		x"ff",	--6236
		x"ff",	--6237
		x"ff",	--6238
		x"ff",	--6239
		x"ff",	--6240
		x"ff",	--6241
		x"ff",	--6242
		x"ff",	--6243
		x"ff",	--6244
		x"ff",	--6245
		x"ff",	--6246
		x"ff",	--6247
		x"ff",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"ff",	--6252
		x"ff",	--6253
		x"ff",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"3c",	--8176
		x"3c",	--8177
		x"3c",	--8178
		x"3c",	--8179
		x"3c",	--8180
		x"3c",	--8181
		x"3c",	--8182
		x"fe",	--8183
		x"80",	--8184
		x"3c",	--8185
		x"3c",	--8186
		x"3c",	--8187
		x"3c",	--8188
		x"3c",	--8189
		x"3c",	--8190
		x"00");	--8191
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"e9",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"ce",	--44
		x"12",	--45
		x"c8",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"e6",	--50
		x"12",	--51
		x"cd",	--52
		x"53",	--53
		x"40",	--54
		x"e7",	--55
		x"40",	--56
		x"c5",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"c9",	--61
		x"40",	--62
		x"e7",	--63
		x"40",	--64
		x"c6",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"c9",	--69
		x"40",	--70
		x"e7",	--71
		x"40",	--72
		x"c6",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"c9",	--77
		x"40",	--78
		x"e7",	--79
		x"40",	--80
		x"c3",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"c9",	--85
		x"40",	--86
		x"e7",	--87
		x"40",	--88
		x"c4",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"c9",	--93
		x"40",	--94
		x"e7",	--95
		x"40",	--96
		x"c2",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"c9",	--101
		x"40",	--102
		x"e7",	--103
		x"40",	--104
		x"c2",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"c9",	--109
		x"40",	--110
		x"e7",	--111
		x"40",	--112
		x"c2",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"c9",	--117
		x"43",	--118
		x"43",	--119
		x"12",	--120
		x"c8",	--121
		x"43",	--122
		x"40",	--123
		x"4e",	--124
		x"40",	--125
		x"01",	--126
		x"41",	--127
		x"50",	--128
		x"00",	--129
		x"12",	--130
		x"c7",	--131
		x"41",	--132
		x"50",	--133
		x"00",	--134
		x"12",	--135
		x"c8",	--136
		x"43",	--137
		x"40",	--138
		x"4e",	--139
		x"40",	--140
		x"01",	--141
		x"41",	--142
		x"52",	--143
		x"12",	--144
		x"c7",	--145
		x"41",	--146
		x"52",	--147
		x"12",	--148
		x"c8",	--149
		x"41",	--150
		x"52",	--151
		x"41",	--152
		x"50",	--153
		x"00",	--154
		x"12",	--155
		x"c3",	--156
		x"40",	--157
		x"01",	--158
		x"41",	--159
		x"53",	--160
		x"12",	--161
		x"cb",	--162
		x"40",	--163
		x"01",	--164
		x"41",	--165
		x"12",	--166
		x"cb",	--167
		x"41",	--168
		x"41",	--169
		x"53",	--170
		x"12",	--171
		x"c4",	--172
		x"41",	--173
		x"52",	--174
		x"41",	--175
		x"50",	--176
		x"00",	--177
		x"12",	--178
		x"c4",	--179
		x"12",	--180
		x"c9",	--181
		x"40",	--182
		x"00",	--183
		x"40",	--184
		x"c5",	--185
		x"12",	--186
		x"ca",	--187
		x"43",	--188
		x"40",	--189
		x"03",	--190
		x"12",	--191
		x"ca",	--192
		x"43",	--193
		x"43",	--194
		x"43",	--195
		x"41",	--196
		x"50",	--197
		x"00",	--198
		x"12",	--199
		x"c3",	--200
		x"43",	--201
		x"43",	--202
		x"43",	--203
		x"41",	--204
		x"50",	--205
		x"00",	--206
		x"12",	--207
		x"c3",	--208
		x"41",	--209
		x"50",	--210
		x"00",	--211
		x"41",	--212
		x"50",	--213
		x"00",	--214
		x"12",	--215
		x"c2",	--216
		x"40",	--217
		x"ff",	--218
		x"00",	--219
		x"d2",	--220
		x"43",	--221
		x"12",	--222
		x"ce",	--223
		x"93",	--224
		x"27",	--225
		x"12",	--226
		x"ce",	--227
		x"92",	--228
		x"24",	--229
		x"90",	--230
		x"00",	--231
		x"20",	--232
		x"12",	--233
		x"e7",	--234
		x"12",	--235
		x"cd",	--236
		x"53",	--237
		x"40",	--238
		x"00",	--239
		x"51",	--240
		x"5f",	--241
		x"43",	--242
		x"00",	--243
		x"4f",	--244
		x"41",	--245
		x"00",	--246
		x"12",	--247
		x"c9",	--248
		x"43",	--249
		x"3f",	--250
		x"93",	--251
		x"27",	--252
		x"53",	--253
		x"12",	--254
		x"e7",	--255
		x"12",	--256
		x"cd",	--257
		x"53",	--258
		x"3f",	--259
		x"90",	--260
		x"00",	--261
		x"2f",	--262
		x"93",	--263
		x"02",	--264
		x"24",	--265
		x"4f",	--266
		x"11",	--267
		x"12",	--268
		x"12",	--269
		x"e7",	--270
		x"4f",	--271
		x"00",	--272
		x"12",	--273
		x"cd",	--274
		x"52",	--275
		x"41",	--276
		x"00",	--277
		x"40",	--278
		x"00",	--279
		x"51",	--280
		x"5b",	--281
		x"4f",	--282
		x"00",	--283
		x"53",	--284
		x"3f",	--285
		x"40",	--286
		x"e6",	--287
		x"4e",	--288
		x"00",	--289
		x"4d",	--290
		x"00",	--291
		x"4c",	--292
		x"00",	--293
		x"43",	--294
		x"00",	--295
		x"43",	--296
		x"00",	--297
		x"43",	--298
		x"00",	--299
		x"41",	--300
		x"43",	--301
		x"00",	--302
		x"43",	--303
		x"00",	--304
		x"43",	--305
		x"00",	--306
		x"41",	--307
		x"4e",	--308
		x"00",	--309
		x"41",	--310
		x"4e",	--311
		x"00",	--312
		x"41",	--313
		x"4e",	--314
		x"00",	--315
		x"41",	--316
		x"4e",	--317
		x"00",	--318
		x"41",	--319
		x"4f",	--320
		x"00",	--321
		x"8e",	--322
		x"4d",	--323
		x"5f",	--324
		x"00",	--325
		x"4d",	--326
		x"00",	--327
		x"12",	--328
		x"c2",	--329
		x"43",	--330
		x"4e",	--331
		x"01",	--332
		x"4f",	--333
		x"01",	--334
		x"42",	--335
		x"01",	--336
		x"41",	--337
		x"12",	--338
		x"c2",	--339
		x"43",	--340
		x"4d",	--341
		x"01",	--342
		x"4f",	--343
		x"00",	--344
		x"01",	--345
		x"42",	--346
		x"01",	--347
		x"41",	--348
		x"5c",	--349
		x"8f",	--350
		x"00",	--351
		x"12",	--352
		x"c2",	--353
		x"43",	--354
		x"4e",	--355
		x"01",	--356
		x"4f",	--357
		x"00",	--358
		x"01",	--359
		x"42",	--360
		x"01",	--361
		x"41",	--362
		x"5d",	--363
		x"41",	--364
		x"41",	--365
		x"43",	--366
		x"41",	--367
		x"43",	--368
		x"41",	--369
		x"40",	--370
		x"c0",	--371
		x"01",	--372
		x"40",	--373
		x"00",	--374
		x"01",	--375
		x"40",	--376
		x"02",	--377
		x"01",	--378
		x"12",	--379
		x"e6",	--380
		x"12",	--381
		x"cd",	--382
		x"43",	--383
		x"01",	--384
		x"40",	--385
		x"e6",	--386
		x"00",	--387
		x"12",	--388
		x"cd",	--389
		x"53",	--390
		x"43",	--391
		x"41",	--392
		x"12",	--393
		x"c2",	--394
		x"41",	--395
		x"12",	--396
		x"12",	--397
		x"43",	--398
		x"40",	--399
		x"3f",	--400
		x"4a",	--401
		x"4b",	--402
		x"42",	--403
		x"02",	--404
		x"12",	--405
		x"c8",	--406
		x"4a",	--407
		x"4b",	--408
		x"42",	--409
		x"02",	--410
		x"12",	--411
		x"c8",	--412
		x"12",	--413
		x"e6",	--414
		x"12",	--415
		x"cd",	--416
		x"53",	--417
		x"41",	--418
		x"41",	--419
		x"41",	--420
		x"4f",	--421
		x"02",	--422
		x"4e",	--423
		x"02",	--424
		x"41",	--425
		x"12",	--426
		x"12",	--427
		x"83",	--428
		x"4f",	--429
		x"4e",	--430
		x"93",	--431
		x"02",	--432
		x"24",	--433
		x"90",	--434
		x"00",	--435
		x"38",	--436
		x"20",	--437
		x"41",	--438
		x"4b",	--439
		x"00",	--440
		x"12",	--441
		x"c6",	--442
		x"4f",	--443
		x"41",	--444
		x"4b",	--445
		x"00",	--446
		x"12",	--447
		x"c6",	--448
		x"4f",	--449
		x"12",	--450
		x"12",	--451
		x"12",	--452
		x"e6",	--453
		x"12",	--454
		x"cd",	--455
		x"50",	--456
		x"00",	--457
		x"4a",	--458
		x"43",	--459
		x"12",	--460
		x"d6",	--461
		x"43",	--462
		x"40",	--463
		x"42",	--464
		x"12",	--465
		x"d4",	--466
		x"4e",	--467
		x"4f",	--468
		x"43",	--469
		x"40",	--470
		x"3f",	--471
		x"12",	--472
		x"d1",	--473
		x"4e",	--474
		x"4f",	--475
		x"42",	--476
		x"02",	--477
		x"12",	--478
		x"c8",	--479
		x"4b",	--480
		x"43",	--481
		x"12",	--482
		x"d6",	--483
		x"43",	--484
		x"40",	--485
		x"42",	--486
		x"12",	--487
		x"d4",	--488
		x"4e",	--489
		x"4f",	--490
		x"42",	--491
		x"02",	--492
		x"12",	--493
		x"c8",	--494
		x"43",	--495
		x"53",	--496
		x"41",	--497
		x"41",	--498
		x"41",	--499
		x"41",	--500
		x"4b",	--501
		x"00",	--502
		x"12",	--503
		x"c6",	--504
		x"43",	--505
		x"4f",	--506
		x"42",	--507
		x"02",	--508
		x"12",	--509
		x"ca",	--510
		x"3f",	--511
		x"43",	--512
		x"40",	--513
		x"c3",	--514
		x"12",	--515
		x"ca",	--516
		x"4f",	--517
		x"02",	--518
		x"3f",	--519
		x"12",	--520
		x"e6",	--521
		x"12",	--522
		x"cd",	--523
		x"40",	--524
		x"e6",	--525
		x"00",	--526
		x"12",	--527
		x"cd",	--528
		x"4b",	--529
		x"00",	--530
		x"12",	--531
		x"e6",	--532
		x"12",	--533
		x"cd",	--534
		x"52",	--535
		x"43",	--536
		x"3f",	--537
		x"12",	--538
		x"12",	--539
		x"42",	--540
		x"02",	--541
		x"12",	--542
		x"cb",	--543
		x"4e",	--544
		x"4f",	--545
		x"42",	--546
		x"02",	--547
		x"12",	--548
		x"cb",	--549
		x"12",	--550
		x"12",	--551
		x"e3",	--552
		x"e3",	--553
		x"53",	--554
		x"63",	--555
		x"12",	--556
		x"12",	--557
		x"12",	--558
		x"e6",	--559
		x"12",	--560
		x"02",	--561
		x"12",	--562
		x"db",	--563
		x"50",	--564
		x"00",	--565
		x"12",	--566
		x"02",	--567
		x"12",	--568
		x"e6",	--569
		x"12",	--570
		x"cd",	--571
		x"52",	--572
		x"41",	--573
		x"41",	--574
		x"41",	--575
		x"4f",	--576
		x"02",	--577
		x"4e",	--578
		x"02",	--579
		x"41",	--580
		x"4f",	--581
		x"02",	--582
		x"4e",	--583
		x"02",	--584
		x"41",	--585
		x"12",	--586
		x"12",	--587
		x"12",	--588
		x"12",	--589
		x"83",	--590
		x"4f",	--591
		x"4e",	--592
		x"43",	--593
		x"00",	--594
		x"93",	--595
		x"24",	--596
		x"93",	--597
		x"02",	--598
		x"24",	--599
		x"43",	--600
		x"02",	--601
		x"41",	--602
		x"4b",	--603
		x"00",	--604
		x"12",	--605
		x"c6",	--606
		x"4f",	--607
		x"90",	--608
		x"00",	--609
		x"34",	--610
		x"43",	--611
		x"49",	--612
		x"48",	--613
		x"42",	--614
		x"02",	--615
		x"12",	--616
		x"ca",	--617
		x"43",	--618
		x"53",	--619
		x"41",	--620
		x"41",	--621
		x"41",	--622
		x"41",	--623
		x"41",	--624
		x"93",	--625
		x"02",	--626
		x"24",	--627
		x"43",	--628
		x"02",	--629
		x"42",	--630
		x"02",	--631
		x"12",	--632
		x"ca",	--633
		x"43",	--634
		x"53",	--635
		x"41",	--636
		x"41",	--637
		x"41",	--638
		x"41",	--639
		x"41",	--640
		x"41",	--641
		x"4b",	--642
		x"00",	--643
		x"12",	--644
		x"c6",	--645
		x"4f",	--646
		x"90",	--647
		x"00",	--648
		x"3b",	--649
		x"41",	--650
		x"4b",	--651
		x"00",	--652
		x"12",	--653
		x"c6",	--654
		x"4f",	--655
		x"41",	--656
		x"4b",	--657
		x"00",	--658
		x"12",	--659
		x"c6",	--660
		x"4f",	--661
		x"12",	--662
		x"12",	--663
		x"12",	--664
		x"e6",	--665
		x"12",	--666
		x"cd",	--667
		x"50",	--668
		x"00",	--669
		x"4a",	--670
		x"43",	--671
		x"12",	--672
		x"d6",	--673
		x"43",	--674
		x"40",	--675
		x"42",	--676
		x"12",	--677
		x"d4",	--678
		x"4e",	--679
		x"4f",	--680
		x"42",	--681
		x"02",	--682
		x"12",	--683
		x"c8",	--684
		x"4b",	--685
		x"43",	--686
		x"12",	--687
		x"d6",	--688
		x"43",	--689
		x"40",	--690
		x"42",	--691
		x"12",	--692
		x"d4",	--693
		x"4e",	--694
		x"4f",	--695
		x"42",	--696
		x"02",	--697
		x"12",	--698
		x"c8",	--699
		x"3f",	--700
		x"43",	--701
		x"12",	--702
		x"c4",	--703
		x"43",	--704
		x"53",	--705
		x"41",	--706
		x"41",	--707
		x"41",	--708
		x"41",	--709
		x"41",	--710
		x"43",	--711
		x"40",	--712
		x"c4",	--713
		x"12",	--714
		x"ca",	--715
		x"4f",	--716
		x"02",	--717
		x"3f",	--718
		x"42",	--719
		x"00",	--720
		x"4e",	--721
		x"be",	--722
		x"20",	--723
		x"df",	--724
		x"00",	--725
		x"41",	--726
		x"cf",	--727
		x"00",	--728
		x"41",	--729
		x"43",	--730
		x"93",	--731
		x"02",	--732
		x"24",	--733
		x"43",	--734
		x"4f",	--735
		x"02",	--736
		x"43",	--737
		x"41",	--738
		x"42",	--739
		x"02",	--740
		x"92",	--741
		x"2c",	--742
		x"4e",	--743
		x"5f",	--744
		x"4f",	--745
		x"e6",	--746
		x"43",	--747
		x"00",	--748
		x"90",	--749
		x"00",	--750
		x"38",	--751
		x"43",	--752
		x"02",	--753
		x"41",	--754
		x"53",	--755
		x"4e",	--756
		x"02",	--757
		x"41",	--758
		x"40",	--759
		x"00",	--760
		x"00",	--761
		x"3f",	--762
		x"40",	--763
		x"00",	--764
		x"00",	--765
		x"3f",	--766
		x"42",	--767
		x"00",	--768
		x"3f",	--769
		x"40",	--770
		x"00",	--771
		x"00",	--772
		x"3f",	--773
		x"40",	--774
		x"00",	--775
		x"00",	--776
		x"3f",	--777
		x"40",	--778
		x"00",	--779
		x"00",	--780
		x"3f",	--781
		x"40",	--782
		x"00",	--783
		x"00",	--784
		x"3f",	--785
		x"12",	--786
		x"12",	--787
		x"83",	--788
		x"4f",	--789
		x"4e",	--790
		x"12",	--791
		x"e7",	--792
		x"12",	--793
		x"cd",	--794
		x"53",	--795
		x"90",	--796
		x"00",	--797
		x"38",	--798
		x"41",	--799
		x"4b",	--800
		x"00",	--801
		x"12",	--802
		x"c6",	--803
		x"4f",	--804
		x"41",	--805
		x"4b",	--806
		x"00",	--807
		x"12",	--808
		x"c6",	--809
		x"4f",	--810
		x"12",	--811
		x"12",	--812
		x"12",	--813
		x"e7",	--814
		x"12",	--815
		x"cd",	--816
		x"50",	--817
		x"00",	--818
		x"4b",	--819
		x"00",	--820
		x"43",	--821
		x"53",	--822
		x"41",	--823
		x"41",	--824
		x"41",	--825
		x"12",	--826
		x"e7",	--827
		x"12",	--828
		x"cd",	--829
		x"40",	--830
		x"e7",	--831
		x"00",	--832
		x"12",	--833
		x"cd",	--834
		x"4b",	--835
		x"00",	--836
		x"12",	--837
		x"e7",	--838
		x"12",	--839
		x"cd",	--840
		x"52",	--841
		x"43",	--842
		x"3f",	--843
		x"12",	--844
		x"83",	--845
		x"4e",	--846
		x"93",	--847
		x"24",	--848
		x"38",	--849
		x"12",	--850
		x"e7",	--851
		x"12",	--852
		x"cd",	--853
		x"53",	--854
		x"41",	--855
		x"4b",	--856
		x"00",	--857
		x"12",	--858
		x"c6",	--859
		x"12",	--860
		x"12",	--861
		x"12",	--862
		x"e7",	--863
		x"12",	--864
		x"cd",	--865
		x"50",	--866
		x"00",	--867
		x"43",	--868
		x"53",	--869
		x"41",	--870
		x"41",	--871
		x"12",	--872
		x"e7",	--873
		x"12",	--874
		x"cd",	--875
		x"40",	--876
		x"e7",	--877
		x"00",	--878
		x"12",	--879
		x"cd",	--880
		x"4b",	--881
		x"00",	--882
		x"12",	--883
		x"e7",	--884
		x"12",	--885
		x"cd",	--886
		x"52",	--887
		x"43",	--888
		x"3f",	--889
		x"12",	--890
		x"12",	--891
		x"43",	--892
		x"00",	--893
		x"4f",	--894
		x"93",	--895
		x"24",	--896
		x"53",	--897
		x"43",	--898
		x"43",	--899
		x"3c",	--900
		x"90",	--901
		x"00",	--902
		x"2c",	--903
		x"5c",	--904
		x"5c",	--905
		x"5c",	--906
		x"5c",	--907
		x"11",	--908
		x"5d",	--909
		x"50",	--910
		x"ff",	--911
		x"43",	--912
		x"4f",	--913
		x"93",	--914
		x"24",	--915
		x"90",	--916
		x"00",	--917
		x"24",	--918
		x"4d",	--919
		x"50",	--920
		x"ff",	--921
		x"93",	--922
		x"23",	--923
		x"90",	--924
		x"00",	--925
		x"2c",	--926
		x"5c",	--927
		x"4c",	--928
		x"5b",	--929
		x"5b",	--930
		x"5b",	--931
		x"11",	--932
		x"5d",	--933
		x"50",	--934
		x"ff",	--935
		x"4f",	--936
		x"93",	--937
		x"23",	--938
		x"43",	--939
		x"00",	--940
		x"4c",	--941
		x"41",	--942
		x"41",	--943
		x"41",	--944
		x"43",	--945
		x"3f",	--946
		x"4d",	--947
		x"50",	--948
		x"ff",	--949
		x"90",	--950
		x"00",	--951
		x"2c",	--952
		x"5c",	--953
		x"5c",	--954
		x"5c",	--955
		x"5c",	--956
		x"11",	--957
		x"5d",	--958
		x"50",	--959
		x"ff",	--960
		x"43",	--961
		x"3f",	--962
		x"4d",	--963
		x"50",	--964
		x"ff",	--965
		x"90",	--966
		x"00",	--967
		x"2c",	--968
		x"5c",	--969
		x"5c",	--970
		x"5c",	--971
		x"5c",	--972
		x"11",	--973
		x"5d",	--974
		x"50",	--975
		x"ff",	--976
		x"43",	--977
		x"3f",	--978
		x"11",	--979
		x"12",	--980
		x"12",	--981
		x"e7",	--982
		x"12",	--983
		x"cd",	--984
		x"52",	--985
		x"43",	--986
		x"4c",	--987
		x"41",	--988
		x"41",	--989
		x"41",	--990
		x"43",	--991
		x"3f",	--992
		x"12",	--993
		x"12",	--994
		x"4e",	--995
		x"4c",	--996
		x"4e",	--997
		x"00",	--998
		x"4d",	--999
		x"00",	--1000
		x"4c",	--1001
		x"00",	--1002
		x"4d",	--1003
		x"43",	--1004
		x"40",	--1005
		x"36",	--1006
		x"40",	--1007
		x"01",	--1008
		x"12",	--1009
		x"e4",	--1010
		x"4e",	--1011
		x"00",	--1012
		x"12",	--1013
		x"c2",	--1014
		x"43",	--1015
		x"4a",	--1016
		x"01",	--1017
		x"40",	--1018
		x"00",	--1019
		x"01",	--1020
		x"42",	--1021
		x"01",	--1022
		x"00",	--1023
		x"41",	--1024
		x"43",	--1025
		x"41",	--1026
		x"41",	--1027
		x"41",	--1028
		x"12",	--1029
		x"12",	--1030
		x"12",	--1031
		x"43",	--1032
		x"00",	--1033
		x"40",	--1034
		x"3f",	--1035
		x"00",	--1036
		x"4f",	--1037
		x"4b",	--1038
		x"00",	--1039
		x"43",	--1040
		x"12",	--1041
		x"d6",	--1042
		x"43",	--1043
		x"40",	--1044
		x"3f",	--1045
		x"12",	--1046
		x"d2",	--1047
		x"4e",	--1048
		x"4f",	--1049
		x"4b",	--1050
		x"00",	--1051
		x"43",	--1052
		x"12",	--1053
		x"d6",	--1054
		x"4e",	--1055
		x"4f",	--1056
		x"48",	--1057
		x"49",	--1058
		x"12",	--1059
		x"d1",	--1060
		x"12",	--1061
		x"ce",	--1062
		x"4e",	--1063
		x"00",	--1064
		x"43",	--1065
		x"00",	--1066
		x"41",	--1067
		x"41",	--1068
		x"41",	--1069
		x"41",	--1070
		x"12",	--1071
		x"12",	--1072
		x"12",	--1073
		x"4d",	--1074
		x"4e",	--1075
		x"4d",	--1076
		x"00",	--1077
		x"4e",	--1078
		x"00",	--1079
		x"4f",	--1080
		x"49",	--1081
		x"00",	--1082
		x"43",	--1083
		x"12",	--1084
		x"d6",	--1085
		x"4e",	--1086
		x"4f",	--1087
		x"4a",	--1088
		x"4b",	--1089
		x"12",	--1090
		x"d2",	--1091
		x"4e",	--1092
		x"4f",	--1093
		x"49",	--1094
		x"00",	--1095
		x"43",	--1096
		x"12",	--1097
		x"d6",	--1098
		x"4e",	--1099
		x"4f",	--1100
		x"4a",	--1101
		x"4b",	--1102
		x"12",	--1103
		x"d1",	--1104
		x"12",	--1105
		x"ce",	--1106
		x"4e",	--1107
		x"00",	--1108
		x"41",	--1109
		x"41",	--1110
		x"41",	--1111
		x"41",	--1112
		x"4f",	--1113
		x"4e",	--1114
		x"00",	--1115
		x"41",	--1116
		x"12",	--1117
		x"12",	--1118
		x"93",	--1119
		x"02",	--1120
		x"38",	--1121
		x"40",	--1122
		x"02",	--1123
		x"43",	--1124
		x"12",	--1125
		x"4b",	--1126
		x"ff",	--1127
		x"11",	--1128
		x"12",	--1129
		x"12",	--1130
		x"e7",	--1131
		x"12",	--1132
		x"cd",	--1133
		x"50",	--1134
		x"00",	--1135
		x"53",	--1136
		x"50",	--1137
		x"00",	--1138
		x"92",	--1139
		x"02",	--1140
		x"3b",	--1141
		x"43",	--1142
		x"41",	--1143
		x"41",	--1144
		x"41",	--1145
		x"42",	--1146
		x"02",	--1147
		x"90",	--1148
		x"00",	--1149
		x"34",	--1150
		x"4e",	--1151
		x"5f",	--1152
		x"5e",	--1153
		x"5f",	--1154
		x"50",	--1155
		x"02",	--1156
		x"40",	--1157
		x"00",	--1158
		x"00",	--1159
		x"40",	--1160
		x"c8",	--1161
		x"00",	--1162
		x"40",	--1163
		x"02",	--1164
		x"00",	--1165
		x"53",	--1166
		x"4e",	--1167
		x"02",	--1168
		x"41",	--1169
		x"12",	--1170
		x"42",	--1171
		x"02",	--1172
		x"90",	--1173
		x"00",	--1174
		x"34",	--1175
		x"4b",	--1176
		x"5c",	--1177
		x"5b",	--1178
		x"5c",	--1179
		x"50",	--1180
		x"02",	--1181
		x"4f",	--1182
		x"00",	--1183
		x"4e",	--1184
		x"00",	--1185
		x"4d",	--1186
		x"00",	--1187
		x"53",	--1188
		x"4b",	--1189
		x"02",	--1190
		x"43",	--1191
		x"41",	--1192
		x"41",	--1193
		x"43",	--1194
		x"3f",	--1195
		x"12",	--1196
		x"50",	--1197
		x"ff",	--1198
		x"42",	--1199
		x"02",	--1200
		x"93",	--1201
		x"38",	--1202
		x"92",	--1203
		x"02",	--1204
		x"24",	--1205
		x"40",	--1206
		x"02",	--1207
		x"43",	--1208
		x"3c",	--1209
		x"50",	--1210
		x"00",	--1211
		x"9f",	--1212
		x"ff",	--1213
		x"24",	--1214
		x"53",	--1215
		x"9b",	--1216
		x"23",	--1217
		x"12",	--1218
		x"e7",	--1219
		x"12",	--1220
		x"cd",	--1221
		x"53",	--1222
		x"43",	--1223
		x"50",	--1224
		x"00",	--1225
		x"41",	--1226
		x"41",	--1227
		x"43",	--1228
		x"4e",	--1229
		x"00",	--1230
		x"4e",	--1231
		x"93",	--1232
		x"24",	--1233
		x"53",	--1234
		x"43",	--1235
		x"3c",	--1236
		x"4e",	--1237
		x"93",	--1238
		x"24",	--1239
		x"53",	--1240
		x"92",	--1241
		x"34",	--1242
		x"90",	--1243
		x"00",	--1244
		x"23",	--1245
		x"43",	--1246
		x"ff",	--1247
		x"4f",	--1248
		x"5d",	--1249
		x"51",	--1250
		x"4e",	--1251
		x"00",	--1252
		x"53",	--1253
		x"4e",	--1254
		x"93",	--1255
		x"23",	--1256
		x"4c",	--1257
		x"5e",	--1258
		x"5e",	--1259
		x"5c",	--1260
		x"50",	--1261
		x"02",	--1262
		x"41",	--1263
		x"12",	--1264
		x"00",	--1265
		x"50",	--1266
		x"00",	--1267
		x"41",	--1268
		x"41",	--1269
		x"43",	--1270
		x"3f",	--1271
		x"d0",	--1272
		x"02",	--1273
		x"01",	--1274
		x"40",	--1275
		x"0b",	--1276
		x"01",	--1277
		x"43",	--1278
		x"41",	--1279
		x"12",	--1280
		x"4f",	--1281
		x"42",	--1282
		x"02",	--1283
		x"90",	--1284
		x"00",	--1285
		x"34",	--1286
		x"4f",	--1287
		x"5c",	--1288
		x"4c",	--1289
		x"5d",	--1290
		x"5d",	--1291
		x"5d",	--1292
		x"8c",	--1293
		x"50",	--1294
		x"03",	--1295
		x"43",	--1296
		x"00",	--1297
		x"43",	--1298
		x"00",	--1299
		x"43",	--1300
		x"00",	--1301
		x"4b",	--1302
		x"00",	--1303
		x"4e",	--1304
		x"00",	--1305
		x"4f",	--1306
		x"53",	--1307
		x"4e",	--1308
		x"02",	--1309
		x"41",	--1310
		x"41",	--1311
		x"43",	--1312
		x"3f",	--1313
		x"5f",	--1314
		x"4f",	--1315
		x"5c",	--1316
		x"5c",	--1317
		x"5c",	--1318
		x"8f",	--1319
		x"50",	--1320
		x"03",	--1321
		x"43",	--1322
		x"00",	--1323
		x"4e",	--1324
		x"00",	--1325
		x"43",	--1326
		x"00",	--1327
		x"4d",	--1328
		x"00",	--1329
		x"43",	--1330
		x"00",	--1331
		x"43",	--1332
		x"41",	--1333
		x"5f",	--1334
		x"4f",	--1335
		x"5e",	--1336
		x"5e",	--1337
		x"5e",	--1338
		x"8f",	--1339
		x"43",	--1340
		x"03",	--1341
		x"43",	--1342
		x"41",	--1343
		x"12",	--1344
		x"12",	--1345
		x"12",	--1346
		x"12",	--1347
		x"12",	--1348
		x"12",	--1349
		x"12",	--1350
		x"12",	--1351
		x"12",	--1352
		x"93",	--1353
		x"02",	--1354
		x"38",	--1355
		x"40",	--1356
		x"03",	--1357
		x"4a",	--1358
		x"53",	--1359
		x"4a",	--1360
		x"52",	--1361
		x"4a",	--1362
		x"50",	--1363
		x"00",	--1364
		x"43",	--1365
		x"3c",	--1366
		x"53",	--1367
		x"4f",	--1368
		x"00",	--1369
		x"53",	--1370
		x"50",	--1371
		x"00",	--1372
		x"50",	--1373
		x"00",	--1374
		x"50",	--1375
		x"00",	--1376
		x"50",	--1377
		x"00",	--1378
		x"92",	--1379
		x"02",	--1380
		x"34",	--1381
		x"93",	--1382
		x"00",	--1383
		x"27",	--1384
		x"4b",	--1385
		x"9b",	--1386
		x"00",	--1387
		x"2b",	--1388
		x"43",	--1389
		x"00",	--1390
		x"4b",	--1391
		x"00",	--1392
		x"12",	--1393
		x"00",	--1394
		x"93",	--1395
		x"00",	--1396
		x"27",	--1397
		x"47",	--1398
		x"53",	--1399
		x"4f",	--1400
		x"00",	--1401
		x"98",	--1402
		x"2b",	--1403
		x"43",	--1404
		x"00",	--1405
		x"3f",	--1406
		x"f0",	--1407
		x"ff",	--1408
		x"01",	--1409
		x"41",	--1410
		x"41",	--1411
		x"41",	--1412
		x"41",	--1413
		x"41",	--1414
		x"41",	--1415
		x"41",	--1416
		x"41",	--1417
		x"41",	--1418
		x"13",	--1419
		x"4e",	--1420
		x"00",	--1421
		x"43",	--1422
		x"41",	--1423
		x"4f",	--1424
		x"4f",	--1425
		x"4f",	--1426
		x"00",	--1427
		x"41",	--1428
		x"42",	--1429
		x"00",	--1430
		x"f2",	--1431
		x"23",	--1432
		x"4f",	--1433
		x"00",	--1434
		x"43",	--1435
		x"41",	--1436
		x"f0",	--1437
		x"00",	--1438
		x"4f",	--1439
		x"e8",	--1440
		x"11",	--1441
		x"12",	--1442
		x"cb",	--1443
		x"41",	--1444
		x"12",	--1445
		x"4f",	--1446
		x"4f",	--1447
		x"11",	--1448
		x"11",	--1449
		x"11",	--1450
		x"11",	--1451
		x"4e",	--1452
		x"12",	--1453
		x"cb",	--1454
		x"4b",	--1455
		x"12",	--1456
		x"cb",	--1457
		x"41",	--1458
		x"41",	--1459
		x"12",	--1460
		x"12",	--1461
		x"4f",	--1462
		x"40",	--1463
		x"00",	--1464
		x"4a",	--1465
		x"4b",	--1466
		x"f0",	--1467
		x"00",	--1468
		x"24",	--1469
		x"11",	--1470
		x"53",	--1471
		x"23",	--1472
		x"f3",	--1473
		x"24",	--1474
		x"40",	--1475
		x"00",	--1476
		x"12",	--1477
		x"cb",	--1478
		x"53",	--1479
		x"93",	--1480
		x"23",	--1481
		x"41",	--1482
		x"41",	--1483
		x"41",	--1484
		x"40",	--1485
		x"00",	--1486
		x"3f",	--1487
		x"12",	--1488
		x"4f",	--1489
		x"4f",	--1490
		x"10",	--1491
		x"11",	--1492
		x"4e",	--1493
		x"12",	--1494
		x"cb",	--1495
		x"4b",	--1496
		x"12",	--1497
		x"cb",	--1498
		x"41",	--1499
		x"41",	--1500
		x"12",	--1501
		x"12",	--1502
		x"4e",	--1503
		x"4f",	--1504
		x"4f",	--1505
		x"10",	--1506
		x"11",	--1507
		x"4d",	--1508
		x"12",	--1509
		x"cb",	--1510
		x"4b",	--1511
		x"12",	--1512
		x"cb",	--1513
		x"4b",	--1514
		x"4a",	--1515
		x"10",	--1516
		x"10",	--1517
		x"ec",	--1518
		x"ec",	--1519
		x"4d",	--1520
		x"12",	--1521
		x"cb",	--1522
		x"4a",	--1523
		x"12",	--1524
		x"cb",	--1525
		x"41",	--1526
		x"41",	--1527
		x"41",	--1528
		x"12",	--1529
		x"12",	--1530
		x"12",	--1531
		x"4f",	--1532
		x"93",	--1533
		x"24",	--1534
		x"4e",	--1535
		x"53",	--1536
		x"43",	--1537
		x"4a",	--1538
		x"5b",	--1539
		x"4d",	--1540
		x"11",	--1541
		x"12",	--1542
		x"cb",	--1543
		x"99",	--1544
		x"24",	--1545
		x"53",	--1546
		x"b0",	--1547
		x"00",	--1548
		x"20",	--1549
		x"40",	--1550
		x"00",	--1551
		x"12",	--1552
		x"cb",	--1553
		x"3f",	--1554
		x"40",	--1555
		x"00",	--1556
		x"12",	--1557
		x"cb",	--1558
		x"3f",	--1559
		x"41",	--1560
		x"41",	--1561
		x"41",	--1562
		x"41",	--1563
		x"12",	--1564
		x"12",	--1565
		x"12",	--1566
		x"4f",	--1567
		x"93",	--1568
		x"24",	--1569
		x"4e",	--1570
		x"53",	--1571
		x"43",	--1572
		x"4a",	--1573
		x"11",	--1574
		x"12",	--1575
		x"cb",	--1576
		x"99",	--1577
		x"24",	--1578
		x"53",	--1579
		x"b0",	--1580
		x"00",	--1581
		x"23",	--1582
		x"40",	--1583
		x"00",	--1584
		x"12",	--1585
		x"cb",	--1586
		x"4a",	--1587
		x"11",	--1588
		x"12",	--1589
		x"cb",	--1590
		x"99",	--1591
		x"23",	--1592
		x"41",	--1593
		x"41",	--1594
		x"41",	--1595
		x"41",	--1596
		x"12",	--1597
		x"12",	--1598
		x"12",	--1599
		x"50",	--1600
		x"ff",	--1601
		x"4f",	--1602
		x"93",	--1603
		x"38",	--1604
		x"90",	--1605
		x"00",	--1606
		x"38",	--1607
		x"43",	--1608
		x"41",	--1609
		x"59",	--1610
		x"40",	--1611
		x"00",	--1612
		x"4b",	--1613
		x"12",	--1614
		x"e4",	--1615
		x"50",	--1616
		x"00",	--1617
		x"4f",	--1618
		x"00",	--1619
		x"53",	--1620
		x"40",	--1621
		x"00",	--1622
		x"4b",	--1623
		x"12",	--1624
		x"e4",	--1625
		x"4f",	--1626
		x"90",	--1627
		x"00",	--1628
		x"37",	--1629
		x"49",	--1630
		x"53",	--1631
		x"51",	--1632
		x"40",	--1633
		x"00",	--1634
		x"4b",	--1635
		x"12",	--1636
		x"e4",	--1637
		x"50",	--1638
		x"00",	--1639
		x"4f",	--1640
		x"00",	--1641
		x"53",	--1642
		x"41",	--1643
		x"5a",	--1644
		x"4f",	--1645
		x"11",	--1646
		x"12",	--1647
		x"cb",	--1648
		x"93",	--1649
		x"23",	--1650
		x"50",	--1651
		x"00",	--1652
		x"41",	--1653
		x"41",	--1654
		x"41",	--1655
		x"41",	--1656
		x"40",	--1657
		x"00",	--1658
		x"12",	--1659
		x"cb",	--1660
		x"e3",	--1661
		x"53",	--1662
		x"3f",	--1663
		x"43",	--1664
		x"43",	--1665
		x"3f",	--1666
		x"12",	--1667
		x"12",	--1668
		x"12",	--1669
		x"41",	--1670
		x"52",	--1671
		x"4b",	--1672
		x"49",	--1673
		x"93",	--1674
		x"20",	--1675
		x"3c",	--1676
		x"11",	--1677
		x"12",	--1678
		x"cb",	--1679
		x"49",	--1680
		x"4a",	--1681
		x"53",	--1682
		x"4a",	--1683
		x"00",	--1684
		x"93",	--1685
		x"24",	--1686
		x"90",	--1687
		x"00",	--1688
		x"23",	--1689
		x"49",	--1690
		x"53",	--1691
		x"49",	--1692
		x"00",	--1693
		x"50",	--1694
		x"ff",	--1695
		x"90",	--1696
		x"00",	--1697
		x"2f",	--1698
		x"4f",	--1699
		x"5f",	--1700
		x"4f",	--1701
		x"e8",	--1702
		x"41",	--1703
		x"41",	--1704
		x"41",	--1705
		x"41",	--1706
		x"4b",	--1707
		x"52",	--1708
		x"4b",	--1709
		x"00",	--1710
		x"4b",	--1711
		x"12",	--1712
		x"cb",	--1713
		x"49",	--1714
		x"3f",	--1715
		x"4b",	--1716
		x"53",	--1717
		x"4b",	--1718
		x"12",	--1719
		x"cb",	--1720
		x"49",	--1721
		x"3f",	--1722
		x"4b",	--1723
		x"53",	--1724
		x"4f",	--1725
		x"49",	--1726
		x"93",	--1727
		x"27",	--1728
		x"53",	--1729
		x"11",	--1730
		x"12",	--1731
		x"cb",	--1732
		x"49",	--1733
		x"93",	--1734
		x"23",	--1735
		x"3f",	--1736
		x"4b",	--1737
		x"52",	--1738
		x"4b",	--1739
		x"00",	--1740
		x"4b",	--1741
		x"12",	--1742
		x"cc",	--1743
		x"49",	--1744
		x"3f",	--1745
		x"4b",	--1746
		x"53",	--1747
		x"4b",	--1748
		x"4e",	--1749
		x"10",	--1750
		x"11",	--1751
		x"10",	--1752
		x"11",	--1753
		x"12",	--1754
		x"cb",	--1755
		x"49",	--1756
		x"3f",	--1757
		x"4b",	--1758
		x"53",	--1759
		x"4b",	--1760
		x"12",	--1761
		x"cc",	--1762
		x"49",	--1763
		x"3f",	--1764
		x"4b",	--1765
		x"53",	--1766
		x"4b",	--1767
		x"12",	--1768
		x"cb",	--1769
		x"49",	--1770
		x"3f",	--1771
		x"4b",	--1772
		x"53",	--1773
		x"4b",	--1774
		x"12",	--1775
		x"cb",	--1776
		x"49",	--1777
		x"3f",	--1778
		x"4b",	--1779
		x"53",	--1780
		x"4b",	--1781
		x"12",	--1782
		x"cb",	--1783
		x"49",	--1784
		x"3f",	--1785
		x"40",	--1786
		x"00",	--1787
		x"12",	--1788
		x"cb",	--1789
		x"3f",	--1790
		x"12",	--1791
		x"12",	--1792
		x"42",	--1793
		x"02",	--1794
		x"42",	--1795
		x"00",	--1796
		x"04",	--1797
		x"42",	--1798
		x"02",	--1799
		x"90",	--1800
		x"00",	--1801
		x"34",	--1802
		x"53",	--1803
		x"02",	--1804
		x"42",	--1805
		x"02",	--1806
		x"42",	--1807
		x"02",	--1808
		x"9f",	--1809
		x"20",	--1810
		x"53",	--1811
		x"02",	--1812
		x"40",	--1813
		x"00",	--1814
		x"00",	--1815
		x"41",	--1816
		x"41",	--1817
		x"c0",	--1818
		x"00",	--1819
		x"00",	--1820
		x"13",	--1821
		x"43",	--1822
		x"02",	--1823
		x"3f",	--1824
		x"4e",	--1825
		x"4f",	--1826
		x"40",	--1827
		x"36",	--1828
		x"40",	--1829
		x"01",	--1830
		x"12",	--1831
		x"e4",	--1832
		x"53",	--1833
		x"4e",	--1834
		x"00",	--1835
		x"40",	--1836
		x"00",	--1837
		x"00",	--1838
		x"41",	--1839
		x"42",	--1840
		x"02",	--1841
		x"42",	--1842
		x"02",	--1843
		x"9f",	--1844
		x"38",	--1845
		x"42",	--1846
		x"02",	--1847
		x"82",	--1848
		x"02",	--1849
		x"41",	--1850
		x"42",	--1851
		x"02",	--1852
		x"42",	--1853
		x"02",	--1854
		x"40",	--1855
		x"00",	--1856
		x"8d",	--1857
		x"8e",	--1858
		x"41",	--1859
		x"42",	--1860
		x"02",	--1861
		x"4f",	--1862
		x"04",	--1863
		x"42",	--1864
		x"02",	--1865
		x"42",	--1866
		x"02",	--1867
		x"9e",	--1868
		x"24",	--1869
		x"42",	--1870
		x"02",	--1871
		x"90",	--1872
		x"00",	--1873
		x"38",	--1874
		x"43",	--1875
		x"02",	--1876
		x"41",	--1877
		x"53",	--1878
		x"02",	--1879
		x"41",	--1880
		x"43",	--1881
		x"41",	--1882
		x"12",	--1883
		x"12",	--1884
		x"4e",	--1885
		x"4f",	--1886
		x"43",	--1887
		x"40",	--1888
		x"4f",	--1889
		x"12",	--1890
		x"d5",	--1891
		x"93",	--1892
		x"34",	--1893
		x"4a",	--1894
		x"4b",	--1895
		x"12",	--1896
		x"d5",	--1897
		x"41",	--1898
		x"41",	--1899
		x"41",	--1900
		x"43",	--1901
		x"40",	--1902
		x"4f",	--1903
		x"4a",	--1904
		x"4b",	--1905
		x"12",	--1906
		x"d1",	--1907
		x"12",	--1908
		x"d5",	--1909
		x"53",	--1910
		x"60",	--1911
		x"80",	--1912
		x"41",	--1913
		x"41",	--1914
		x"41",	--1915
		x"12",	--1916
		x"12",	--1917
		x"12",	--1918
		x"12",	--1919
		x"12",	--1920
		x"12",	--1921
		x"12",	--1922
		x"12",	--1923
		x"50",	--1924
		x"ff",	--1925
		x"4d",	--1926
		x"4f",	--1927
		x"93",	--1928
		x"28",	--1929
		x"4e",	--1930
		x"93",	--1931
		x"28",	--1932
		x"92",	--1933
		x"20",	--1934
		x"40",	--1935
		x"d1",	--1936
		x"92",	--1937
		x"24",	--1938
		x"93",	--1939
		x"24",	--1940
		x"93",	--1941
		x"24",	--1942
		x"4f",	--1943
		x"00",	--1944
		x"00",	--1945
		x"4e",	--1946
		x"00",	--1947
		x"4f",	--1948
		x"00",	--1949
		x"4f",	--1950
		x"00",	--1951
		x"4e",	--1952
		x"00",	--1953
		x"4e",	--1954
		x"00",	--1955
		x"41",	--1956
		x"8b",	--1957
		x"4c",	--1958
		x"93",	--1959
		x"38",	--1960
		x"90",	--1961
		x"00",	--1962
		x"34",	--1963
		x"93",	--1964
		x"38",	--1965
		x"46",	--1966
		x"00",	--1967
		x"47",	--1968
		x"00",	--1969
		x"49",	--1970
		x"f0",	--1971
		x"00",	--1972
		x"24",	--1973
		x"46",	--1974
		x"47",	--1975
		x"c3",	--1976
		x"10",	--1977
		x"10",	--1978
		x"53",	--1979
		x"23",	--1980
		x"4a",	--1981
		x"00",	--1982
		x"4b",	--1983
		x"00",	--1984
		x"43",	--1985
		x"43",	--1986
		x"f0",	--1987
		x"00",	--1988
		x"24",	--1989
		x"5c",	--1990
		x"6d",	--1991
		x"53",	--1992
		x"23",	--1993
		x"53",	--1994
		x"63",	--1995
		x"f6",	--1996
		x"f7",	--1997
		x"43",	--1998
		x"43",	--1999
		x"93",	--2000
		x"20",	--2001
		x"93",	--2002
		x"24",	--2003
		x"41",	--2004
		x"00",	--2005
		x"41",	--2006
		x"00",	--2007
		x"da",	--2008
		x"db",	--2009
		x"4f",	--2010
		x"00",	--2011
		x"9e",	--2012
		x"00",	--2013
		x"20",	--2014
		x"4f",	--2015
		x"00",	--2016
		x"41",	--2017
		x"00",	--2018
		x"46",	--2019
		x"47",	--2020
		x"54",	--2021
		x"65",	--2022
		x"4e",	--2023
		x"00",	--2024
		x"4f",	--2025
		x"00",	--2026
		x"40",	--2027
		x"00",	--2028
		x"00",	--2029
		x"93",	--2030
		x"38",	--2031
		x"48",	--2032
		x"50",	--2033
		x"00",	--2034
		x"41",	--2035
		x"41",	--2036
		x"41",	--2037
		x"41",	--2038
		x"41",	--2039
		x"41",	--2040
		x"41",	--2041
		x"41",	--2042
		x"41",	--2043
		x"91",	--2044
		x"38",	--2045
		x"4b",	--2046
		x"00",	--2047
		x"43",	--2048
		x"43",	--2049
		x"4f",	--2050
		x"00",	--2051
		x"9e",	--2052
		x"00",	--2053
		x"27",	--2054
		x"93",	--2055
		x"24",	--2056
		x"46",	--2057
		x"47",	--2058
		x"84",	--2059
		x"75",	--2060
		x"93",	--2061
		x"38",	--2062
		x"43",	--2063
		x"00",	--2064
		x"41",	--2065
		x"00",	--2066
		x"4e",	--2067
		x"00",	--2068
		x"4f",	--2069
		x"00",	--2070
		x"4e",	--2071
		x"4f",	--2072
		x"53",	--2073
		x"63",	--2074
		x"90",	--2075
		x"3f",	--2076
		x"28",	--2077
		x"90",	--2078
		x"40",	--2079
		x"2c",	--2080
		x"93",	--2081
		x"2c",	--2082
		x"48",	--2083
		x"00",	--2084
		x"53",	--2085
		x"5e",	--2086
		x"6f",	--2087
		x"4b",	--2088
		x"53",	--2089
		x"4e",	--2090
		x"4f",	--2091
		x"53",	--2092
		x"63",	--2093
		x"90",	--2094
		x"3f",	--2095
		x"2b",	--2096
		x"24",	--2097
		x"4e",	--2098
		x"00",	--2099
		x"4f",	--2100
		x"00",	--2101
		x"4a",	--2102
		x"00",	--2103
		x"40",	--2104
		x"00",	--2105
		x"00",	--2106
		x"93",	--2107
		x"37",	--2108
		x"4e",	--2109
		x"4f",	--2110
		x"f3",	--2111
		x"f3",	--2112
		x"c3",	--2113
		x"10",	--2114
		x"10",	--2115
		x"4c",	--2116
		x"4d",	--2117
		x"de",	--2118
		x"df",	--2119
		x"4a",	--2120
		x"00",	--2121
		x"4b",	--2122
		x"00",	--2123
		x"53",	--2124
		x"00",	--2125
		x"48",	--2126
		x"3f",	--2127
		x"93",	--2128
		x"23",	--2129
		x"4f",	--2130
		x"00",	--2131
		x"4f",	--2132
		x"00",	--2133
		x"00",	--2134
		x"4f",	--2135
		x"00",	--2136
		x"00",	--2137
		x"4f",	--2138
		x"00",	--2139
		x"00",	--2140
		x"4e",	--2141
		x"00",	--2142
		x"ff",	--2143
		x"00",	--2144
		x"4e",	--2145
		x"00",	--2146
		x"4d",	--2147
		x"3f",	--2148
		x"43",	--2149
		x"43",	--2150
		x"3f",	--2151
		x"e3",	--2152
		x"53",	--2153
		x"90",	--2154
		x"00",	--2155
		x"37",	--2156
		x"3f",	--2157
		x"93",	--2158
		x"2b",	--2159
		x"3f",	--2160
		x"44",	--2161
		x"45",	--2162
		x"86",	--2163
		x"77",	--2164
		x"3f",	--2165
		x"4e",	--2166
		x"3f",	--2167
		x"43",	--2168
		x"00",	--2169
		x"41",	--2170
		x"00",	--2171
		x"e3",	--2172
		x"e3",	--2173
		x"53",	--2174
		x"63",	--2175
		x"4e",	--2176
		x"00",	--2177
		x"4f",	--2178
		x"00",	--2179
		x"3f",	--2180
		x"93",	--2181
		x"27",	--2182
		x"59",	--2183
		x"00",	--2184
		x"44",	--2185
		x"00",	--2186
		x"45",	--2187
		x"00",	--2188
		x"49",	--2189
		x"f0",	--2190
		x"00",	--2191
		x"24",	--2192
		x"4d",	--2193
		x"44",	--2194
		x"45",	--2195
		x"c3",	--2196
		x"10",	--2197
		x"10",	--2198
		x"53",	--2199
		x"23",	--2200
		x"4c",	--2201
		x"00",	--2202
		x"4d",	--2203
		x"00",	--2204
		x"43",	--2205
		x"43",	--2206
		x"f0",	--2207
		x"00",	--2208
		x"24",	--2209
		x"5c",	--2210
		x"6d",	--2211
		x"53",	--2212
		x"23",	--2213
		x"53",	--2214
		x"63",	--2215
		x"f4",	--2216
		x"f5",	--2217
		x"43",	--2218
		x"43",	--2219
		x"93",	--2220
		x"20",	--2221
		x"93",	--2222
		x"20",	--2223
		x"43",	--2224
		x"43",	--2225
		x"41",	--2226
		x"00",	--2227
		x"41",	--2228
		x"00",	--2229
		x"da",	--2230
		x"db",	--2231
		x"3f",	--2232
		x"43",	--2233
		x"43",	--2234
		x"3f",	--2235
		x"92",	--2236
		x"23",	--2237
		x"9e",	--2238
		x"00",	--2239
		x"00",	--2240
		x"27",	--2241
		x"40",	--2242
		x"e8",	--2243
		x"3f",	--2244
		x"50",	--2245
		x"ff",	--2246
		x"4e",	--2247
		x"00",	--2248
		x"4f",	--2249
		x"00",	--2250
		x"4c",	--2251
		x"00",	--2252
		x"4d",	--2253
		x"00",	--2254
		x"41",	--2255
		x"50",	--2256
		x"00",	--2257
		x"41",	--2258
		x"52",	--2259
		x"12",	--2260
		x"d9",	--2261
		x"41",	--2262
		x"50",	--2263
		x"00",	--2264
		x"41",	--2265
		x"12",	--2266
		x"d9",	--2267
		x"41",	--2268
		x"52",	--2269
		x"41",	--2270
		x"50",	--2271
		x"00",	--2272
		x"41",	--2273
		x"50",	--2274
		x"00",	--2275
		x"12",	--2276
		x"ce",	--2277
		x"12",	--2278
		x"d7",	--2279
		x"50",	--2280
		x"00",	--2281
		x"41",	--2282
		x"50",	--2283
		x"ff",	--2284
		x"4e",	--2285
		x"00",	--2286
		x"4f",	--2287
		x"00",	--2288
		x"4c",	--2289
		x"00",	--2290
		x"4d",	--2291
		x"00",	--2292
		x"41",	--2293
		x"50",	--2294
		x"00",	--2295
		x"41",	--2296
		x"52",	--2297
		x"12",	--2298
		x"d9",	--2299
		x"41",	--2300
		x"50",	--2301
		x"00",	--2302
		x"41",	--2303
		x"12",	--2304
		x"d9",	--2305
		x"e3",	--2306
		x"00",	--2307
		x"41",	--2308
		x"52",	--2309
		x"41",	--2310
		x"50",	--2311
		x"00",	--2312
		x"41",	--2313
		x"50",	--2314
		x"00",	--2315
		x"12",	--2316
		x"ce",	--2317
		x"12",	--2318
		x"d7",	--2319
		x"50",	--2320
		x"00",	--2321
		x"41",	--2322
		x"12",	--2323
		x"12",	--2324
		x"12",	--2325
		x"12",	--2326
		x"12",	--2327
		x"12",	--2328
		x"12",	--2329
		x"12",	--2330
		x"50",	--2331
		x"ff",	--2332
		x"4e",	--2333
		x"00",	--2334
		x"4f",	--2335
		x"00",	--2336
		x"4c",	--2337
		x"00",	--2338
		x"4d",	--2339
		x"00",	--2340
		x"41",	--2341
		x"50",	--2342
		x"00",	--2343
		x"41",	--2344
		x"52",	--2345
		x"12",	--2346
		x"d9",	--2347
		x"41",	--2348
		x"50",	--2349
		x"00",	--2350
		x"41",	--2351
		x"12",	--2352
		x"d9",	--2353
		x"41",	--2354
		x"00",	--2355
		x"93",	--2356
		x"28",	--2357
		x"41",	--2358
		x"00",	--2359
		x"93",	--2360
		x"28",	--2361
		x"92",	--2362
		x"24",	--2363
		x"92",	--2364
		x"24",	--2365
		x"93",	--2366
		x"24",	--2367
		x"93",	--2368
		x"24",	--2369
		x"41",	--2370
		x"00",	--2371
		x"41",	--2372
		x"00",	--2373
		x"41",	--2374
		x"00",	--2375
		x"41",	--2376
		x"00",	--2377
		x"40",	--2378
		x"00",	--2379
		x"43",	--2380
		x"43",	--2381
		x"43",	--2382
		x"43",	--2383
		x"43",	--2384
		x"00",	--2385
		x"43",	--2386
		x"00",	--2387
		x"43",	--2388
		x"43",	--2389
		x"4c",	--2390
		x"00",	--2391
		x"3c",	--2392
		x"58",	--2393
		x"69",	--2394
		x"c3",	--2395
		x"10",	--2396
		x"10",	--2397
		x"53",	--2398
		x"00",	--2399
		x"24",	--2400
		x"b3",	--2401
		x"24",	--2402
		x"58",	--2403
		x"69",	--2404
		x"56",	--2405
		x"67",	--2406
		x"43",	--2407
		x"43",	--2408
		x"99",	--2409
		x"28",	--2410
		x"24",	--2411
		x"43",	--2412
		x"43",	--2413
		x"5c",	--2414
		x"6d",	--2415
		x"56",	--2416
		x"67",	--2417
		x"93",	--2418
		x"37",	--2419
		x"d3",	--2420
		x"d3",	--2421
		x"3f",	--2422
		x"98",	--2423
		x"2b",	--2424
		x"3f",	--2425
		x"4a",	--2426
		x"00",	--2427
		x"4b",	--2428
		x"00",	--2429
		x"4f",	--2430
		x"41",	--2431
		x"00",	--2432
		x"51",	--2433
		x"00",	--2434
		x"4a",	--2435
		x"53",	--2436
		x"46",	--2437
		x"00",	--2438
		x"43",	--2439
		x"91",	--2440
		x"00",	--2441
		x"00",	--2442
		x"24",	--2443
		x"4d",	--2444
		x"00",	--2445
		x"93",	--2446
		x"38",	--2447
		x"90",	--2448
		x"40",	--2449
		x"2c",	--2450
		x"41",	--2451
		x"00",	--2452
		x"53",	--2453
		x"41",	--2454
		x"00",	--2455
		x"41",	--2456
		x"00",	--2457
		x"4d",	--2458
		x"5e",	--2459
		x"6f",	--2460
		x"93",	--2461
		x"38",	--2462
		x"5a",	--2463
		x"6b",	--2464
		x"53",	--2465
		x"90",	--2466
		x"40",	--2467
		x"2b",	--2468
		x"4a",	--2469
		x"00",	--2470
		x"4b",	--2471
		x"00",	--2472
		x"4c",	--2473
		x"00",	--2474
		x"4e",	--2475
		x"4f",	--2476
		x"f0",	--2477
		x"00",	--2478
		x"f3",	--2479
		x"90",	--2480
		x"00",	--2481
		x"24",	--2482
		x"4e",	--2483
		x"00",	--2484
		x"4f",	--2485
		x"00",	--2486
		x"40",	--2487
		x"00",	--2488
		x"00",	--2489
		x"41",	--2490
		x"52",	--2491
		x"12",	--2492
		x"d7",	--2493
		x"50",	--2494
		x"00",	--2495
		x"41",	--2496
		x"41",	--2497
		x"41",	--2498
		x"41",	--2499
		x"41",	--2500
		x"41",	--2501
		x"41",	--2502
		x"41",	--2503
		x"41",	--2504
		x"d3",	--2505
		x"d3",	--2506
		x"3f",	--2507
		x"50",	--2508
		x"00",	--2509
		x"4a",	--2510
		x"b3",	--2511
		x"24",	--2512
		x"41",	--2513
		x"00",	--2514
		x"41",	--2515
		x"00",	--2516
		x"c3",	--2517
		x"10",	--2518
		x"10",	--2519
		x"4c",	--2520
		x"4d",	--2521
		x"d3",	--2522
		x"d0",	--2523
		x"80",	--2524
		x"46",	--2525
		x"00",	--2526
		x"47",	--2527
		x"00",	--2528
		x"c3",	--2529
		x"10",	--2530
		x"10",	--2531
		x"53",	--2532
		x"93",	--2533
		x"3b",	--2534
		x"48",	--2535
		x"00",	--2536
		x"3f",	--2537
		x"93",	--2538
		x"24",	--2539
		x"43",	--2540
		x"91",	--2541
		x"00",	--2542
		x"00",	--2543
		x"24",	--2544
		x"4f",	--2545
		x"00",	--2546
		x"41",	--2547
		x"50",	--2548
		x"00",	--2549
		x"3f",	--2550
		x"93",	--2551
		x"23",	--2552
		x"4e",	--2553
		x"4f",	--2554
		x"f0",	--2555
		x"00",	--2556
		x"f3",	--2557
		x"93",	--2558
		x"23",	--2559
		x"93",	--2560
		x"23",	--2561
		x"93",	--2562
		x"00",	--2563
		x"20",	--2564
		x"93",	--2565
		x"00",	--2566
		x"27",	--2567
		x"50",	--2568
		x"00",	--2569
		x"63",	--2570
		x"f0",	--2571
		x"ff",	--2572
		x"f3",	--2573
		x"3f",	--2574
		x"43",	--2575
		x"3f",	--2576
		x"43",	--2577
		x"3f",	--2578
		x"43",	--2579
		x"91",	--2580
		x"00",	--2581
		x"00",	--2582
		x"24",	--2583
		x"4f",	--2584
		x"00",	--2585
		x"41",	--2586
		x"50",	--2587
		x"00",	--2588
		x"3f",	--2589
		x"43",	--2590
		x"3f",	--2591
		x"93",	--2592
		x"23",	--2593
		x"40",	--2594
		x"e8",	--2595
		x"3f",	--2596
		x"12",	--2597
		x"12",	--2598
		x"12",	--2599
		x"12",	--2600
		x"12",	--2601
		x"50",	--2602
		x"ff",	--2603
		x"4e",	--2604
		x"00",	--2605
		x"4f",	--2606
		x"00",	--2607
		x"4c",	--2608
		x"00",	--2609
		x"4d",	--2610
		x"00",	--2611
		x"41",	--2612
		x"50",	--2613
		x"00",	--2614
		x"41",	--2615
		x"52",	--2616
		x"12",	--2617
		x"d9",	--2618
		x"41",	--2619
		x"52",	--2620
		x"41",	--2621
		x"12",	--2622
		x"d9",	--2623
		x"41",	--2624
		x"00",	--2625
		x"93",	--2626
		x"28",	--2627
		x"41",	--2628
		x"00",	--2629
		x"93",	--2630
		x"28",	--2631
		x"e1",	--2632
		x"00",	--2633
		x"00",	--2634
		x"92",	--2635
		x"24",	--2636
		x"93",	--2637
		x"24",	--2638
		x"92",	--2639
		x"24",	--2640
		x"93",	--2641
		x"24",	--2642
		x"41",	--2643
		x"00",	--2644
		x"81",	--2645
		x"00",	--2646
		x"4d",	--2647
		x"00",	--2648
		x"41",	--2649
		x"00",	--2650
		x"41",	--2651
		x"00",	--2652
		x"41",	--2653
		x"00",	--2654
		x"41",	--2655
		x"00",	--2656
		x"99",	--2657
		x"2c",	--2658
		x"5e",	--2659
		x"6f",	--2660
		x"53",	--2661
		x"4d",	--2662
		x"00",	--2663
		x"40",	--2664
		x"00",	--2665
		x"43",	--2666
		x"40",	--2667
		x"40",	--2668
		x"43",	--2669
		x"43",	--2670
		x"3c",	--2671
		x"dc",	--2672
		x"dd",	--2673
		x"88",	--2674
		x"79",	--2675
		x"c3",	--2676
		x"10",	--2677
		x"10",	--2678
		x"5e",	--2679
		x"6f",	--2680
		x"53",	--2681
		x"24",	--2682
		x"99",	--2683
		x"2b",	--2684
		x"23",	--2685
		x"98",	--2686
		x"2b",	--2687
		x"3f",	--2688
		x"9f",	--2689
		x"2b",	--2690
		x"98",	--2691
		x"2f",	--2692
		x"3f",	--2693
		x"4a",	--2694
		x"4b",	--2695
		x"f0",	--2696
		x"00",	--2697
		x"f3",	--2698
		x"90",	--2699
		x"00",	--2700
		x"24",	--2701
		x"4a",	--2702
		x"00",	--2703
		x"4b",	--2704
		x"00",	--2705
		x"41",	--2706
		x"50",	--2707
		x"00",	--2708
		x"12",	--2709
		x"d7",	--2710
		x"50",	--2711
		x"00",	--2712
		x"41",	--2713
		x"41",	--2714
		x"41",	--2715
		x"41",	--2716
		x"41",	--2717
		x"41",	--2718
		x"42",	--2719
		x"00",	--2720
		x"41",	--2721
		x"50",	--2722
		x"00",	--2723
		x"3f",	--2724
		x"9e",	--2725
		x"23",	--2726
		x"40",	--2727
		x"e8",	--2728
		x"3f",	--2729
		x"93",	--2730
		x"23",	--2731
		x"4a",	--2732
		x"4b",	--2733
		x"f0",	--2734
		x"00",	--2735
		x"f3",	--2736
		x"93",	--2737
		x"23",	--2738
		x"93",	--2739
		x"23",	--2740
		x"93",	--2741
		x"20",	--2742
		x"93",	--2743
		x"27",	--2744
		x"50",	--2745
		x"00",	--2746
		x"63",	--2747
		x"f0",	--2748
		x"ff",	--2749
		x"f3",	--2750
		x"3f",	--2751
		x"43",	--2752
		x"00",	--2753
		x"43",	--2754
		x"00",	--2755
		x"43",	--2756
		x"00",	--2757
		x"41",	--2758
		x"50",	--2759
		x"00",	--2760
		x"3f",	--2761
		x"41",	--2762
		x"52",	--2763
		x"3f",	--2764
		x"50",	--2765
		x"ff",	--2766
		x"4e",	--2767
		x"00",	--2768
		x"4f",	--2769
		x"00",	--2770
		x"4c",	--2771
		x"00",	--2772
		x"4d",	--2773
		x"00",	--2774
		x"41",	--2775
		x"50",	--2776
		x"00",	--2777
		x"41",	--2778
		x"52",	--2779
		x"12",	--2780
		x"d9",	--2781
		x"41",	--2782
		x"52",	--2783
		x"41",	--2784
		x"12",	--2785
		x"d9",	--2786
		x"93",	--2787
		x"00",	--2788
		x"28",	--2789
		x"93",	--2790
		x"00",	--2791
		x"28",	--2792
		x"41",	--2793
		x"52",	--2794
		x"41",	--2795
		x"50",	--2796
		x"00",	--2797
		x"12",	--2798
		x"da",	--2799
		x"50",	--2800
		x"00",	--2801
		x"41",	--2802
		x"43",	--2803
		x"3f",	--2804
		x"50",	--2805
		x"ff",	--2806
		x"4e",	--2807
		x"00",	--2808
		x"4f",	--2809
		x"00",	--2810
		x"41",	--2811
		x"52",	--2812
		x"41",	--2813
		x"12",	--2814
		x"d9",	--2815
		x"41",	--2816
		x"00",	--2817
		x"93",	--2818
		x"24",	--2819
		x"28",	--2820
		x"92",	--2821
		x"24",	--2822
		x"41",	--2823
		x"00",	--2824
		x"93",	--2825
		x"38",	--2826
		x"90",	--2827
		x"00",	--2828
		x"38",	--2829
		x"93",	--2830
		x"00",	--2831
		x"20",	--2832
		x"43",	--2833
		x"40",	--2834
		x"7f",	--2835
		x"50",	--2836
		x"00",	--2837
		x"41",	--2838
		x"41",	--2839
		x"00",	--2840
		x"41",	--2841
		x"00",	--2842
		x"40",	--2843
		x"00",	--2844
		x"8d",	--2845
		x"4c",	--2846
		x"f0",	--2847
		x"00",	--2848
		x"20",	--2849
		x"93",	--2850
		x"00",	--2851
		x"27",	--2852
		x"e3",	--2853
		x"e3",	--2854
		x"53",	--2855
		x"63",	--2856
		x"50",	--2857
		x"00",	--2858
		x"41",	--2859
		x"43",	--2860
		x"43",	--2861
		x"50",	--2862
		x"00",	--2863
		x"41",	--2864
		x"c3",	--2865
		x"10",	--2866
		x"10",	--2867
		x"53",	--2868
		x"23",	--2869
		x"3f",	--2870
		x"43",	--2871
		x"40",	--2872
		x"80",	--2873
		x"50",	--2874
		x"00",	--2875
		x"41",	--2876
		x"12",	--2877
		x"12",	--2878
		x"12",	--2879
		x"12",	--2880
		x"82",	--2881
		x"4e",	--2882
		x"4f",	--2883
		x"43",	--2884
		x"00",	--2885
		x"93",	--2886
		x"20",	--2887
		x"93",	--2888
		x"20",	--2889
		x"43",	--2890
		x"00",	--2891
		x"41",	--2892
		x"12",	--2893
		x"d7",	--2894
		x"52",	--2895
		x"41",	--2896
		x"41",	--2897
		x"41",	--2898
		x"41",	--2899
		x"41",	--2900
		x"40",	--2901
		x"00",	--2902
		x"00",	--2903
		x"40",	--2904
		x"00",	--2905
		x"00",	--2906
		x"4a",	--2907
		x"00",	--2908
		x"4b",	--2909
		x"00",	--2910
		x"4a",	--2911
		x"4b",	--2912
		x"12",	--2913
		x"d7",	--2914
		x"53",	--2915
		x"93",	--2916
		x"38",	--2917
		x"27",	--2918
		x"4a",	--2919
		x"00",	--2920
		x"4b",	--2921
		x"00",	--2922
		x"4f",	--2923
		x"f0",	--2924
		x"00",	--2925
		x"20",	--2926
		x"40",	--2927
		x"00",	--2928
		x"8f",	--2929
		x"4e",	--2930
		x"00",	--2931
		x"3f",	--2932
		x"51",	--2933
		x"00",	--2934
		x"00",	--2935
		x"61",	--2936
		x"00",	--2937
		x"00",	--2938
		x"53",	--2939
		x"23",	--2940
		x"3f",	--2941
		x"4f",	--2942
		x"e3",	--2943
		x"53",	--2944
		x"43",	--2945
		x"43",	--2946
		x"4e",	--2947
		x"f0",	--2948
		x"00",	--2949
		x"24",	--2950
		x"5c",	--2951
		x"6d",	--2952
		x"53",	--2953
		x"23",	--2954
		x"53",	--2955
		x"63",	--2956
		x"fa",	--2957
		x"fb",	--2958
		x"43",	--2959
		x"43",	--2960
		x"93",	--2961
		x"20",	--2962
		x"93",	--2963
		x"20",	--2964
		x"43",	--2965
		x"43",	--2966
		x"f0",	--2967
		x"00",	--2968
		x"20",	--2969
		x"48",	--2970
		x"49",	--2971
		x"da",	--2972
		x"db",	--2973
		x"4d",	--2974
		x"00",	--2975
		x"4e",	--2976
		x"00",	--2977
		x"40",	--2978
		x"00",	--2979
		x"8f",	--2980
		x"4e",	--2981
		x"00",	--2982
		x"3f",	--2983
		x"c3",	--2984
		x"10",	--2985
		x"10",	--2986
		x"53",	--2987
		x"23",	--2988
		x"3f",	--2989
		x"12",	--2990
		x"12",	--2991
		x"12",	--2992
		x"93",	--2993
		x"2c",	--2994
		x"90",	--2995
		x"01",	--2996
		x"28",	--2997
		x"40",	--2998
		x"00",	--2999
		x"43",	--3000
		x"42",	--3001
		x"4e",	--3002
		x"4f",	--3003
		x"49",	--3004
		x"93",	--3005
		x"20",	--3006
		x"50",	--3007
		x"e8",	--3008
		x"4c",	--3009
		x"43",	--3010
		x"8e",	--3011
		x"7f",	--3012
		x"4a",	--3013
		x"41",	--3014
		x"41",	--3015
		x"41",	--3016
		x"41",	--3017
		x"90",	--3018
		x"01",	--3019
		x"28",	--3020
		x"42",	--3021
		x"43",	--3022
		x"40",	--3023
		x"00",	--3024
		x"4e",	--3025
		x"4f",	--3026
		x"49",	--3027
		x"93",	--3028
		x"27",	--3029
		x"c3",	--3030
		x"10",	--3031
		x"10",	--3032
		x"53",	--3033
		x"23",	--3034
		x"3f",	--3035
		x"40",	--3036
		x"00",	--3037
		x"43",	--3038
		x"40",	--3039
		x"00",	--3040
		x"3f",	--3041
		x"40",	--3042
		x"00",	--3043
		x"43",	--3044
		x"43",	--3045
		x"3f",	--3046
		x"12",	--3047
		x"12",	--3048
		x"12",	--3049
		x"12",	--3050
		x"12",	--3051
		x"4f",	--3052
		x"4f",	--3053
		x"00",	--3054
		x"4f",	--3055
		x"00",	--3056
		x"4d",	--3057
		x"00",	--3058
		x"4d",	--3059
		x"93",	--3060
		x"28",	--3061
		x"92",	--3062
		x"24",	--3063
		x"93",	--3064
		x"24",	--3065
		x"93",	--3066
		x"24",	--3067
		x"4d",	--3068
		x"00",	--3069
		x"90",	--3070
		x"ff",	--3071
		x"38",	--3072
		x"90",	--3073
		x"00",	--3074
		x"34",	--3075
		x"4e",	--3076
		x"4f",	--3077
		x"f0",	--3078
		x"00",	--3079
		x"f3",	--3080
		x"90",	--3081
		x"00",	--3082
		x"24",	--3083
		x"50",	--3084
		x"00",	--3085
		x"63",	--3086
		x"93",	--3087
		x"38",	--3088
		x"4b",	--3089
		x"50",	--3090
		x"00",	--3091
		x"c3",	--3092
		x"10",	--3093
		x"10",	--3094
		x"c3",	--3095
		x"10",	--3096
		x"10",	--3097
		x"c3",	--3098
		x"10",	--3099
		x"10",	--3100
		x"c3",	--3101
		x"10",	--3102
		x"10",	--3103
		x"c3",	--3104
		x"10",	--3105
		x"10",	--3106
		x"c3",	--3107
		x"10",	--3108
		x"10",	--3109
		x"c3",	--3110
		x"10",	--3111
		x"10",	--3112
		x"f3",	--3113
		x"f0",	--3114
		x"00",	--3115
		x"4d",	--3116
		x"3c",	--3117
		x"93",	--3118
		x"23",	--3119
		x"43",	--3120
		x"43",	--3121
		x"43",	--3122
		x"4d",	--3123
		x"5d",	--3124
		x"5d",	--3125
		x"5d",	--3126
		x"5d",	--3127
		x"5d",	--3128
		x"5d",	--3129
		x"5d",	--3130
		x"4f",	--3131
		x"f0",	--3132
		x"00",	--3133
		x"dd",	--3134
		x"4a",	--3135
		x"11",	--3136
		x"43",	--3137
		x"10",	--3138
		x"4c",	--3139
		x"df",	--3140
		x"4d",	--3141
		x"41",	--3142
		x"41",	--3143
		x"41",	--3144
		x"41",	--3145
		x"41",	--3146
		x"41",	--3147
		x"93",	--3148
		x"23",	--3149
		x"4e",	--3150
		x"4f",	--3151
		x"f0",	--3152
		x"00",	--3153
		x"f3",	--3154
		x"93",	--3155
		x"20",	--3156
		x"93",	--3157
		x"27",	--3158
		x"50",	--3159
		x"00",	--3160
		x"63",	--3161
		x"3f",	--3162
		x"c3",	--3163
		x"10",	--3164
		x"10",	--3165
		x"4b",	--3166
		x"50",	--3167
		x"00",	--3168
		x"3f",	--3169
		x"43",	--3170
		x"43",	--3171
		x"43",	--3172
		x"3f",	--3173
		x"d3",	--3174
		x"d0",	--3175
		x"00",	--3176
		x"f3",	--3177
		x"f0",	--3178
		x"00",	--3179
		x"43",	--3180
		x"3f",	--3181
		x"40",	--3182
		x"ff",	--3183
		x"8b",	--3184
		x"90",	--3185
		x"00",	--3186
		x"34",	--3187
		x"4e",	--3188
		x"4f",	--3189
		x"47",	--3190
		x"f0",	--3191
		x"00",	--3192
		x"24",	--3193
		x"c3",	--3194
		x"10",	--3195
		x"10",	--3196
		x"53",	--3197
		x"23",	--3198
		x"43",	--3199
		x"43",	--3200
		x"f0",	--3201
		x"00",	--3202
		x"24",	--3203
		x"58",	--3204
		x"69",	--3205
		x"53",	--3206
		x"23",	--3207
		x"53",	--3208
		x"63",	--3209
		x"fe",	--3210
		x"ff",	--3211
		x"43",	--3212
		x"43",	--3213
		x"93",	--3214
		x"20",	--3215
		x"93",	--3216
		x"20",	--3217
		x"43",	--3218
		x"43",	--3219
		x"4e",	--3220
		x"4f",	--3221
		x"dc",	--3222
		x"dd",	--3223
		x"48",	--3224
		x"49",	--3225
		x"f0",	--3226
		x"00",	--3227
		x"f3",	--3228
		x"90",	--3229
		x"00",	--3230
		x"24",	--3231
		x"50",	--3232
		x"00",	--3233
		x"63",	--3234
		x"48",	--3235
		x"49",	--3236
		x"c3",	--3237
		x"10",	--3238
		x"10",	--3239
		x"c3",	--3240
		x"10",	--3241
		x"10",	--3242
		x"c3",	--3243
		x"10",	--3244
		x"10",	--3245
		x"c3",	--3246
		x"10",	--3247
		x"10",	--3248
		x"c3",	--3249
		x"10",	--3250
		x"10",	--3251
		x"c3",	--3252
		x"10",	--3253
		x"10",	--3254
		x"c3",	--3255
		x"10",	--3256
		x"10",	--3257
		x"f3",	--3258
		x"f0",	--3259
		x"00",	--3260
		x"43",	--3261
		x"90",	--3262
		x"40",	--3263
		x"2f",	--3264
		x"43",	--3265
		x"3f",	--3266
		x"43",	--3267
		x"43",	--3268
		x"3f",	--3269
		x"93",	--3270
		x"23",	--3271
		x"48",	--3272
		x"49",	--3273
		x"f0",	--3274
		x"00",	--3275
		x"f3",	--3276
		x"93",	--3277
		x"24",	--3278
		x"50",	--3279
		x"00",	--3280
		x"63",	--3281
		x"3f",	--3282
		x"93",	--3283
		x"27",	--3284
		x"3f",	--3285
		x"12",	--3286
		x"12",	--3287
		x"4f",	--3288
		x"4f",	--3289
		x"00",	--3290
		x"f0",	--3291
		x"00",	--3292
		x"4f",	--3293
		x"00",	--3294
		x"c3",	--3295
		x"10",	--3296
		x"c3",	--3297
		x"10",	--3298
		x"c3",	--3299
		x"10",	--3300
		x"c3",	--3301
		x"10",	--3302
		x"c3",	--3303
		x"10",	--3304
		x"c3",	--3305
		x"10",	--3306
		x"c3",	--3307
		x"10",	--3308
		x"4d",	--3309
		x"4f",	--3310
		x"00",	--3311
		x"b0",	--3312
		x"00",	--3313
		x"43",	--3314
		x"6f",	--3315
		x"4f",	--3316
		x"00",	--3317
		x"93",	--3318
		x"20",	--3319
		x"93",	--3320
		x"24",	--3321
		x"40",	--3322
		x"ff",	--3323
		x"00",	--3324
		x"4a",	--3325
		x"4b",	--3326
		x"5c",	--3327
		x"6d",	--3328
		x"5c",	--3329
		x"6d",	--3330
		x"5c",	--3331
		x"6d",	--3332
		x"5c",	--3333
		x"6d",	--3334
		x"5c",	--3335
		x"6d",	--3336
		x"5c",	--3337
		x"6d",	--3338
		x"5c",	--3339
		x"6d",	--3340
		x"40",	--3341
		x"00",	--3342
		x"00",	--3343
		x"90",	--3344
		x"40",	--3345
		x"2c",	--3346
		x"40",	--3347
		x"ff",	--3348
		x"5c",	--3349
		x"6d",	--3350
		x"4f",	--3351
		x"53",	--3352
		x"90",	--3353
		x"40",	--3354
		x"2b",	--3355
		x"4a",	--3356
		x"00",	--3357
		x"4c",	--3358
		x"00",	--3359
		x"4d",	--3360
		x"00",	--3361
		x"41",	--3362
		x"41",	--3363
		x"41",	--3364
		x"90",	--3365
		x"00",	--3366
		x"24",	--3367
		x"50",	--3368
		x"ff",	--3369
		x"4d",	--3370
		x"00",	--3371
		x"40",	--3372
		x"00",	--3373
		x"00",	--3374
		x"4a",	--3375
		x"4b",	--3376
		x"5c",	--3377
		x"6d",	--3378
		x"5c",	--3379
		x"6d",	--3380
		x"5c",	--3381
		x"6d",	--3382
		x"5c",	--3383
		x"6d",	--3384
		x"5c",	--3385
		x"6d",	--3386
		x"5c",	--3387
		x"6d",	--3388
		x"5c",	--3389
		x"6d",	--3390
		x"4c",	--3391
		x"4d",	--3392
		x"d3",	--3393
		x"d0",	--3394
		x"40",	--3395
		x"4a",	--3396
		x"00",	--3397
		x"4b",	--3398
		x"00",	--3399
		x"41",	--3400
		x"41",	--3401
		x"41",	--3402
		x"93",	--3403
		x"23",	--3404
		x"43",	--3405
		x"00",	--3406
		x"41",	--3407
		x"41",	--3408
		x"41",	--3409
		x"93",	--3410
		x"24",	--3411
		x"4a",	--3412
		x"4b",	--3413
		x"f3",	--3414
		x"f0",	--3415
		x"00",	--3416
		x"93",	--3417
		x"20",	--3418
		x"93",	--3419
		x"24",	--3420
		x"43",	--3421
		x"00",	--3422
		x"3f",	--3423
		x"93",	--3424
		x"23",	--3425
		x"42",	--3426
		x"00",	--3427
		x"3f",	--3428
		x"43",	--3429
		x"00",	--3430
		x"3f",	--3431
		x"12",	--3432
		x"4f",	--3433
		x"93",	--3434
		x"28",	--3435
		x"4e",	--3436
		x"93",	--3437
		x"28",	--3438
		x"92",	--3439
		x"24",	--3440
		x"92",	--3441
		x"24",	--3442
		x"93",	--3443
		x"24",	--3444
		x"93",	--3445
		x"24",	--3446
		x"4f",	--3447
		x"00",	--3448
		x"9e",	--3449
		x"00",	--3450
		x"24",	--3451
		x"93",	--3452
		x"20",	--3453
		x"43",	--3454
		x"4e",	--3455
		x"41",	--3456
		x"41",	--3457
		x"93",	--3458
		x"24",	--3459
		x"93",	--3460
		x"00",	--3461
		x"23",	--3462
		x"43",	--3463
		x"4e",	--3464
		x"41",	--3465
		x"41",	--3466
		x"93",	--3467
		x"00",	--3468
		x"27",	--3469
		x"43",	--3470
		x"3f",	--3471
		x"4f",	--3472
		x"00",	--3473
		x"4e",	--3474
		x"00",	--3475
		x"9b",	--3476
		x"3b",	--3477
		x"9c",	--3478
		x"38",	--3479
		x"4f",	--3480
		x"00",	--3481
		x"4f",	--3482
		x"00",	--3483
		x"4e",	--3484
		x"00",	--3485
		x"4e",	--3486
		x"00",	--3487
		x"9f",	--3488
		x"2b",	--3489
		x"9e",	--3490
		x"28",	--3491
		x"9b",	--3492
		x"2b",	--3493
		x"9e",	--3494
		x"28",	--3495
		x"9f",	--3496
		x"28",	--3497
		x"9c",	--3498
		x"28",	--3499
		x"43",	--3500
		x"3f",	--3501
		x"93",	--3502
		x"23",	--3503
		x"43",	--3504
		x"3f",	--3505
		x"92",	--3506
		x"23",	--3507
		x"4e",	--3508
		x"00",	--3509
		x"4f",	--3510
		x"00",	--3511
		x"8f",	--3512
		x"3f",	--3513
		x"42",	--3514
		x"02",	--3515
		x"93",	--3516
		x"38",	--3517
		x"42",	--3518
		x"02",	--3519
		x"4f",	--3520
		x"00",	--3521
		x"53",	--3522
		x"4d",	--3523
		x"02",	--3524
		x"53",	--3525
		x"4e",	--3526
		x"02",	--3527
		x"41",	--3528
		x"43",	--3529
		x"41",	--3530
		x"12",	--3531
		x"12",	--3532
		x"83",	--3533
		x"4e",	--3534
		x"00",	--3535
		x"42",	--3536
		x"02",	--3537
		x"42",	--3538
		x"02",	--3539
		x"4e",	--3540
		x"4f",	--3541
		x"40",	--3542
		x"db",	--3543
		x"12",	--3544
		x"dd",	--3545
		x"9b",	--3546
		x"38",	--3547
		x"4a",	--3548
		x"5b",	--3549
		x"43",	--3550
		x"ff",	--3551
		x"3c",	--3552
		x"42",	--3553
		x"02",	--3554
		x"43",	--3555
		x"00",	--3556
		x"53",	--3557
		x"41",	--3558
		x"41",	--3559
		x"41",	--3560
		x"41",	--3561
		x"00",	--3562
		x"02",	--3563
		x"40",	--3564
		x"7f",	--3565
		x"02",	--3566
		x"41",	--3567
		x"50",	--3568
		x"00",	--3569
		x"41",	--3570
		x"00",	--3571
		x"12",	--3572
		x"db",	--3573
		x"41",	--3574
		x"41",	--3575
		x"00",	--3576
		x"02",	--3577
		x"41",	--3578
		x"00",	--3579
		x"02",	--3580
		x"41",	--3581
		x"52",	--3582
		x"41",	--3583
		x"00",	--3584
		x"12",	--3585
		x"db",	--3586
		x"41",	--3587
		x"4e",	--3588
		x"4f",	--3589
		x"02",	--3590
		x"40",	--3591
		x"7f",	--3592
		x"02",	--3593
		x"4d",	--3594
		x"4c",	--3595
		x"12",	--3596
		x"db",	--3597
		x"41",	--3598
		x"4f",	--3599
		x"02",	--3600
		x"4e",	--3601
		x"02",	--3602
		x"4c",	--3603
		x"4d",	--3604
		x"12",	--3605
		x"db",	--3606
		x"41",	--3607
		x"12",	--3608
		x"12",	--3609
		x"12",	--3610
		x"12",	--3611
		x"12",	--3612
		x"12",	--3613
		x"12",	--3614
		x"12",	--3615
		x"82",	--3616
		x"4f",	--3617
		x"4e",	--3618
		x"00",	--3619
		x"4d",	--3620
		x"41",	--3621
		x"00",	--3622
		x"41",	--3623
		x"00",	--3624
		x"4d",	--3625
		x"4d",	--3626
		x"10",	--3627
		x"44",	--3628
		x"4f",	--3629
		x"b0",	--3630
		x"00",	--3631
		x"24",	--3632
		x"40",	--3633
		x"00",	--3634
		x"00",	--3635
		x"4f",	--3636
		x"10",	--3637
		x"f3",	--3638
		x"24",	--3639
		x"40",	--3640
		x"00",	--3641
		x"3c",	--3642
		x"40",	--3643
		x"00",	--3644
		x"4e",	--3645
		x"00",	--3646
		x"41",	--3647
		x"53",	--3648
		x"3c",	--3649
		x"f0",	--3650
		x"00",	--3651
		x"24",	--3652
		x"40",	--3653
		x"00",	--3654
		x"00",	--3655
		x"3c",	--3656
		x"93",	--3657
		x"24",	--3658
		x"4d",	--3659
		x"00",	--3660
		x"41",	--3661
		x"53",	--3662
		x"3c",	--3663
		x"41",	--3664
		x"4c",	--3665
		x"10",	--3666
		x"11",	--3667
		x"10",	--3668
		x"11",	--3669
		x"4c",	--3670
		x"41",	--3671
		x"41",	--3672
		x"10",	--3673
		x"11",	--3674
		x"10",	--3675
		x"11",	--3676
		x"4c",	--3677
		x"86",	--3678
		x"77",	--3679
		x"4f",	--3680
		x"10",	--3681
		x"4e",	--3682
		x"00",	--3683
		x"f2",	--3684
		x"24",	--3685
		x"45",	--3686
		x"3c",	--3687
		x"43",	--3688
		x"4f",	--3689
		x"b0",	--3690
		x"00",	--3691
		x"20",	--3692
		x"41",	--3693
		x"00",	--3694
		x"53",	--3695
		x"53",	--3696
		x"93",	--3697
		x"00",	--3698
		x"23",	--3699
		x"81",	--3700
		x"00",	--3701
		x"9a",	--3702
		x"28",	--3703
		x"8a",	--3704
		x"3c",	--3705
		x"43",	--3706
		x"b3",	--3707
		x"00",	--3708
		x"24",	--3709
		x"95",	--3710
		x"28",	--3711
		x"85",	--3712
		x"3c",	--3713
		x"43",	--3714
		x"4d",	--3715
		x"9d",	--3716
		x"2c",	--3717
		x"47",	--3718
		x"93",	--3719
		x"38",	--3720
		x"40",	--3721
		x"00",	--3722
		x"00",	--3723
		x"43",	--3724
		x"43",	--3725
		x"3c",	--3726
		x"41",	--3727
		x"56",	--3728
		x"4f",	--3729
		x"11",	--3730
		x"53",	--3731
		x"12",	--3732
		x"3c",	--3733
		x"43",	--3734
		x"9a",	--3735
		x"3b",	--3736
		x"4a",	--3737
		x"40",	--3738
		x"00",	--3739
		x"00",	--3740
		x"8b",	--3741
		x"3c",	--3742
		x"41",	--3743
		x"00",	--3744
		x"11",	--3745
		x"12",	--3746
		x"53",	--3747
		x"45",	--3748
		x"5b",	--3749
		x"99",	--3750
		x"2b",	--3751
		x"3c",	--3752
		x"43",	--3753
		x"43",	--3754
		x"3c",	--3755
		x"53",	--3756
		x"41",	--3757
		x"56",	--3758
		x"4f",	--3759
		x"11",	--3760
		x"53",	--3761
		x"12",	--3762
		x"9a",	--3763
		x"3b",	--3764
		x"b3",	--3765
		x"00",	--3766
		x"24",	--3767
		x"44",	--3768
		x"3c",	--3769
		x"41",	--3770
		x"00",	--3771
		x"8b",	--3772
		x"3c",	--3773
		x"40",	--3774
		x"00",	--3775
		x"12",	--3776
		x"53",	--3777
		x"93",	--3778
		x"23",	--3779
		x"44",	--3780
		x"54",	--3781
		x"3f",	--3782
		x"53",	--3783
		x"11",	--3784
		x"12",	--3785
		x"53",	--3786
		x"4a",	--3787
		x"5b",	--3788
		x"4f",	--3789
		x"93",	--3790
		x"24",	--3791
		x"93",	--3792
		x"23",	--3793
		x"3c",	--3794
		x"40",	--3795
		x"00",	--3796
		x"12",	--3797
		x"53",	--3798
		x"99",	--3799
		x"2b",	--3800
		x"4b",	--3801
		x"52",	--3802
		x"41",	--3803
		x"41",	--3804
		x"41",	--3805
		x"41",	--3806
		x"41",	--3807
		x"41",	--3808
		x"41",	--3809
		x"41",	--3810
		x"41",	--3811
		x"12",	--3812
		x"12",	--3813
		x"12",	--3814
		x"12",	--3815
		x"12",	--3816
		x"12",	--3817
		x"12",	--3818
		x"12",	--3819
		x"50",	--3820
		x"ff",	--3821
		x"4f",	--3822
		x"00",	--3823
		x"4e",	--3824
		x"4d",	--3825
		x"4e",	--3826
		x"00",	--3827
		x"43",	--3828
		x"00",	--3829
		x"43",	--3830
		x"00",	--3831
		x"43",	--3832
		x"00",	--3833
		x"43",	--3834
		x"00",	--3835
		x"43",	--3836
		x"00",	--3837
		x"43",	--3838
		x"00",	--3839
		x"43",	--3840
		x"43",	--3841
		x"00",	--3842
		x"41",	--3843
		x"50",	--3844
		x"00",	--3845
		x"4e",	--3846
		x"00",	--3847
		x"40",	--3848
		x"e4",	--3849
		x"46",	--3850
		x"53",	--3851
		x"4f",	--3852
		x"00",	--3853
		x"93",	--3854
		x"20",	--3855
		x"90",	--3856
		x"00",	--3857
		x"20",	--3858
		x"43",	--3859
		x"00",	--3860
		x"43",	--3861
		x"00",	--3862
		x"46",	--3863
		x"00",	--3864
		x"43",	--3865
		x"00",	--3866
		x"43",	--3867
		x"00",	--3868
		x"43",	--3869
		x"00",	--3870
		x"43",	--3871
		x"00",	--3872
		x"43",	--3873
		x"00",	--3874
		x"40",	--3875
		x"e4",	--3876
		x"47",	--3877
		x"11",	--3878
		x"4e",	--3879
		x"12",	--3880
		x"00",	--3881
		x"53",	--3882
		x"00",	--3883
		x"40",	--3884
		x"e4",	--3885
		x"90",	--3886
		x"00",	--3887
		x"24",	--3888
		x"90",	--3889
		x"00",	--3890
		x"34",	--3891
		x"90",	--3892
		x"00",	--3893
		x"24",	--3894
		x"90",	--3895
		x"00",	--3896
		x"34",	--3897
		x"90",	--3898
		x"00",	--3899
		x"24",	--3900
		x"90",	--3901
		x"00",	--3902
		x"34",	--3903
		x"90",	--3904
		x"00",	--3905
		x"24",	--3906
		x"90",	--3907
		x"00",	--3908
		x"27",	--3909
		x"90",	--3910
		x"00",	--3911
		x"20",	--3912
		x"3c",	--3913
		x"90",	--3914
		x"00",	--3915
		x"24",	--3916
		x"90",	--3917
		x"00",	--3918
		x"24",	--3919
		x"90",	--3920
		x"00",	--3921
		x"20",	--3922
		x"3c",	--3923
		x"90",	--3924
		x"00",	--3925
		x"38",	--3926
		x"90",	--3927
		x"00",	--3928
		x"20",	--3929
		x"3c",	--3930
		x"90",	--3931
		x"00",	--3932
		x"24",	--3933
		x"90",	--3934
		x"00",	--3935
		x"34",	--3936
		x"90",	--3937
		x"00",	--3938
		x"24",	--3939
		x"90",	--3940
		x"00",	--3941
		x"24",	--3942
		x"90",	--3943
		x"00",	--3944
		x"20",	--3945
		x"3c",	--3946
		x"90",	--3947
		x"00",	--3948
		x"24",	--3949
		x"90",	--3950
		x"00",	--3951
		x"34",	--3952
		x"90",	--3953
		x"00",	--3954
		x"20",	--3955
		x"3c",	--3956
		x"90",	--3957
		x"00",	--3958
		x"24",	--3959
		x"90",	--3960
		x"00",	--3961
		x"24",	--3962
		x"41",	--3963
		x"00",	--3964
		x"41",	--3965
		x"00",	--3966
		x"89",	--3967
		x"40",	--3968
		x"e4",	--3969
		x"42",	--3970
		x"00",	--3971
		x"3c",	--3972
		x"d2",	--3973
		x"00",	--3974
		x"40",	--3975
		x"e4",	--3976
		x"41",	--3977
		x"f3",	--3978
		x"41",	--3979
		x"24",	--3980
		x"f0",	--3981
		x"ff",	--3982
		x"d3",	--3983
		x"3c",	--3984
		x"d3",	--3985
		x"4e",	--3986
		x"00",	--3987
		x"40",	--3988
		x"e4",	--3989
		x"d0",	--3990
		x"00",	--3991
		x"00",	--3992
		x"40",	--3993
		x"e4",	--3994
		x"40",	--3995
		x"00",	--3996
		x"00",	--3997
		x"40",	--3998
		x"e4",	--3999
		x"90",	--4000
		x"00",	--4001
		x"00",	--4002
		x"20",	--4003
		x"40",	--4004
		x"e4",	--4005
		x"40",	--4006
		x"00",	--4007
		x"00",	--4008
		x"40",	--4009
		x"e4",	--4010
		x"93",	--4011
		x"00",	--4012
		x"24",	--4013
		x"40",	--4014
		x"e4",	--4015
		x"43",	--4016
		x"00",	--4017
		x"40",	--4018
		x"e4",	--4019
		x"45",	--4020
		x"53",	--4021
		x"45",	--4022
		x"93",	--4023
		x"38",	--4024
		x"4a",	--4025
		x"00",	--4026
		x"3c",	--4027
		x"93",	--4028
		x"00",	--4029
		x"24",	--4030
		x"40",	--4031
		x"e4",	--4032
		x"d0",	--4033
		x"00",	--4034
		x"00",	--4035
		x"e3",	--4036
		x"4a",	--4037
		x"00",	--4038
		x"53",	--4039
		x"00",	--4040
		x"4e",	--4041
		x"3c",	--4042
		x"93",	--4043
		x"00",	--4044
		x"20",	--4045
		x"93",	--4046
		x"00",	--4047
		x"20",	--4048
		x"41",	--4049
		x"f0",	--4050
		x"00",	--4051
		x"43",	--4052
		x"24",	--4053
		x"43",	--4054
		x"4e",	--4055
		x"11",	--4056
		x"43",	--4057
		x"10",	--4058
		x"41",	--4059
		x"f0",	--4060
		x"00",	--4061
		x"de",	--4062
		x"4a",	--4063
		x"00",	--4064
		x"40",	--4065
		x"e4",	--4066
		x"41",	--4067
		x"00",	--4068
		x"5a",	--4069
		x"4a",	--4070
		x"5c",	--4071
		x"5c",	--4072
		x"5c",	--4073
		x"4a",	--4074
		x"00",	--4075
		x"50",	--4076
		x"ff",	--4077
		x"00",	--4078
		x"11",	--4079
		x"5e",	--4080
		x"00",	--4081
		x"43",	--4082
		x"00",	--4083
		x"40",	--4084
		x"e4",	--4085
		x"45",	--4086
		x"53",	--4087
		x"45",	--4088
		x"93",	--4089
		x"00",	--4090
		x"20",	--4091
		x"93",	--4092
		x"00",	--4093
		x"27",	--4094
		x"4e",	--4095
		x"00",	--4096
		x"43",	--4097
		x"00",	--4098
		x"41",	--4099
		x"52",	--4100
		x"3c",	--4101
		x"45",	--4102
		x"53",	--4103
		x"45",	--4104
		x"93",	--4105
		x"00",	--4106
		x"24",	--4107
		x"d2",	--4108
		x"00",	--4109
		x"41",	--4110
		x"00",	--4111
		x"4f",	--4112
		x"00",	--4113
		x"3c",	--4114
		x"93",	--4115
		x"00",	--4116
		x"24",	--4117
		x"41",	--4118
		x"00",	--4119
		x"00",	--4120
		x"93",	--4121
		x"20",	--4122
		x"40",	--4123
		x"e9",	--4124
		x"12",	--4125
		x"00",	--4126
		x"12",	--4127
		x"00",	--4128
		x"41",	--4129
		x"00",	--4130
		x"41",	--4131
		x"00",	--4132
		x"12",	--4133
		x"dc",	--4134
		x"52",	--4135
		x"5f",	--4136
		x"00",	--4137
		x"47",	--4138
		x"40",	--4139
		x"e4",	--4140
		x"45",	--4141
		x"53",	--4142
		x"45",	--4143
		x"49",	--4144
		x"00",	--4145
		x"43",	--4146
		x"93",	--4147
		x"20",	--4148
		x"43",	--4149
		x"5e",	--4150
		x"5e",	--4151
		x"5e",	--4152
		x"41",	--4153
		x"f0",	--4154
		x"ff",	--4155
		x"de",	--4156
		x"4a",	--4157
		x"00",	--4158
		x"47",	--4159
		x"40",	--4160
		x"00",	--4161
		x"00",	--4162
		x"3c",	--4163
		x"d3",	--4164
		x"00",	--4165
		x"3c",	--4166
		x"d2",	--4167
		x"00",	--4168
		x"40",	--4169
		x"00",	--4170
		x"00",	--4171
		x"3c",	--4172
		x"40",	--4173
		x"00",	--4174
		x"00",	--4175
		x"41",	--4176
		x"b3",	--4177
		x"24",	--4178
		x"45",	--4179
		x"52",	--4180
		x"45",	--4181
		x"45",	--4182
		x"00",	--4183
		x"45",	--4184
		x"00",	--4185
		x"45",	--4186
		x"00",	--4187
		x"48",	--4188
		x"00",	--4189
		x"47",	--4190
		x"00",	--4191
		x"46",	--4192
		x"00",	--4193
		x"4b",	--4194
		x"00",	--4195
		x"43",	--4196
		x"00",	--4197
		x"93",	--4198
		x"20",	--4199
		x"93",	--4200
		x"20",	--4201
		x"93",	--4202
		x"20",	--4203
		x"93",	--4204
		x"24",	--4205
		x"43",	--4206
		x"00",	--4207
		x"5b",	--4208
		x"43",	--4209
		x"6b",	--4210
		x"4b",	--4211
		x"00",	--4212
		x"4c",	--4213
		x"3c",	--4214
		x"f3",	--4215
		x"45",	--4216
		x"24",	--4217
		x"52",	--4218
		x"45",	--4219
		x"45",	--4220
		x"00",	--4221
		x"48",	--4222
		x"00",	--4223
		x"4b",	--4224
		x"00",	--4225
		x"43",	--4226
		x"00",	--4227
		x"93",	--4228
		x"20",	--4229
		x"3c",	--4230
		x"53",	--4231
		x"45",	--4232
		x"4b",	--4233
		x"00",	--4234
		x"43",	--4235
		x"00",	--4236
		x"93",	--4237
		x"24",	--4238
		x"43",	--4239
		x"00",	--4240
		x"5b",	--4241
		x"43",	--4242
		x"6b",	--4243
		x"4b",	--4244
		x"00",	--4245
		x"47",	--4246
		x"b2",	--4247
		x"00",	--4248
		x"24",	--4249
		x"93",	--4250
		x"00",	--4251
		x"20",	--4252
		x"41",	--4253
		x"90",	--4254
		x"00",	--4255
		x"00",	--4256
		x"20",	--4257
		x"d0",	--4258
		x"00",	--4259
		x"3c",	--4260
		x"92",	--4261
		x"00",	--4262
		x"20",	--4263
		x"d0",	--4264
		x"00",	--4265
		x"48",	--4266
		x"00",	--4267
		x"41",	--4268
		x"b2",	--4269
		x"24",	--4270
		x"93",	--4271
		x"00",	--4272
		x"24",	--4273
		x"40",	--4274
		x"00",	--4275
		x"00",	--4276
		x"b3",	--4277
		x"24",	--4278
		x"e3",	--4279
		x"00",	--4280
		x"e3",	--4281
		x"00",	--4282
		x"e3",	--4283
		x"00",	--4284
		x"e3",	--4285
		x"00",	--4286
		x"53",	--4287
		x"00",	--4288
		x"63",	--4289
		x"00",	--4290
		x"63",	--4291
		x"00",	--4292
		x"63",	--4293
		x"00",	--4294
		x"3c",	--4295
		x"b3",	--4296
		x"24",	--4297
		x"41",	--4298
		x"00",	--4299
		x"41",	--4300
		x"00",	--4301
		x"e3",	--4302
		x"e3",	--4303
		x"4a",	--4304
		x"4b",	--4305
		x"53",	--4306
		x"63",	--4307
		x"4e",	--4308
		x"00",	--4309
		x"4f",	--4310
		x"00",	--4311
		x"3c",	--4312
		x"41",	--4313
		x"00",	--4314
		x"e3",	--4315
		x"53",	--4316
		x"4a",	--4317
		x"00",	--4318
		x"43",	--4319
		x"00",	--4320
		x"b3",	--4321
		x"24",	--4322
		x"41",	--4323
		x"00",	--4324
		x"41",	--4325
		x"00",	--4326
		x"00",	--4327
		x"41",	--4328
		x"00",	--4329
		x"41",	--4330
		x"00",	--4331
		x"41",	--4332
		x"50",	--4333
		x"00",	--4334
		x"46",	--4335
		x"41",	--4336
		x"00",	--4337
		x"00",	--4338
		x"41",	--4339
		x"00",	--4340
		x"10",	--4341
		x"11",	--4342
		x"10",	--4343
		x"11",	--4344
		x"4b",	--4345
		x"00",	--4346
		x"4b",	--4347
		x"00",	--4348
		x"4b",	--4349
		x"00",	--4350
		x"12",	--4351
		x"00",	--4352
		x"12",	--4353
		x"00",	--4354
		x"12",	--4355
		x"00",	--4356
		x"12",	--4357
		x"00",	--4358
		x"49",	--4359
		x"41",	--4360
		x"00",	--4361
		x"48",	--4362
		x"44",	--4363
		x"12",	--4364
		x"e5",	--4365
		x"52",	--4366
		x"4c",	--4367
		x"90",	--4368
		x"00",	--4369
		x"34",	--4370
		x"50",	--4371
		x"00",	--4372
		x"4b",	--4373
		x"00",	--4374
		x"3c",	--4375
		x"4c",	--4376
		x"b3",	--4377
		x"00",	--4378
		x"24",	--4379
		x"40",	--4380
		x"00",	--4381
		x"3c",	--4382
		x"40",	--4383
		x"00",	--4384
		x"5b",	--4385
		x"4a",	--4386
		x"00",	--4387
		x"47",	--4388
		x"53",	--4389
		x"12",	--4390
		x"00",	--4391
		x"12",	--4392
		x"00",	--4393
		x"12",	--4394
		x"00",	--4395
		x"12",	--4396
		x"00",	--4397
		x"49",	--4398
		x"41",	--4399
		x"00",	--4400
		x"48",	--4401
		x"44",	--4402
		x"12",	--4403
		x"e5",	--4404
		x"52",	--4405
		x"4c",	--4406
		x"4d",	--4407
		x"00",	--4408
		x"4e",	--4409
		x"4f",	--4410
		x"53",	--4411
		x"93",	--4412
		x"23",	--4413
		x"93",	--4414
		x"23",	--4415
		x"93",	--4416
		x"23",	--4417
		x"93",	--4418
		x"23",	--4419
		x"43",	--4420
		x"00",	--4421
		x"43",	--4422
		x"00",	--4423
		x"43",	--4424
		x"00",	--4425
		x"43",	--4426
		x"00",	--4427
		x"3c",	--4428
		x"b3",	--4429
		x"24",	--4430
		x"41",	--4431
		x"00",	--4432
		x"41",	--4433
		x"00",	--4434
		x"41",	--4435
		x"50",	--4436
		x"00",	--4437
		x"41",	--4438
		x"00",	--4439
		x"10",	--4440
		x"11",	--4441
		x"10",	--4442
		x"11",	--4443
		x"41",	--4444
		x"00",	--4445
		x"49",	--4446
		x"44",	--4447
		x"47",	--4448
		x"12",	--4449
		x"e4",	--4450
		x"4e",	--4451
		x"90",	--4452
		x"00",	--4453
		x"34",	--4454
		x"50",	--4455
		x"00",	--4456
		x"4b",	--4457
		x"00",	--4458
		x"3c",	--4459
		x"4e",	--4460
		x"b3",	--4461
		x"00",	--4462
		x"24",	--4463
		x"40",	--4464
		x"00",	--4465
		x"3c",	--4466
		x"40",	--4467
		x"00",	--4468
		x"5b",	--4469
		x"4a",	--4470
		x"00",	--4471
		x"48",	--4472
		x"53",	--4473
		x"41",	--4474
		x"00",	--4475
		x"49",	--4476
		x"44",	--4477
		x"47",	--4478
		x"12",	--4479
		x"e4",	--4480
		x"4e",	--4481
		x"4f",	--4482
		x"53",	--4483
		x"93",	--4484
		x"23",	--4485
		x"93",	--4486
		x"23",	--4487
		x"43",	--4488
		x"00",	--4489
		x"43",	--4490
		x"00",	--4491
		x"3c",	--4492
		x"41",	--4493
		x"00",	--4494
		x"41",	--4495
		x"50",	--4496
		x"00",	--4497
		x"41",	--4498
		x"00",	--4499
		x"47",	--4500
		x"12",	--4501
		x"e5",	--4502
		x"4f",	--4503
		x"90",	--4504
		x"00",	--4505
		x"34",	--4506
		x"50",	--4507
		x"00",	--4508
		x"4d",	--4509
		x"00",	--4510
		x"3c",	--4511
		x"4f",	--4512
		x"b3",	--4513
		x"00",	--4514
		x"24",	--4515
		x"40",	--4516
		x"00",	--4517
		x"3c",	--4518
		x"40",	--4519
		x"00",	--4520
		x"5d",	--4521
		x"4c",	--4522
		x"00",	--4523
		x"48",	--4524
		x"53",	--4525
		x"41",	--4526
		x"00",	--4527
		x"47",	--4528
		x"12",	--4529
		x"e5",	--4530
		x"4f",	--4531
		x"53",	--4532
		x"93",	--4533
		x"23",	--4534
		x"43",	--4535
		x"00",	--4536
		x"90",	--4537
		x"00",	--4538
		x"00",	--4539
		x"24",	--4540
		x"43",	--4541
		x"00",	--4542
		x"93",	--4543
		x"00",	--4544
		x"24",	--4545
		x"41",	--4546
		x"50",	--4547
		x"00",	--4548
		x"4f",	--4549
		x"00",	--4550
		x"41",	--4551
		x"00",	--4552
		x"10",	--4553
		x"11",	--4554
		x"10",	--4555
		x"11",	--4556
		x"4a",	--4557
		x"00",	--4558
		x"46",	--4559
		x"00",	--4560
		x"46",	--4561
		x"10",	--4562
		x"11",	--4563
		x"10",	--4564
		x"11",	--4565
		x"4a",	--4566
		x"00",	--4567
		x"41",	--4568
		x"00",	--4569
		x"41",	--4570
		x"00",	--4571
		x"81",	--4572
		x"00",	--4573
		x"71",	--4574
		x"00",	--4575
		x"83",	--4576
		x"91",	--4577
		x"00",	--4578
		x"2c",	--4579
		x"d3",	--4580
		x"00",	--4581
		x"41",	--4582
		x"00",	--4583
		x"8c",	--4584
		x"4e",	--4585
		x"00",	--4586
		x"3c",	--4587
		x"93",	--4588
		x"00",	--4589
		x"24",	--4590
		x"41",	--4591
		x"00",	--4592
		x"00",	--4593
		x"12",	--4594
		x"00",	--4595
		x"12",	--4596
		x"00",	--4597
		x"41",	--4598
		x"00",	--4599
		x"46",	--4600
		x"53",	--4601
		x"41",	--4602
		x"00",	--4603
		x"12",	--4604
		x"dc",	--4605
		x"52",	--4606
		x"5f",	--4607
		x"00",	--4608
		x"3c",	--4609
		x"49",	--4610
		x"11",	--4611
		x"12",	--4612
		x"00",	--4613
		x"49",	--4614
		x"58",	--4615
		x"91",	--4616
		x"00",	--4617
		x"2b",	--4618
		x"49",	--4619
		x"00",	--4620
		x"4e",	--4621
		x"00",	--4622
		x"43",	--4623
		x"3c",	--4624
		x"41",	--4625
		x"00",	--4626
		x"00",	--4627
		x"43",	--4628
		x"00",	--4629
		x"43",	--4630
		x"00",	--4631
		x"3c",	--4632
		x"4e",	--4633
		x"43",	--4634
		x"00",	--4635
		x"43",	--4636
		x"00",	--4637
		x"43",	--4638
		x"41",	--4639
		x"00",	--4640
		x"46",	--4641
		x"93",	--4642
		x"24",	--4643
		x"40",	--4644
		x"de",	--4645
		x"41",	--4646
		x"00",	--4647
		x"50",	--4648
		x"00",	--4649
		x"41",	--4650
		x"41",	--4651
		x"41",	--4652
		x"41",	--4653
		x"41",	--4654
		x"41",	--4655
		x"41",	--4656
		x"41",	--4657
		x"41",	--4658
		x"43",	--4659
		x"93",	--4660
		x"34",	--4661
		x"40",	--4662
		x"00",	--4663
		x"e3",	--4664
		x"53",	--4665
		x"93",	--4666
		x"34",	--4667
		x"e3",	--4668
		x"e3",	--4669
		x"53",	--4670
		x"12",	--4671
		x"12",	--4672
		x"e5",	--4673
		x"41",	--4674
		x"b3",	--4675
		x"24",	--4676
		x"e3",	--4677
		x"53",	--4678
		x"b3",	--4679
		x"24",	--4680
		x"e3",	--4681
		x"53",	--4682
		x"41",	--4683
		x"12",	--4684
		x"e4",	--4685
		x"4e",	--4686
		x"41",	--4687
		x"12",	--4688
		x"12",	--4689
		x"12",	--4690
		x"40",	--4691
		x"00",	--4692
		x"4c",	--4693
		x"4d",	--4694
		x"43",	--4695
		x"43",	--4696
		x"5e",	--4697
		x"6f",	--4698
		x"6c",	--4699
		x"6d",	--4700
		x"9b",	--4701
		x"28",	--4702
		x"20",	--4703
		x"9a",	--4704
		x"28",	--4705
		x"8a",	--4706
		x"7b",	--4707
		x"d3",	--4708
		x"83",	--4709
		x"23",	--4710
		x"41",	--4711
		x"41",	--4712
		x"41",	--4713
		x"41",	--4714
		x"12",	--4715
		x"e4",	--4716
		x"4c",	--4717
		x"4d",	--4718
		x"41",	--4719
		x"12",	--4720
		x"43",	--4721
		x"93",	--4722
		x"34",	--4723
		x"40",	--4724
		x"00",	--4725
		x"e3",	--4726
		x"e3",	--4727
		x"53",	--4728
		x"63",	--4729
		x"93",	--4730
		x"34",	--4731
		x"e3",	--4732
		x"e3",	--4733
		x"e3",	--4734
		x"53",	--4735
		x"63",	--4736
		x"12",	--4737
		x"e4",	--4738
		x"b3",	--4739
		x"24",	--4740
		x"e3",	--4741
		x"e3",	--4742
		x"53",	--4743
		x"63",	--4744
		x"b3",	--4745
		x"24",	--4746
		x"e3",	--4747
		x"e3",	--4748
		x"53",	--4749
		x"63",	--4750
		x"41",	--4751
		x"41",	--4752
		x"12",	--4753
		x"e4",	--4754
		x"4c",	--4755
		x"4d",	--4756
		x"41",	--4757
		x"40",	--4758
		x"00",	--4759
		x"4e",	--4760
		x"43",	--4761
		x"5f",	--4762
		x"6e",	--4763
		x"9d",	--4764
		x"28",	--4765
		x"8d",	--4766
		x"d3",	--4767
		x"83",	--4768
		x"23",	--4769
		x"41",	--4770
		x"12",	--4771
		x"e5",	--4772
		x"4e",	--4773
		x"41",	--4774
		x"12",	--4775
		x"12",	--4776
		x"12",	--4777
		x"12",	--4778
		x"12",	--4779
		x"00",	--4780
		x"48",	--4781
		x"49",	--4782
		x"4a",	--4783
		x"4b",	--4784
		x"43",	--4785
		x"43",	--4786
		x"43",	--4787
		x"43",	--4788
		x"5c",	--4789
		x"6d",	--4790
		x"6e",	--4791
		x"6f",	--4792
		x"68",	--4793
		x"69",	--4794
		x"6a",	--4795
		x"6b",	--4796
		x"97",	--4797
		x"28",	--4798
		x"20",	--4799
		x"96",	--4800
		x"28",	--4801
		x"20",	--4802
		x"95",	--4803
		x"28",	--4804
		x"20",	--4805
		x"94",	--4806
		x"28",	--4807
		x"84",	--4808
		x"75",	--4809
		x"76",	--4810
		x"77",	--4811
		x"d3",	--4812
		x"83",	--4813
		x"00",	--4814
		x"23",	--4815
		x"53",	--4816
		x"41",	--4817
		x"41",	--4818
		x"41",	--4819
		x"41",	--4820
		x"41",	--4821
		x"12",	--4822
		x"12",	--4823
		x"12",	--4824
		x"12",	--4825
		x"41",	--4826
		x"00",	--4827
		x"41",	--4828
		x"00",	--4829
		x"41",	--4830
		x"00",	--4831
		x"41",	--4832
		x"00",	--4833
		x"12",	--4834
		x"e5",	--4835
		x"41",	--4836
		x"41",	--4837
		x"41",	--4838
		x"41",	--4839
		x"41",	--4840
		x"12",	--4841
		x"12",	--4842
		x"12",	--4843
		x"12",	--4844
		x"41",	--4845
		x"00",	--4846
		x"41",	--4847
		x"00",	--4848
		x"41",	--4849
		x"00",	--4850
		x"41",	--4851
		x"00",	--4852
		x"12",	--4853
		x"e5",	--4854
		x"48",	--4855
		x"49",	--4856
		x"4a",	--4857
		x"4b",	--4858
		x"41",	--4859
		x"41",	--4860
		x"41",	--4861
		x"41",	--4862
		x"41",	--4863
		x"12",	--4864
		x"12",	--4865
		x"12",	--4866
		x"12",	--4867
		x"12",	--4868
		x"41",	--4869
		x"00",	--4870
		x"41",	--4871
		x"00",	--4872
		x"41",	--4873
		x"00",	--4874
		x"41",	--4875
		x"00",	--4876
		x"12",	--4877
		x"e5",	--4878
		x"41",	--4879
		x"00",	--4880
		x"48",	--4881
		x"00",	--4882
		x"49",	--4883
		x"00",	--4884
		x"4a",	--4885
		x"00",	--4886
		x"4b",	--4887
		x"00",	--4888
		x"41",	--4889
		x"41",	--4890
		x"41",	--4891
		x"41",	--4892
		x"41",	--4893
		x"41",	--4894
		x"13",	--4895
		x"d0",	--4896
		x"00",	--4897
		x"3f",	--4898
		x"61",	--4899
		x"74",	--4900
		x"6e",	--4901
		x"20",	--4902
		x"6f",	--4903
		x"20",	--4904
		x"20",	--4905
		x"65",	--4906
		x"20",	--4907
		x"62",	--4908
		x"6e",	--4909
		x"66",	--4910
		x"6c",	--4911
		x"0d",	--4912
		x"00",	--4913
		x"65",	--4914
		x"73",	--4915
		x"6f",	--4916
		x"6c",	--4917
		x"20",	--4918
		x"6f",	--4919
		x"20",	--4920
		x"65",	--4921
		x"20",	--4922
		x"68",	--4923
		x"74",	--4924
		x"0a",	--4925
		x"53",	--4926
		x"6f",	--4927
		x"0d",	--4928
		x"00",	--4929
		x"72",	--4930
		x"6f",	--4931
		x"3a",	--4932
		x"6d",	--4933
		x"73",	--4934
		x"69",	--4935
		x"67",	--4936
		x"61",	--4937
		x"67",	--4938
		x"6d",	--4939
		x"6e",	--4940
		x"0d",	--4941
		x"00",	--4942
		x"6f",	--4943
		x"72",	--4944
		x"63",	--4945
		x"20",	--4946
		x"73",	--4947
		x"67",	--4948
		x"3a",	--4949
		x"0a",	--4950
		x"09",	--4951
		x"73",	--4952
		x"4c",	--4953
		x"46",	--4954
		x"20",	--4955
		x"49",	--4956
		x"48",	--4957
		x"20",	--4958
		x"54",	--4959
		x"4d",	--4960
		x"4f",	--4961
		x"54",	--4962
		x"0d",	--4963
		x"00",	--4964
		x"64",	--4965
		x"25",	--4966
		x"0d",	--4967
		x"00",	--4968
		x"6c",	--4969
		x"20",	--4970
		x"6c",	--4971
		x"00",	--4972
		x"73",	--4973
		x"0a",	--4974
		x"25",	--4975
		x"20",	--4976
		x"64",	--4977
		x"0a",	--4978
		x"00",	--4979
		x"c5",	--4980
		x"c5",	--4981
		x"c6",	--4982
		x"c6",	--4983
		x"c6",	--4984
		x"c6",	--4985
		x"c5",	--4986
		x"c5",	--4987
		x"0a",	--4988
		x"3d",	--4989
		x"3d",	--4990
		x"3d",	--4991
		x"4d",	--4992
		x"72",	--4993
		x"65",	--4994
		x"20",	--4995
		x"43",	--4996
		x"20",	--4997
		x"3d",	--4998
		x"3d",	--4999
		x"3d",	--5000
		x"0a",	--5001
		x"69",	--5002
		x"74",	--5003
		x"72",	--5004
		x"63",	--5005
		x"69",	--5006
		x"65",	--5007
		x"6d",	--5008
		x"64",	--5009
		x"00",	--5010
		x"72",	--5011
		x"74",	--5012
		x"00",	--5013
		x"65",	--5014
		x"64",	--5015
		x"70",	--5016
		x"6d",	--5017
		x"65",	--5018
		x"63",	--5019
		x"64",	--5020
		x"72",	--5021
		x"73",	--5022
		x"65",	--5023
		x"64",	--5024
		x"63",	--5025
		x"6e",	--5026
		x"72",	--5027
		x"6c",	--5028
		x"65",	--5029
		x"00",	--5030
		x"70",	--5031
		x"65",	--5032
		x"20",	--5033
		x"6f",	--5034
		x"66",	--5035
		x"67",	--5036
		x"72",	--5037
		x"74",	--5038
		x"6f",	--5039
		x"00",	--5040
		x"6f",	--5041
		x"74",	--5042
		x"6f",	--5043
		x"64",	--5044
		x"72",	--5045
		x"0d",	--5046
		x"00",	--5047
		x"20",	--5048
		x"00",	--5049
		x"63",	--5050
		x"00",	--5051
		x"72",	--5052
		x"74",	--5053
		x"0a",	--5054
		x"00",	--5055
		x"72",	--5056
		x"6f",	--5057
		x"3a",	--5058
		x"6d",	--5059
		x"73",	--5060
		x"69",	--5061
		x"67",	--5062
		x"61",	--5063
		x"67",	--5064
		x"6d",	--5065
		x"6e",	--5066
		x"0d",	--5067
		x"00",	--5068
		x"6f",	--5069
		x"72",	--5070
		x"63",	--5071
		x"20",	--5072
		x"73",	--5073
		x"67",	--5074
		x"3a",	--5075
		x"0a",	--5076
		x"09",	--5077
		x"73",	--5078
		x"52",	--5079
		x"47",	--5080
		x"53",	--5081
		x"45",	--5082
		x"20",	--5083
		x"41",	--5084
		x"55",	--5085
		x"0d",	--5086
		x"00",	--5087
		x"3d",	--5088
		x"64",	--5089
		x"76",	--5090
		x"25",	--5091
		x"0d",	--5092
		x"00",	--5093
		x"25",	--5094
		x"20",	--5095
		x"45",	--5096
		x"49",	--5097
		x"54",	--5098
		x"52",	--5099
		x"0a",	--5100
		x"72",	--5101
		x"61",	--5102
		x"0a",	--5103
		x"00",	--5104
		x"63",	--5105
		x"69",	--5106
		x"20",	--5107
		x"6f",	--5108
		x"20",	--5109
		x"20",	--5110
		x"75",	--5111
		x"62",	--5112
		x"72",	--5113
		x"0a",	--5114
		x"25",	--5115
		x"20",	--5116
		x"73",	--5117
		x"0a",	--5118
		x"25",	--5119
		x"3a",	--5120
		x"6e",	--5121
		x"20",	--5122
		x"75",	--5123
		x"68",	--5124
		x"63",	--5125
		x"6d",	--5126
		x"61",	--5127
		x"64",	--5128
		x"0a",	--5129
		x"00",	--5130
		x"cd",	--5131
		x"cd",	--5132
		x"cd",	--5133
		x"cd",	--5134
		x"cd",	--5135
		x"cd",	--5136
		x"cd",	--5137
		x"cd",	--5138
		x"cd",	--5139
		x"cd",	--5140
		x"cd",	--5141
		x"cd",	--5142
		x"cd",	--5143
		x"cd",	--5144
		x"cd",	--5145
		x"cd",	--5146
		x"cd",	--5147
		x"cd",	--5148
		x"cd",	--5149
		x"cd",	--5150
		x"cd",	--5151
		x"cd",	--5152
		x"cd",	--5153
		x"cd",	--5154
		x"cd",	--5155
		x"cd",	--5156
		x"cd",	--5157
		x"cd",	--5158
		x"cd",	--5159
		x"cd",	--5160
		x"cd",	--5161
		x"cd",	--5162
		x"cd",	--5163
		x"cd",	--5164
		x"cd",	--5165
		x"cd",	--5166
		x"cd",	--5167
		x"cd",	--5168
		x"cd",	--5169
		x"cd",	--5170
		x"cd",	--5171
		x"cd",	--5172
		x"cd",	--5173
		x"cd",	--5174
		x"cd",	--5175
		x"cd",	--5176
		x"cd",	--5177
		x"cd",	--5178
		x"cd",	--5179
		x"cd",	--5180
		x"cd",	--5181
		x"cd",	--5182
		x"cd",	--5183
		x"cd",	--5184
		x"cd",	--5185
		x"cd",	--5186
		x"cd",	--5187
		x"cd",	--5188
		x"cd",	--5189
		x"cd",	--5190
		x"cd",	--5191
		x"cd",	--5192
		x"cd",	--5193
		x"cd",	--5194
		x"cd",	--5195
		x"cd",	--5196
		x"cd",	--5197
		x"cd",	--5198
		x"cd",	--5199
		x"cd",	--5200
		x"cd",	--5201
		x"cd",	--5202
		x"cd",	--5203
		x"cd",	--5204
		x"cd",	--5205
		x"cd",	--5206
		x"cd",	--5207
		x"cd",	--5208
		x"cd",	--5209
		x"cd",	--5210
		x"cd",	--5211
		x"cd",	--5212
		x"cd",	--5213
		x"cd",	--5214
		x"31",	--5215
		x"33",	--5216
		x"35",	--5217
		x"37",	--5218
		x"39",	--5219
		x"62",	--5220
		x"64",	--5221
		x"66",	--5222
		x"00",	--5223
		x"00",	--5224
		x"00",	--5225
		x"00",	--5226
		x"00",	--5227
		x"01",	--5228
		x"02",	--5229
		x"03",	--5230
		x"03",	--5231
		x"04",	--5232
		x"04",	--5233
		x"04",	--5234
		x"04",	--5235
		x"05",	--5236
		x"05",	--5237
		x"05",	--5238
		x"05",	--5239
		x"05",	--5240
		x"05",	--5241
		x"05",	--5242
		x"05",	--5243
		x"06",	--5244
		x"06",	--5245
		x"06",	--5246
		x"06",	--5247
		x"06",	--5248
		x"06",	--5249
		x"06",	--5250
		x"06",	--5251
		x"06",	--5252
		x"06",	--5253
		x"06",	--5254
		x"06",	--5255
		x"06",	--5256
		x"06",	--5257
		x"06",	--5258
		x"06",	--5259
		x"07",	--5260
		x"07",	--5261
		x"07",	--5262
		x"07",	--5263
		x"07",	--5264
		x"07",	--5265
		x"07",	--5266
		x"07",	--5267
		x"07",	--5268
		x"07",	--5269
		x"07",	--5270
		x"07",	--5271
		x"07",	--5272
		x"07",	--5273
		x"07",	--5274
		x"07",	--5275
		x"07",	--5276
		x"07",	--5277
		x"07",	--5278
		x"07",	--5279
		x"07",	--5280
		x"07",	--5281
		x"07",	--5282
		x"07",	--5283
		x"07",	--5284
		x"07",	--5285
		x"07",	--5286
		x"07",	--5287
		x"07",	--5288
		x"07",	--5289
		x"07",	--5290
		x"07",	--5291
		x"08",	--5292
		x"08",	--5293
		x"08",	--5294
		x"08",	--5295
		x"08",	--5296
		x"08",	--5297
		x"08",	--5298
		x"08",	--5299
		x"08",	--5300
		x"08",	--5301
		x"08",	--5302
		x"08",	--5303
		x"08",	--5304
		x"08",	--5305
		x"08",	--5306
		x"08",	--5307
		x"08",	--5308
		x"08",	--5309
		x"08",	--5310
		x"08",	--5311
		x"08",	--5312
		x"08",	--5313
		x"08",	--5314
		x"08",	--5315
		x"08",	--5316
		x"08",	--5317
		x"08",	--5318
		x"08",	--5319
		x"08",	--5320
		x"08",	--5321
		x"08",	--5322
		x"08",	--5323
		x"08",	--5324
		x"08",	--5325
		x"08",	--5326
		x"08",	--5327
		x"08",	--5328
		x"08",	--5329
		x"08",	--5330
		x"08",	--5331
		x"08",	--5332
		x"08",	--5333
		x"08",	--5334
		x"08",	--5335
		x"08",	--5336
		x"08",	--5337
		x"08",	--5338
		x"08",	--5339
		x"08",	--5340
		x"08",	--5341
		x"08",	--5342
		x"08",	--5343
		x"08",	--5344
		x"08",	--5345
		x"08",	--5346
		x"08",	--5347
		x"08",	--5348
		x"08",	--5349
		x"08",	--5350
		x"08",	--5351
		x"08",	--5352
		x"08",	--5353
		x"08",	--5354
		x"08",	--5355
		x"6e",	--5356
		x"6c",	--5357
		x"29",	--5358
		x"00",	--5359
		x"ff",	--5360
		x"ff",	--5361
		x"65",	--5362
		x"70",	--5363
		x"00",	--5364
		x"ff",	--5365
		x"ff",	--5366
		x"ff",	--5367
		x"ff",	--5368
		x"ff",	--5369
		x"ff",	--5370
		x"ff",	--5371
		x"ff",	--5372
		x"ff",	--5373
		x"ff",	--5374
		x"ff",	--5375
		x"ff",	--5376
		x"ff",	--5377
		x"ff",	--5378
		x"ff",	--5379
		x"ff",	--5380
		x"ff",	--5381
		x"ff",	--5382
		x"ff",	--5383
		x"ff",	--5384
		x"ff",	--5385
		x"ff",	--5386
		x"ff",	--5387
		x"ff",	--5388
		x"ff",	--5389
		x"ff",	--5390
		x"ff",	--5391
		x"ff",	--5392
		x"ff",	--5393
		x"ff",	--5394
		x"ff",	--5395
		x"ff",	--5396
		x"ff",	--5397
		x"ff",	--5398
		x"ff",	--5399
		x"ff",	--5400
		x"ff",	--5401
		x"ff",	--5402
		x"ff",	--5403
		x"ff",	--5404
		x"ff",	--5405
		x"ff",	--5406
		x"ff",	--5407
		x"ff",	--5408
		x"ff",	--5409
		x"ff",	--5410
		x"ff",	--5411
		x"ff",	--5412
		x"ff",	--5413
		x"ff",	--5414
		x"ff",	--5415
		x"ff",	--5416
		x"ff",	--5417
		x"ff",	--5418
		x"ff",	--5419
		x"ff",	--5420
		x"ff",	--5421
		x"ff",	--5422
		x"ff",	--5423
		x"ff",	--5424
		x"ff",	--5425
		x"ff",	--5426
		x"ff",	--5427
		x"ff",	--5428
		x"ff",	--5429
		x"ff",	--5430
		x"ff",	--5431
		x"ff",	--5432
		x"ff",	--5433
		x"ff",	--5434
		x"ff",	--5435
		x"ff",	--5436
		x"ff",	--5437
		x"ff",	--5438
		x"ff",	--5439
		x"ff",	--5440
		x"ff",	--5441
		x"ff",	--5442
		x"ff",	--5443
		x"ff",	--5444
		x"ff",	--5445
		x"ff",	--5446
		x"ff",	--5447
		x"ff",	--5448
		x"ff",	--5449
		x"ff",	--5450
		x"ff",	--5451
		x"ff",	--5452
		x"ff",	--5453
		x"ff",	--5454
		x"ff",	--5455
		x"ff",	--5456
		x"ff",	--5457
		x"ff",	--5458
		x"ff",	--5459
		x"ff",	--5460
		x"ff",	--5461
		x"ff",	--5462
		x"ff",	--5463
		x"ff",	--5464
		x"ff",	--5465
		x"ff",	--5466
		x"ff",	--5467
		x"ff",	--5468
		x"ff",	--5469
		x"ff",	--5470
		x"ff",	--5471
		x"ff",	--5472
		x"ff",	--5473
		x"ff",	--5474
		x"ff",	--5475
		x"ff",	--5476
		x"ff",	--5477
		x"ff",	--5478
		x"ff",	--5479
		x"ff",	--5480
		x"ff",	--5481
		x"ff",	--5482
		x"ff",	--5483
		x"ff",	--5484
		x"ff",	--5485
		x"ff",	--5486
		x"ff",	--5487
		x"ff",	--5488
		x"ff",	--5489
		x"ff",	--5490
		x"ff",	--5491
		x"ff",	--5492
		x"ff",	--5493
		x"ff",	--5494
		x"ff",	--5495
		x"ff",	--5496
		x"ff",	--5497
		x"ff",	--5498
		x"ff",	--5499
		x"ff",	--5500
		x"ff",	--5501
		x"ff",	--5502
		x"ff",	--5503
		x"ff",	--5504
		x"ff",	--5505
		x"ff",	--5506
		x"ff",	--5507
		x"ff",	--5508
		x"ff",	--5509
		x"ff",	--5510
		x"ff",	--5511
		x"ff",	--5512
		x"ff",	--5513
		x"ff",	--5514
		x"ff",	--5515
		x"ff",	--5516
		x"ff",	--5517
		x"ff",	--5518
		x"ff",	--5519
		x"ff",	--5520
		x"ff",	--5521
		x"ff",	--5522
		x"ff",	--5523
		x"ff",	--5524
		x"ff",	--5525
		x"ff",	--5526
		x"ff",	--5527
		x"ff",	--5528
		x"ff",	--5529
		x"ff",	--5530
		x"ff",	--5531
		x"ff",	--5532
		x"ff",	--5533
		x"ff",	--5534
		x"ff",	--5535
		x"ff",	--5536
		x"ff",	--5537
		x"ff",	--5538
		x"ff",	--5539
		x"ff",	--5540
		x"ff",	--5541
		x"ff",	--5542
		x"ff",	--5543
		x"ff",	--5544
		x"ff",	--5545
		x"ff",	--5546
		x"ff",	--5547
		x"ff",	--5548
		x"ff",	--5549
		x"ff",	--5550
		x"ff",	--5551
		x"ff",	--5552
		x"ff",	--5553
		x"ff",	--5554
		x"ff",	--5555
		x"ff",	--5556
		x"ff",	--5557
		x"ff",	--5558
		x"ff",	--5559
		x"ff",	--5560
		x"ff",	--5561
		x"ff",	--5562
		x"ff",	--5563
		x"ff",	--5564
		x"ff",	--5565
		x"ff",	--5566
		x"ff",	--5567
		x"ff",	--5568
		x"ff",	--5569
		x"ff",	--5570
		x"ff",	--5571
		x"ff",	--5572
		x"ff",	--5573
		x"ff",	--5574
		x"ff",	--5575
		x"ff",	--5576
		x"ff",	--5577
		x"ff",	--5578
		x"ff",	--5579
		x"ff",	--5580
		x"ff",	--5581
		x"ff",	--5582
		x"ff",	--5583
		x"ff",	--5584
		x"ff",	--5585
		x"ff",	--5586
		x"ff",	--5587
		x"ff",	--5588
		x"ff",	--5589
		x"ff",	--5590
		x"ff",	--5591
		x"ff",	--5592
		x"ff",	--5593
		x"ff",	--5594
		x"ff",	--5595
		x"ff",	--5596
		x"ff",	--5597
		x"ff",	--5598
		x"ff",	--5599
		x"ff",	--5600
		x"ff",	--5601
		x"ff",	--5602
		x"ff",	--5603
		x"ff",	--5604
		x"ff",	--5605
		x"ff",	--5606
		x"ff",	--5607
		x"ff",	--5608
		x"ff",	--5609
		x"ff",	--5610
		x"ff",	--5611
		x"ff",	--5612
		x"ff",	--5613
		x"ff",	--5614
		x"ff",	--5615
		x"ff",	--5616
		x"ff",	--5617
		x"ff",	--5618
		x"ff",	--5619
		x"ff",	--5620
		x"ff",	--5621
		x"ff",	--5622
		x"ff",	--5623
		x"ff",	--5624
		x"ff",	--5625
		x"ff",	--5626
		x"ff",	--5627
		x"ff",	--5628
		x"ff",	--5629
		x"ff",	--5630
		x"ff",	--5631
		x"ff",	--5632
		x"ff",	--5633
		x"ff",	--5634
		x"ff",	--5635
		x"ff",	--5636
		x"ff",	--5637
		x"ff",	--5638
		x"ff",	--5639
		x"ff",	--5640
		x"ff",	--5641
		x"ff",	--5642
		x"ff",	--5643
		x"ff",	--5644
		x"ff",	--5645
		x"ff",	--5646
		x"ff",	--5647
		x"ff",	--5648
		x"ff",	--5649
		x"ff",	--5650
		x"ff",	--5651
		x"ff",	--5652
		x"ff",	--5653
		x"ff",	--5654
		x"ff",	--5655
		x"ff",	--5656
		x"ff",	--5657
		x"ff",	--5658
		x"ff",	--5659
		x"ff",	--5660
		x"ff",	--5661
		x"ff",	--5662
		x"ff",	--5663
		x"ff",	--5664
		x"ff",	--5665
		x"ff",	--5666
		x"ff",	--5667
		x"ff",	--5668
		x"ff",	--5669
		x"ff",	--5670
		x"ff",	--5671
		x"ff",	--5672
		x"ff",	--5673
		x"ff",	--5674
		x"ff",	--5675
		x"ff",	--5676
		x"ff",	--5677
		x"ff",	--5678
		x"ff",	--5679
		x"ff",	--5680
		x"ff",	--5681
		x"ff",	--5682
		x"ff",	--5683
		x"ff",	--5684
		x"ff",	--5685
		x"ff",	--5686
		x"ff",	--5687
		x"ff",	--5688
		x"ff",	--5689
		x"ff",	--5690
		x"ff",	--5691
		x"ff",	--5692
		x"ff",	--5693
		x"ff",	--5694
		x"ff",	--5695
		x"ff",	--5696
		x"ff",	--5697
		x"ff",	--5698
		x"ff",	--5699
		x"ff",	--5700
		x"ff",	--5701
		x"ff",	--5702
		x"ff",	--5703
		x"ff",	--5704
		x"ff",	--5705
		x"ff",	--5706
		x"ff",	--5707
		x"ff",	--5708
		x"ff",	--5709
		x"ff",	--5710
		x"ff",	--5711
		x"ff",	--5712
		x"ff",	--5713
		x"ff",	--5714
		x"ff",	--5715
		x"ff",	--5716
		x"ff",	--5717
		x"ff",	--5718
		x"ff",	--5719
		x"ff",	--5720
		x"ff",	--5721
		x"ff",	--5722
		x"ff",	--5723
		x"ff",	--5724
		x"ff",	--5725
		x"ff",	--5726
		x"ff",	--5727
		x"ff",	--5728
		x"ff",	--5729
		x"ff",	--5730
		x"ff",	--5731
		x"ff",	--5732
		x"ff",	--5733
		x"ff",	--5734
		x"ff",	--5735
		x"ff",	--5736
		x"ff",	--5737
		x"ff",	--5738
		x"ff",	--5739
		x"ff",	--5740
		x"ff",	--5741
		x"ff",	--5742
		x"ff",	--5743
		x"ff",	--5744
		x"ff",	--5745
		x"ff",	--5746
		x"ff",	--5747
		x"ff",	--5748
		x"ff",	--5749
		x"ff",	--5750
		x"ff",	--5751
		x"ff",	--5752
		x"ff",	--5753
		x"ff",	--5754
		x"ff",	--5755
		x"ff",	--5756
		x"ff",	--5757
		x"ff",	--5758
		x"ff",	--5759
		x"ff",	--5760
		x"ff",	--5761
		x"ff",	--5762
		x"ff",	--5763
		x"ff",	--5764
		x"ff",	--5765
		x"ff",	--5766
		x"ff",	--5767
		x"ff",	--5768
		x"ff",	--5769
		x"ff",	--5770
		x"ff",	--5771
		x"ff",	--5772
		x"ff",	--5773
		x"ff",	--5774
		x"ff",	--5775
		x"ff",	--5776
		x"ff",	--5777
		x"ff",	--5778
		x"ff",	--5779
		x"ff",	--5780
		x"ff",	--5781
		x"ff",	--5782
		x"ff",	--5783
		x"ff",	--5784
		x"ff",	--5785
		x"ff",	--5786
		x"ff",	--5787
		x"ff",	--5788
		x"ff",	--5789
		x"ff",	--5790
		x"ff",	--5791
		x"ff",	--5792
		x"ff",	--5793
		x"ff",	--5794
		x"ff",	--5795
		x"ff",	--5796
		x"ff",	--5797
		x"ff",	--5798
		x"ff",	--5799
		x"ff",	--5800
		x"ff",	--5801
		x"ff",	--5802
		x"ff",	--5803
		x"ff",	--5804
		x"ff",	--5805
		x"ff",	--5806
		x"ff",	--5807
		x"ff",	--5808
		x"ff",	--5809
		x"ff",	--5810
		x"ff",	--5811
		x"ff",	--5812
		x"ff",	--5813
		x"ff",	--5814
		x"ff",	--5815
		x"ff",	--5816
		x"ff",	--5817
		x"ff",	--5818
		x"ff",	--5819
		x"ff",	--5820
		x"ff",	--5821
		x"ff",	--5822
		x"ff",	--5823
		x"ff",	--5824
		x"ff",	--5825
		x"ff",	--5826
		x"ff",	--5827
		x"ff",	--5828
		x"ff",	--5829
		x"ff",	--5830
		x"ff",	--5831
		x"ff",	--5832
		x"ff",	--5833
		x"ff",	--5834
		x"ff",	--5835
		x"ff",	--5836
		x"ff",	--5837
		x"ff",	--5838
		x"ff",	--5839
		x"ff",	--5840
		x"ff",	--5841
		x"ff",	--5842
		x"ff",	--5843
		x"ff",	--5844
		x"ff",	--5845
		x"ff",	--5846
		x"ff",	--5847
		x"ff",	--5848
		x"ff",	--5849
		x"ff",	--5850
		x"ff",	--5851
		x"ff",	--5852
		x"ff",	--5853
		x"ff",	--5854
		x"ff",	--5855
		x"ff",	--5856
		x"ff",	--5857
		x"ff",	--5858
		x"ff",	--5859
		x"ff",	--5860
		x"ff",	--5861
		x"ff",	--5862
		x"ff",	--5863
		x"ff",	--5864
		x"ff",	--5865
		x"ff",	--5866
		x"ff",	--5867
		x"ff",	--5868
		x"ff",	--5869
		x"ff",	--5870
		x"ff",	--5871
		x"ff",	--5872
		x"ff",	--5873
		x"ff",	--5874
		x"ff",	--5875
		x"ff",	--5876
		x"ff",	--5877
		x"ff",	--5878
		x"ff",	--5879
		x"ff",	--5880
		x"ff",	--5881
		x"ff",	--5882
		x"ff",	--5883
		x"ff",	--5884
		x"ff",	--5885
		x"ff",	--5886
		x"ff",	--5887
		x"ff",	--5888
		x"ff",	--5889
		x"ff",	--5890
		x"ff",	--5891
		x"ff",	--5892
		x"ff",	--5893
		x"ff",	--5894
		x"ff",	--5895
		x"ff",	--5896
		x"ff",	--5897
		x"ff",	--5898
		x"ff",	--5899
		x"ff",	--5900
		x"ff",	--5901
		x"ff",	--5902
		x"ff",	--5903
		x"ff",	--5904
		x"ff",	--5905
		x"ff",	--5906
		x"ff",	--5907
		x"ff",	--5908
		x"ff",	--5909
		x"ff",	--5910
		x"ff",	--5911
		x"ff",	--5912
		x"ff",	--5913
		x"ff",	--5914
		x"ff",	--5915
		x"ff",	--5916
		x"ff",	--5917
		x"ff",	--5918
		x"ff",	--5919
		x"ff",	--5920
		x"ff",	--5921
		x"ff",	--5922
		x"ff",	--5923
		x"ff",	--5924
		x"ff",	--5925
		x"ff",	--5926
		x"ff",	--5927
		x"ff",	--5928
		x"ff",	--5929
		x"ff",	--5930
		x"ff",	--5931
		x"ff",	--5932
		x"ff",	--5933
		x"ff",	--5934
		x"ff",	--5935
		x"ff",	--5936
		x"ff",	--5937
		x"ff",	--5938
		x"ff",	--5939
		x"ff",	--5940
		x"ff",	--5941
		x"ff",	--5942
		x"ff",	--5943
		x"ff",	--5944
		x"ff",	--5945
		x"ff",	--5946
		x"ff",	--5947
		x"ff",	--5948
		x"ff",	--5949
		x"ff",	--5950
		x"ff",	--5951
		x"ff",	--5952
		x"ff",	--5953
		x"ff",	--5954
		x"ff",	--5955
		x"ff",	--5956
		x"ff",	--5957
		x"ff",	--5958
		x"ff",	--5959
		x"ff",	--5960
		x"ff",	--5961
		x"ff",	--5962
		x"ff",	--5963
		x"ff",	--5964
		x"ff",	--5965
		x"ff",	--5966
		x"ff",	--5967
		x"ff",	--5968
		x"ff",	--5969
		x"ff",	--5970
		x"ff",	--5971
		x"ff",	--5972
		x"ff",	--5973
		x"ff",	--5974
		x"ff",	--5975
		x"ff",	--5976
		x"ff",	--5977
		x"ff",	--5978
		x"ff",	--5979
		x"ff",	--5980
		x"ff",	--5981
		x"ff",	--5982
		x"ff",	--5983
		x"ff",	--5984
		x"ff",	--5985
		x"ff",	--5986
		x"ff",	--5987
		x"ff",	--5988
		x"ff",	--5989
		x"ff",	--5990
		x"ff",	--5991
		x"ff",	--5992
		x"ff",	--5993
		x"ff",	--5994
		x"ff",	--5995
		x"ff",	--5996
		x"ff",	--5997
		x"ff",	--5998
		x"ff",	--5999
		x"ff",	--6000
		x"ff",	--6001
		x"ff",	--6002
		x"ff",	--6003
		x"ff",	--6004
		x"ff",	--6005
		x"ff",	--6006
		x"ff",	--6007
		x"ff",	--6008
		x"ff",	--6009
		x"ff",	--6010
		x"ff",	--6011
		x"ff",	--6012
		x"ff",	--6013
		x"ff",	--6014
		x"ff",	--6015
		x"ff",	--6016
		x"ff",	--6017
		x"ff",	--6018
		x"ff",	--6019
		x"ff",	--6020
		x"ff",	--6021
		x"ff",	--6022
		x"ff",	--6023
		x"ff",	--6024
		x"ff",	--6025
		x"ff",	--6026
		x"ff",	--6027
		x"ff",	--6028
		x"ff",	--6029
		x"ff",	--6030
		x"ff",	--6031
		x"ff",	--6032
		x"ff",	--6033
		x"ff",	--6034
		x"ff",	--6035
		x"ff",	--6036
		x"ff",	--6037
		x"ff",	--6038
		x"ff",	--6039
		x"ff",	--6040
		x"ff",	--6041
		x"ff",	--6042
		x"ff",	--6043
		x"ff",	--6044
		x"ff",	--6045
		x"ff",	--6046
		x"ff",	--6047
		x"ff",	--6048
		x"ff",	--6049
		x"ff",	--6050
		x"ff",	--6051
		x"ff",	--6052
		x"ff",	--6053
		x"ff",	--6054
		x"ff",	--6055
		x"ff",	--6056
		x"ff",	--6057
		x"ff",	--6058
		x"ff",	--6059
		x"ff",	--6060
		x"ff",	--6061
		x"ff",	--6062
		x"ff",	--6063
		x"ff",	--6064
		x"ff",	--6065
		x"ff",	--6066
		x"ff",	--6067
		x"ff",	--6068
		x"ff",	--6069
		x"ff",	--6070
		x"ff",	--6071
		x"ff",	--6072
		x"ff",	--6073
		x"ff",	--6074
		x"ff",	--6075
		x"ff",	--6076
		x"ff",	--6077
		x"ff",	--6078
		x"ff",	--6079
		x"ff",	--6080
		x"ff",	--6081
		x"ff",	--6082
		x"ff",	--6083
		x"ff",	--6084
		x"ff",	--6085
		x"ff",	--6086
		x"ff",	--6087
		x"ff",	--6088
		x"ff",	--6089
		x"ff",	--6090
		x"ff",	--6091
		x"ff",	--6092
		x"ff",	--6093
		x"ff",	--6094
		x"ff",	--6095
		x"ff",	--6096
		x"ff",	--6097
		x"ff",	--6098
		x"ff",	--6099
		x"ff",	--6100
		x"ff",	--6101
		x"ff",	--6102
		x"ff",	--6103
		x"ff",	--6104
		x"ff",	--6105
		x"ff",	--6106
		x"ff",	--6107
		x"ff",	--6108
		x"ff",	--6109
		x"ff",	--6110
		x"ff",	--6111
		x"ff",	--6112
		x"ff",	--6113
		x"ff",	--6114
		x"ff",	--6115
		x"ff",	--6116
		x"ff",	--6117
		x"ff",	--6118
		x"ff",	--6119
		x"ff",	--6120
		x"ff",	--6121
		x"ff",	--6122
		x"ff",	--6123
		x"ff",	--6124
		x"ff",	--6125
		x"ff",	--6126
		x"ff",	--6127
		x"ff",	--6128
		x"ff",	--6129
		x"ff",	--6130
		x"ff",	--6131
		x"ff",	--6132
		x"ff",	--6133
		x"ff",	--6134
		x"ff",	--6135
		x"ff",	--6136
		x"ff",	--6137
		x"ff",	--6138
		x"ff",	--6139
		x"ff",	--6140
		x"ff",	--6141
		x"ff",	--6142
		x"ff",	--6143
		x"ff",	--6144
		x"ff",	--6145
		x"ff",	--6146
		x"ff",	--6147
		x"ff",	--6148
		x"ff",	--6149
		x"ff",	--6150
		x"ff",	--6151
		x"ff",	--6152
		x"ff",	--6153
		x"ff",	--6154
		x"ff",	--6155
		x"ff",	--6156
		x"ff",	--6157
		x"ff",	--6158
		x"ff",	--6159
		x"ff",	--6160
		x"ff",	--6161
		x"ff",	--6162
		x"ff",	--6163
		x"ff",	--6164
		x"ff",	--6165
		x"ff",	--6166
		x"ff",	--6167
		x"ff",	--6168
		x"ff",	--6169
		x"ff",	--6170
		x"ff",	--6171
		x"ff",	--6172
		x"ff",	--6173
		x"ff",	--6174
		x"ff",	--6175
		x"ff",	--6176
		x"ff",	--6177
		x"ff",	--6178
		x"ff",	--6179
		x"ff",	--6180
		x"ff",	--6181
		x"ff",	--6182
		x"ff",	--6183
		x"ff",	--6184
		x"ff",	--6185
		x"ff",	--6186
		x"ff",	--6187
		x"ff",	--6188
		x"ff",	--6189
		x"ff",	--6190
		x"ff",	--6191
		x"ff",	--6192
		x"ff",	--6193
		x"ff",	--6194
		x"ff",	--6195
		x"ff",	--6196
		x"ff",	--6197
		x"ff",	--6198
		x"ff",	--6199
		x"ff",	--6200
		x"ff",	--6201
		x"ff",	--6202
		x"ff",	--6203
		x"ff",	--6204
		x"ff",	--6205
		x"ff",	--6206
		x"ff",	--6207
		x"ff",	--6208
		x"ff",	--6209
		x"ff",	--6210
		x"ff",	--6211
		x"ff",	--6212
		x"ff",	--6213
		x"ff",	--6214
		x"ff",	--6215
		x"ff",	--6216
		x"ff",	--6217
		x"ff",	--6218
		x"ff",	--6219
		x"ff",	--6220
		x"ff",	--6221
		x"ff",	--6222
		x"ff",	--6223
		x"ff",	--6224
		x"ff",	--6225
		x"ff",	--6226
		x"ff",	--6227
		x"ff",	--6228
		x"ff",	--6229
		x"ff",	--6230
		x"ff",	--6231
		x"ff",	--6232
		x"ff",	--6233
		x"ff",	--6234
		x"ff",	--6235
		x"ff",	--6236
		x"ff",	--6237
		x"ff",	--6238
		x"ff",	--6239
		x"ff",	--6240
		x"ff",	--6241
		x"ff",	--6242
		x"ff",	--6243
		x"ff",	--6244
		x"ff",	--6245
		x"ff",	--6246
		x"ff",	--6247
		x"ff",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"ff",	--6252
		x"ff",	--6253
		x"ff",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"c2",	--8176
		x"c2",	--8177
		x"c2",	--8178
		x"c2",	--8179
		x"c2",	--8180
		x"c2",	--8181
		x"c2",	--8182
		x"cd",	--8183
		x"ca",	--8184
		x"c2",	--8185
		x"c2",	--8186
		x"c2",	--8187
		x"c2",	--8188
		x"c2",	--8189
		x"c2",	--8190
		x"c0");	--8191

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
