library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"28",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"0c",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"28",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"94",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"1c",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"28",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"0c",	--29
		x"f9",	--30
		x"31",	--31
		x"a4",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"f0",	--44
		x"b0",	--45
		x"72",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"a6",	--50
		x"b0",	--51
		x"b4",	--52
		x"21",	--53
		x"3d",	--54
		x"c3",	--55
		x"3e",	--56
		x"82",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"a2",	--61
		x"3d",	--62
		x"d4",	--63
		x"3e",	--64
		x"a2",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"a2",	--69
		x"3d",	--70
		x"da",	--71
		x"3e",	--72
		x"16",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"a2",	--77
		x"3d",	--78
		x"df",	--79
		x"3e",	--80
		x"6a",	--81
		x"7f",	--82
		x"61",	--83
		x"b0",	--84
		x"a2",	--85
		x"3d",	--86
		x"e6",	--87
		x"3e",	--88
		x"38",	--89
		x"7f",	--90
		x"70",	--91
		x"b0",	--92
		x"a2",	--93
		x"3d",	--94
		x"ea",	--95
		x"3e",	--96
		x"78",	--97
		x"7f",	--98
		x"65",	--99
		x"b0",	--100
		x"a2",	--101
		x"3d",	--102
		x"f2",	--103
		x"3e",	--104
		x"c0",	--105
		x"7f",	--106
		x"73",	--107
		x"b0",	--108
		x"a2",	--109
		x"3d",	--110
		x"03",	--111
		x"3e",	--112
		x"c4",	--113
		x"7f",	--114
		x"63",	--115
		x"b0",	--116
		x"a2",	--117
		x"3d",	--118
		x"17",	--119
		x"3e",	--120
		x"c8",	--121
		x"7f",	--122
		x"62",	--123
		x"b0",	--124
		x"a2",	--125
		x"0e",	--126
		x"0f",	--127
		x"b0",	--128
		x"38",	--129
		x"2c",	--130
		x"3d",	--131
		x"20",	--132
		x"3e",	--133
		x"80",	--134
		x"0f",	--135
		x"3f",	--136
		x"10",	--137
		x"b0",	--138
		x"40",	--139
		x"0f",	--140
		x"3f",	--141
		x"10",	--142
		x"b0",	--143
		x"88",	--144
		x"2c",	--145
		x"3d",	--146
		x"20",	--147
		x"3e",	--148
		x"88",	--149
		x"0f",	--150
		x"3f",	--151
		x"06",	--152
		x"b0",	--153
		x"40",	--154
		x"0f",	--155
		x"3f",	--156
		x"06",	--157
		x"b0",	--158
		x"88",	--159
		x"0e",	--160
		x"3e",	--161
		x"06",	--162
		x"0f",	--163
		x"3f",	--164
		x"10",	--165
		x"b0",	--166
		x"2e",	--167
		x"3e",	--168
		x"98",	--169
		x"0f",	--170
		x"2f",	--171
		x"b0",	--172
		x"96",	--173
		x"3e",	--174
		x"9c",	--175
		x"0f",	--176
		x"2f",	--177
		x"b0",	--178
		x"96",	--179
		x"0e",	--180
		x"2e",	--181
		x"0f",	--182
		x"2f",	--183
		x"b0",	--184
		x"64",	--185
		x"0e",	--186
		x"3e",	--187
		x"06",	--188
		x"0f",	--189
		x"3f",	--190
		x"10",	--191
		x"b0",	--192
		x"6e",	--193
		x"b0",	--194
		x"6e",	--195
		x"3e",	--196
		x"a0",	--197
		x"0f",	--198
		x"b0",	--199
		x"ae",	--200
		x"0f",	--201
		x"b0",	--202
		x"64",	--203
		x"3d",	--204
		x"64",	--205
		x"3e",	--206
		x"70",	--207
		x"0f",	--208
		x"b0",	--209
		x"c2",	--210
		x"0c",	--211
		x"0d",	--212
		x"1e",	--213
		x"0f",	--214
		x"3f",	--215
		x"26",	--216
		x"b0",	--217
		x"f6",	--218
		x"0c",	--219
		x"0d",	--220
		x"1e",	--221
		x"0f",	--222
		x"3f",	--223
		x"1a",	--224
		x"b0",	--225
		x"f6",	--226
		x"0e",	--227
		x"3e",	--228
		x"1a",	--229
		x"0f",	--230
		x"3f",	--231
		x"26",	--232
		x"b0",	--233
		x"be",	--234
		x"f2",	--235
		x"80",	--236
		x"19",	--237
		x"32",	--238
		x"0b",	--239
		x"b0",	--240
		x"0e",	--241
		x"0f",	--242
		x"fc",	--243
		x"b0",	--244
		x"36",	--245
		x"7f",	--246
		x"15",	--247
		x"7f",	--248
		x"0d",	--249
		x"1b",	--250
		x"30",	--251
		x"22",	--252
		x"b0",	--253
		x"b4",	--254
		x"21",	--255
		x"3f",	--256
		x"32",	--257
		x"0f",	--258
		x"0b",	--259
		x"cb",	--260
		x"00",	--261
		x"0e",	--262
		x"5f",	--263
		x"32",	--264
		x"b0",	--265
		x"d6",	--266
		x"0b",	--267
		x"e3",	--268
		x"0b",	--269
		x"e1",	--270
		x"3b",	--271
		x"30",	--272
		x"25",	--273
		x"b0",	--274
		x"b4",	--275
		x"21",	--276
		x"da",	--277
		x"3b",	--278
		x"28",	--279
		x"d7",	--280
		x"82",	--281
		x"0e",	--282
		x"0c",	--283
		x"4e",	--284
		x"8e",	--285
		x"0e",	--286
		x"30",	--287
		x"29",	--288
		x"81",	--289
		x"5e",	--290
		x"b0",	--291
		x"b4",	--292
		x"21",	--293
		x"1f",	--294
		x"5a",	--295
		x"3e",	--296
		x"32",	--297
		x"0e",	--298
		x"0e",	--299
		x"ce",	--300
		x"00",	--301
		x"1b",	--302
		x"c0",	--303
		x"30",	--304
		x"ec",	--305
		x"82",	--306
		x"1e",	--307
		x"30",	--308
		x"0b",	--309
		x"0a",	--310
		x"21",	--311
		x"0a",	--312
		x"0b",	--313
		x"2f",	--314
		x"1b",	--315
		x"0e",	--316
		x"1f",	--317
		x"02",	--318
		x"b0",	--319
		x"72",	--320
		x"0d",	--321
		x"2a",	--322
		x"18",	--323
		x"0e",	--324
		x"1f",	--325
		x"04",	--326
		x"81",	--327
		x"02",	--328
		x"b0",	--329
		x"72",	--330
		x"0e",	--331
		x"1d",	--332
		x"02",	--333
		x"1f",	--334
		x"1e",	--335
		x"b0",	--336
		x"c2",	--337
		x"0f",	--338
		x"21",	--339
		x"3a",	--340
		x"3b",	--341
		x"30",	--342
		x"3d",	--343
		x"64",	--344
		x"3e",	--345
		x"70",	--346
		x"f2",	--347
		x"3e",	--348
		x"70",	--349
		x"ef",	--350
		x"30",	--351
		x"0f",	--352
		x"30",	--353
		x"0f",	--354
		x"30",	--355
		x"b2",	--356
		x"00",	--357
		x"92",	--358
		x"b2",	--359
		x"30",	--360
		x"94",	--361
		x"b2",	--362
		x"41",	--363
		x"96",	--364
		x"30",	--365
		x"f4",	--366
		x"b0",	--367
		x"b4",	--368
		x"92",	--369
		x"90",	--370
		x"b1",	--371
		x"12",	--372
		x"00",	--373
		x"b0",	--374
		x"b4",	--375
		x"21",	--376
		x"0f",	--377
		x"30",	--378
		x"b0",	--379
		x"08",	--380
		x"30",	--381
		x"0b",	--382
		x"0a",	--383
		x"0a",	--384
		x"3b",	--385
		x"00",	--386
		x"0d",	--387
		x"0e",	--388
		x"1f",	--389
		x"22",	--390
		x"b0",	--391
		x"dc",	--392
		x"0d",	--393
		x"0e",	--394
		x"1f",	--395
		x"20",	--396
		x"b0",	--397
		x"dc",	--398
		x"30",	--399
		x"2b",	--400
		x"b0",	--401
		x"b4",	--402
		x"21",	--403
		x"3a",	--404
		x"3b",	--405
		x"30",	--406
		x"82",	--407
		x"22",	--408
		x"82",	--409
		x"20",	--410
		x"30",	--411
		x"0b",	--412
		x"0a",	--413
		x"21",	--414
		x"0a",	--415
		x"0b",	--416
		x"b2",	--417
		x"00",	--418
		x"4e",	--419
		x"3a",	--420
		x"03",	--421
		x"53",	--422
		x"3e",	--423
		x"0e",	--424
		x"1f",	--425
		x"02",	--426
		x"b0",	--427
		x"72",	--428
		x"0a",	--429
		x"0e",	--430
		x"1f",	--431
		x"04",	--432
		x"b0",	--433
		x"72",	--434
		x"0b",	--435
		x"0f",	--436
		x"0a",	--437
		x"30",	--438
		x"78",	--439
		x"b0",	--440
		x"b4",	--441
		x"31",	--442
		x"06",	--443
		x"0e",	--444
		x"0f",	--445
		x"b0",	--446
		x"28",	--447
		x"0c",	--448
		x"3d",	--449
		x"c8",	--450
		x"b0",	--451
		x"f8",	--452
		x"0c",	--453
		x"0d",	--454
		x"0e",	--455
		x"3f",	--456
		x"80",	--457
		x"b0",	--458
		x"84",	--459
		x"0d",	--460
		x"0e",	--461
		x"1f",	--462
		x"22",	--463
		x"b0",	--464
		x"dc",	--465
		x"0e",	--466
		x"0f",	--467
		x"b0",	--468
		x"28",	--469
		x"0c",	--470
		x"3d",	--471
		x"c8",	--472
		x"b0",	--473
		x"f8",	--474
		x"0d",	--475
		x"0e",	--476
		x"1f",	--477
		x"20",	--478
		x"b0",	--479
		x"dc",	--480
		x"0f",	--481
		x"21",	--482
		x"3a",	--483
		x"3b",	--484
		x"30",	--485
		x"0e",	--486
		x"1f",	--487
		x"06",	--488
		x"b0",	--489
		x"72",	--490
		x"1d",	--491
		x"0e",	--492
		x"1f",	--493
		x"00",	--494
		x"b0",	--495
		x"c2",	--496
		x"b6",	--497
		x"0e",	--498
		x"3f",	--499
		x"fc",	--500
		x"b0",	--501
		x"7e",	--502
		x"82",	--503
		x"00",	--504
		x"aa",	--505
		x"30",	--506
		x"32",	--507
		x"b0",	--508
		x"b4",	--509
		x"b1",	--510
		x"4c",	--511
		x"00",	--512
		x"b0",	--513
		x"b4",	--514
		x"a1",	--515
		x"00",	--516
		x"30",	--517
		x"5d",	--518
		x"b0",	--519
		x"b4",	--520
		x"21",	--521
		x"3f",	--522
		x"d6",	--523
		x"0b",	--524
		x"0a",	--525
		x"1f",	--526
		x"26",	--527
		x"b0",	--528
		x"9e",	--529
		x"0a",	--530
		x"0b",	--531
		x"1f",	--532
		x"24",	--533
		x"b0",	--534
		x"9e",	--535
		x"0b",	--536
		x"0a",	--537
		x"3e",	--538
		x"3f",	--539
		x"1e",	--540
		x"0f",	--541
		x"0f",	--542
		x"0e",	--543
		x"30",	--544
		x"80",	--545
		x"30",	--546
		x"28",	--547
		x"b0",	--548
		x"80",	--549
		x"31",	--550
		x"0c",	--551
		x"30",	--552
		x"28",	--553
		x"30",	--554
		x"88",	--555
		x"b0",	--556
		x"b4",	--557
		x"21",	--558
		x"3a",	--559
		x"3b",	--560
		x"30",	--561
		x"82",	--562
		x"24",	--563
		x"82",	--564
		x"26",	--565
		x"30",	--566
		x"82",	--567
		x"22",	--568
		x"82",	--569
		x"20",	--570
		x"30",	--571
		x"0b",	--572
		x"0a",	--573
		x"09",	--574
		x"08",	--575
		x"21",	--576
		x"0a",	--577
		x"0b",	--578
		x"81",	--579
		x"00",	--580
		x"1f",	--581
		x"1c",	--582
		x"b2",	--583
		x"02",	--584
		x"6f",	--585
		x"92",	--586
		x"0c",	--587
		x"0e",	--588
		x"1f",	--589
		x"02",	--590
		x"b0",	--591
		x"72",	--592
		x"08",	--593
		x"3a",	--594
		x"03",	--595
		x"1e",	--596
		x"09",	--597
		x"0d",	--598
		x"0e",	--599
		x"1f",	--600
		x"02",	--601
		x"b0",	--602
		x"c2",	--603
		x"0f",	--604
		x"21",	--605
		x"38",	--606
		x"39",	--607
		x"3a",	--608
		x"3b",	--609
		x"30",	--610
		x"82",	--611
		x"0c",	--612
		x"49",	--613
		x"82",	--614
		x"0c",	--615
		x"1f",	--616
		x"02",	--617
		x"b0",	--618
		x"ea",	--619
		x"0f",	--620
		x"21",	--621
		x"38",	--622
		x"39",	--623
		x"3a",	--624
		x"3b",	--625
		x"30",	--626
		x"0e",	--627
		x"1f",	--628
		x"04",	--629
		x"b0",	--630
		x"72",	--631
		x"09",	--632
		x"3a",	--633
		x"05",	--634
		x"da",	--635
		x"0e",	--636
		x"1f",	--637
		x"06",	--638
		x"b0",	--639
		x"72",	--640
		x"0a",	--641
		x"0e",	--642
		x"1f",	--643
		x"08",	--644
		x"b0",	--645
		x"72",	--646
		x"0b",	--647
		x"0f",	--648
		x"0a",	--649
		x"30",	--650
		x"8d",	--651
		x"b0",	--652
		x"b4",	--653
		x"31",	--654
		x"06",	--655
		x"0e",	--656
		x"0f",	--657
		x"b0",	--658
		x"28",	--659
		x"0c",	--660
		x"3d",	--661
		x"c8",	--662
		x"b0",	--663
		x"f8",	--664
		x"0d",	--665
		x"0e",	--666
		x"1f",	--667
		x"22",	--668
		x"b0",	--669
		x"dc",	--670
		x"0e",	--671
		x"0f",	--672
		x"b0",	--673
		x"28",	--674
		x"0c",	--675
		x"3d",	--676
		x"c8",	--677
		x"b0",	--678
		x"f8",	--679
		x"0d",	--680
		x"0e",	--681
		x"1f",	--682
		x"20",	--683
		x"b0",	--684
		x"dc",	--685
		x"a7",	--686
		x"0f",	--687
		x"b0",	--688
		x"18",	--689
		x"0f",	--690
		x"21",	--691
		x"38",	--692
		x"39",	--693
		x"3a",	--694
		x"3b",	--695
		x"30",	--696
		x"0e",	--697
		x"3f",	--698
		x"18",	--699
		x"b0",	--700
		x"7e",	--701
		x"82",	--702
		x"02",	--703
		x"89",	--704
		x"1f",	--705
		x"82",	--706
		x"0e",	--707
		x"01",	--708
		x"0f",	--709
		x"82",	--710
		x"0e",	--711
		x"0f",	--712
		x"30",	--713
		x"5e",	--714
		x"19",	--715
		x"4e",	--716
		x"0f",	--717
		x"03",	--718
		x"c2",	--719
		x"19",	--720
		x"30",	--721
		x"c2",	--722
		x"19",	--723
		x"30",	--724
		x"1e",	--725
		x"10",	--726
		x"3e",	--727
		x"06",	--728
		x"0f",	--729
		x"0f",	--730
		x"10",	--731
		x"96",	--732
		x"c2",	--733
		x"19",	--734
		x"3e",	--735
		x"07",	--736
		x"03",	--737
		x"82",	--738
		x"10",	--739
		x"30",	--740
		x"1e",	--741
		x"82",	--742
		x"10",	--743
		x"30",	--744
		x"f2",	--745
		x"0e",	--746
		x"19",	--747
		x"f2",	--748
		x"f2",	--749
		x"0a",	--750
		x"19",	--751
		x"ee",	--752
		x"e2",	--753
		x"19",	--754
		x"eb",	--755
		x"f2",	--756
		x"0d",	--757
		x"19",	--758
		x"e7",	--759
		x"f2",	--760
		x"09",	--761
		x"19",	--762
		x"e3",	--763
		x"f2",	--764
		x"03",	--765
		x"19",	--766
		x"df",	--767
		x"f2",	--768
		x"07",	--769
		x"19",	--770
		x"db",	--771
		x"8f",	--772
		x"00",	--773
		x"8f",	--774
		x"02",	--775
		x"8f",	--776
		x"04",	--777
		x"8f",	--778
		x"06",	--779
		x"8f",	--780
		x"08",	--781
		x"8f",	--782
		x"0a",	--783
		x"30",	--784
		x"8f",	--785
		x"06",	--786
		x"8f",	--787
		x"08",	--788
		x"8f",	--789
		x"0a",	--790
		x"30",	--791
		x"8f",	--792
		x"00",	--793
		x"30",	--794
		x"8f",	--795
		x"02",	--796
		x"30",	--797
		x"8f",	--798
		x"04",	--799
		x"30",	--800
		x"8f",	--801
		x"06",	--802
		x"30",	--803
		x"1d",	--804
		x"06",	--805
		x"0d",	--806
		x"0e",	--807
		x"1d",	--808
		x"08",	--809
		x"8f",	--810
		x"08",	--811
		x"02",	--812
		x"32",	--813
		x"03",	--814
		x"82",	--815
		x"32",	--816
		x"a2",	--817
		x"38",	--818
		x"1c",	--819
		x"3a",	--820
		x"32",	--821
		x"02",	--822
		x"32",	--823
		x"03",	--824
		x"82",	--825
		x"32",	--826
		x"92",	--827
		x"02",	--828
		x"38",	--829
		x"1d",	--830
		x"3a",	--831
		x"32",	--832
		x"0d",	--833
		x"1e",	--834
		x"0a",	--835
		x"02",	--836
		x"32",	--837
		x"03",	--838
		x"82",	--839
		x"32",	--840
		x"92",	--841
		x"04",	--842
		x"38",	--843
		x"1f",	--844
		x"3a",	--845
		x"32",	--846
		x"0f",	--847
		x"30",	--848
		x"0b",	--849
		x"0a",	--850
		x"21",	--851
		x"0a",	--852
		x"0b",	--853
		x"30",	--854
		x"2c",	--855
		x"b0",	--856
		x"b4",	--857
		x"21",	--858
		x"3a",	--859
		x"03",	--860
		x"1b",	--861
		x"0e",	--862
		x"1f",	--863
		x"02",	--864
		x"b0",	--865
		x"72",	--866
		x"0a",	--867
		x"0e",	--868
		x"1f",	--869
		x"04",	--870
		x"b0",	--871
		x"72",	--872
		x"0b",	--873
		x"0f",	--874
		x"0a",	--875
		x"30",	--876
		x"74",	--877
		x"b0",	--878
		x"b4",	--879
		x"31",	--880
		x"06",	--881
		x"8a",	--882
		x"00",	--883
		x"0f",	--884
		x"21",	--885
		x"3a",	--886
		x"3b",	--887
		x"30",	--888
		x"30",	--889
		x"34",	--890
		x"b0",	--891
		x"b4",	--892
		x"b1",	--893
		x"4e",	--894
		x"00",	--895
		x"b0",	--896
		x"b4",	--897
		x"a1",	--898
		x"00",	--899
		x"30",	--900
		x"5f",	--901
		x"b0",	--902
		x"b4",	--903
		x"21",	--904
		x"3f",	--905
		x"ea",	--906
		x"0b",	--907
		x"21",	--908
		x"0b",	--909
		x"1f",	--910
		x"17",	--911
		x"16",	--912
		x"30",	--913
		x"8f",	--914
		x"b0",	--915
		x"b4",	--916
		x"21",	--917
		x"0e",	--918
		x"1f",	--919
		x"02",	--920
		x"b0",	--921
		x"72",	--922
		x"2f",	--923
		x"0f",	--924
		x"30",	--925
		x"74",	--926
		x"b0",	--927
		x"b4",	--928
		x"31",	--929
		x"06",	--930
		x"0f",	--931
		x"21",	--932
		x"3b",	--933
		x"30",	--934
		x"30",	--935
		x"34",	--936
		x"b0",	--937
		x"b4",	--938
		x"b1",	--939
		x"4e",	--940
		x"00",	--941
		x"b0",	--942
		x"b4",	--943
		x"a1",	--944
		x"00",	--945
		x"30",	--946
		x"80",	--947
		x"b0",	--948
		x"b4",	--949
		x"21",	--950
		x"3f",	--951
		x"eb",	--952
		x"0b",	--953
		x"0a",	--954
		x"8e",	--955
		x"00",	--956
		x"6d",	--957
		x"4d",	--958
		x"5e",	--959
		x"1f",	--960
		x"0a",	--961
		x"0c",	--962
		x"0f",	--963
		x"7b",	--964
		x"0a",	--965
		x"2b",	--966
		x"0c",	--967
		x"0c",	--968
		x"0c",	--969
		x"0c",	--970
		x"8d",	--971
		x"0c",	--972
		x"3c",	--973
		x"d0",	--974
		x"1a",	--975
		x"7d",	--976
		x"4d",	--977
		x"17",	--978
		x"7d",	--979
		x"78",	--980
		x"1a",	--981
		x"4b",	--982
		x"7b",	--983
		x"d0",	--984
		x"0a",	--985
		x"e9",	--986
		x"7b",	--987
		x"0a",	--988
		x"34",	--989
		x"0c",	--990
		x"0b",	--991
		x"0b",	--992
		x"0b",	--993
		x"0c",	--994
		x"8d",	--995
		x"0c",	--996
		x"3c",	--997
		x"d0",	--998
		x"7d",	--999
		x"4d",	--1000
		x"e9",	--1001
		x"9e",	--1002
		x"00",	--1003
		x"0f",	--1004
		x"3a",	--1005
		x"3b",	--1006
		x"30",	--1007
		x"1a",	--1008
		x"de",	--1009
		x"4b",	--1010
		x"7b",	--1011
		x"9f",	--1012
		x"7b",	--1013
		x"06",	--1014
		x"0a",	--1015
		x"0c",	--1016
		x"0c",	--1017
		x"0c",	--1018
		x"0c",	--1019
		x"8d",	--1020
		x"0c",	--1021
		x"3c",	--1022
		x"a9",	--1023
		x"1a",	--1024
		x"ce",	--1025
		x"4b",	--1026
		x"7b",	--1027
		x"bf",	--1028
		x"7b",	--1029
		x"06",	--1030
		x"0a",	--1031
		x"0c",	--1032
		x"0c",	--1033
		x"0c",	--1034
		x"0c",	--1035
		x"8d",	--1036
		x"0c",	--1037
		x"3c",	--1038
		x"c9",	--1039
		x"1a",	--1040
		x"be",	--1041
		x"8d",	--1042
		x"0d",	--1043
		x"30",	--1044
		x"96",	--1045
		x"b0",	--1046
		x"b4",	--1047
		x"21",	--1048
		x"0c",	--1049
		x"0f",	--1050
		x"3a",	--1051
		x"3b",	--1052
		x"30",	--1053
		x"0c",	--1054
		x"ca",	--1055
		x"0b",	--1056
		x"0a",	--1057
		x"0b",	--1058
		x"0a",	--1059
		x"8f",	--1060
		x"00",	--1061
		x"8f",	--1062
		x"02",	--1063
		x"8f",	--1064
		x"04",	--1065
		x"0c",	--1066
		x"0d",	--1067
		x"3e",	--1068
		x"00",	--1069
		x"3f",	--1070
		x"6e",	--1071
		x"b0",	--1072
		x"8e",	--1073
		x"8b",	--1074
		x"02",	--1075
		x"02",	--1076
		x"32",	--1077
		x"03",	--1078
		x"82",	--1079
		x"32",	--1080
		x"b2",	--1081
		x"18",	--1082
		x"38",	--1083
		x"9b",	--1084
		x"3a",	--1085
		x"06",	--1086
		x"32",	--1087
		x"0f",	--1088
		x"3a",	--1089
		x"3b",	--1090
		x"30",	--1091
		x"0b",	--1092
		x"09",	--1093
		x"08",	--1094
		x"8f",	--1095
		x"06",	--1096
		x"bf",	--1097
		x"00",	--1098
		x"08",	--1099
		x"2b",	--1100
		x"1e",	--1101
		x"02",	--1102
		x"0f",	--1103
		x"b0",	--1104
		x"28",	--1105
		x"0c",	--1106
		x"3d",	--1107
		x"00",	--1108
		x"b0",	--1109
		x"d4",	--1110
		x"08",	--1111
		x"09",	--1112
		x"1e",	--1113
		x"06",	--1114
		x"0f",	--1115
		x"b0",	--1116
		x"28",	--1117
		x"0c",	--1118
		x"0d",	--1119
		x"0e",	--1120
		x"0f",	--1121
		x"b0",	--1122
		x"84",	--1123
		x"b0",	--1124
		x"64",	--1125
		x"8b",	--1126
		x"04",	--1127
		x"9b",	--1128
		x"00",	--1129
		x"38",	--1130
		x"39",	--1131
		x"3b",	--1132
		x"30",	--1133
		x"0b",	--1134
		x"0a",	--1135
		x"09",	--1136
		x"0a",	--1137
		x"0b",	--1138
		x"8f",	--1139
		x"06",	--1140
		x"8f",	--1141
		x"08",	--1142
		x"29",	--1143
		x"1e",	--1144
		x"02",	--1145
		x"0f",	--1146
		x"b0",	--1147
		x"28",	--1148
		x"0c",	--1149
		x"0d",	--1150
		x"0e",	--1151
		x"0f",	--1152
		x"b0",	--1153
		x"d4",	--1154
		x"0a",	--1155
		x"0b",	--1156
		x"1e",	--1157
		x"06",	--1158
		x"0f",	--1159
		x"b0",	--1160
		x"28",	--1161
		x"0c",	--1162
		x"0d",	--1163
		x"0e",	--1164
		x"0f",	--1165
		x"b0",	--1166
		x"84",	--1167
		x"b0",	--1168
		x"64",	--1169
		x"89",	--1170
		x"04",	--1171
		x"39",	--1172
		x"3a",	--1173
		x"3b",	--1174
		x"30",	--1175
		x"2f",	--1176
		x"8f",	--1177
		x"04",	--1178
		x"30",	--1179
		x"0b",	--1180
		x"0a",	--1181
		x"92",	--1182
		x"12",	--1183
		x"14",	--1184
		x"3b",	--1185
		x"6c",	--1186
		x"0a",	--1187
		x"2b",	--1188
		x"5f",	--1189
		x"fc",	--1190
		x"8f",	--1191
		x"0f",	--1192
		x"30",	--1193
		x"ab",	--1194
		x"b0",	--1195
		x"b4",	--1196
		x"31",	--1197
		x"06",	--1198
		x"1a",	--1199
		x"3b",	--1200
		x"06",	--1201
		x"1a",	--1202
		x"12",	--1203
		x"ef",	--1204
		x"0f",	--1205
		x"3a",	--1206
		x"3b",	--1207
		x"30",	--1208
		x"1e",	--1209
		x"12",	--1210
		x"3e",	--1211
		x"20",	--1212
		x"12",	--1213
		x"0f",	--1214
		x"0f",	--1215
		x"0f",	--1216
		x"0f",	--1217
		x"3f",	--1218
		x"68",	--1219
		x"ff",	--1220
		x"68",	--1221
		x"00",	--1222
		x"bf",	--1223
		x"38",	--1224
		x"02",	--1225
		x"bf",	--1226
		x"04",	--1227
		x"04",	--1228
		x"1e",	--1229
		x"82",	--1230
		x"12",	--1231
		x"30",	--1232
		x"0b",	--1233
		x"1b",	--1234
		x"12",	--1235
		x"3b",	--1236
		x"20",	--1237
		x"12",	--1238
		x"0c",	--1239
		x"0c",	--1240
		x"0c",	--1241
		x"0c",	--1242
		x"3c",	--1243
		x"68",	--1244
		x"cc",	--1245
		x"00",	--1246
		x"8c",	--1247
		x"02",	--1248
		x"8c",	--1249
		x"04",	--1250
		x"1b",	--1251
		x"82",	--1252
		x"12",	--1253
		x"0f",	--1254
		x"3b",	--1255
		x"30",	--1256
		x"3f",	--1257
		x"fc",	--1258
		x"0b",	--1259
		x"31",	--1260
		x"f0",	--1261
		x"1b",	--1262
		x"12",	--1263
		x"1b",	--1264
		x"0f",	--1265
		x"5f",	--1266
		x"68",	--1267
		x"16",	--1268
		x"3d",	--1269
		x"6e",	--1270
		x"0c",	--1271
		x"05",	--1272
		x"3d",	--1273
		x"06",	--1274
		x"cd",	--1275
		x"fa",	--1276
		x"0e",	--1277
		x"1c",	--1278
		x"0c",	--1279
		x"f8",	--1280
		x"30",	--1281
		x"b3",	--1282
		x"b0",	--1283
		x"b4",	--1284
		x"21",	--1285
		x"3f",	--1286
		x"31",	--1287
		x"10",	--1288
		x"3b",	--1289
		x"30",	--1290
		x"0c",	--1291
		x"81",	--1292
		x"00",	--1293
		x"6d",	--1294
		x"4d",	--1295
		x"24",	--1296
		x"1e",	--1297
		x"1f",	--1298
		x"06",	--1299
		x"6d",	--1300
		x"4d",	--1301
		x"11",	--1302
		x"1e",	--1303
		x"3f",	--1304
		x"0e",	--1305
		x"7d",	--1306
		x"20",	--1307
		x"f7",	--1308
		x"ce",	--1309
		x"ff",	--1310
		x"0d",	--1311
		x"0d",	--1312
		x"0d",	--1313
		x"8d",	--1314
		x"00",	--1315
		x"1f",	--1316
		x"6d",	--1317
		x"4d",	--1318
		x"ef",	--1319
		x"0e",	--1320
		x"0e",	--1321
		x"0c",	--1322
		x"0c",	--1323
		x"3c",	--1324
		x"68",	--1325
		x"0e",	--1326
		x"9c",	--1327
		x"02",	--1328
		x"31",	--1329
		x"10",	--1330
		x"3b",	--1331
		x"30",	--1332
		x"1f",	--1333
		x"f1",	--1334
		x"b2",	--1335
		x"d2",	--1336
		x"60",	--1337
		x"b2",	--1338
		x"b8",	--1339
		x"72",	--1340
		x"0f",	--1341
		x"30",	--1342
		x"0b",	--1343
		x"0b",	--1344
		x"1f",	--1345
		x"14",	--1346
		x"3f",	--1347
		x"20",	--1348
		x"19",	--1349
		x"0c",	--1350
		x"0c",	--1351
		x"0d",	--1352
		x"0d",	--1353
		x"0d",	--1354
		x"0d",	--1355
		x"0d",	--1356
		x"3d",	--1357
		x"28",	--1358
		x"8d",	--1359
		x"00",	--1360
		x"8d",	--1361
		x"02",	--1362
		x"8d",	--1363
		x"08",	--1364
		x"8d",	--1365
		x"0a",	--1366
		x"8d",	--1367
		x"0c",	--1368
		x"0e",	--1369
		x"1e",	--1370
		x"82",	--1371
		x"14",	--1372
		x"3b",	--1373
		x"30",	--1374
		x"3f",	--1375
		x"fc",	--1376
		x"0f",	--1377
		x"0c",	--1378
		x"0c",	--1379
		x"0c",	--1380
		x"0c",	--1381
		x"0c",	--1382
		x"3c",	--1383
		x"28",	--1384
		x"8c",	--1385
		x"02",	--1386
		x"8c",	--1387
		x"04",	--1388
		x"8c",	--1389
		x"06",	--1390
		x"8c",	--1391
		x"08",	--1392
		x"9c",	--1393
		x"00",	--1394
		x"0f",	--1395
		x"30",	--1396
		x"0f",	--1397
		x"0e",	--1398
		x"0e",	--1399
		x"0e",	--1400
		x"0e",	--1401
		x"0e",	--1402
		x"8e",	--1403
		x"28",	--1404
		x"0f",	--1405
		x"30",	--1406
		x"0f",	--1407
		x"0e",	--1408
		x"0d",	--1409
		x"0c",	--1410
		x"0b",	--1411
		x"0a",	--1412
		x"09",	--1413
		x"08",	--1414
		x"07",	--1415
		x"92",	--1416
		x"14",	--1417
		x"33",	--1418
		x"3a",	--1419
		x"28",	--1420
		x"0b",	--1421
		x"2b",	--1422
		x"08",	--1423
		x"38",	--1424
		x"07",	--1425
		x"37",	--1426
		x"06",	--1427
		x"09",	--1428
		x"0f",	--1429
		x"1f",	--1430
		x"8b",	--1431
		x"00",	--1432
		x"19",	--1433
		x"3a",	--1434
		x"0e",	--1435
		x"3b",	--1436
		x"0e",	--1437
		x"38",	--1438
		x"0e",	--1439
		x"37",	--1440
		x"0e",	--1441
		x"19",	--1442
		x"14",	--1443
		x"19",	--1444
		x"8a",	--1445
		x"00",	--1446
		x"f1",	--1447
		x"2f",	--1448
		x"1f",	--1449
		x"02",	--1450
		x"ea",	--1451
		x"8b",	--1452
		x"00",	--1453
		x"1f",	--1454
		x"0a",	--1455
		x"9b",	--1456
		x"08",	--1457
		x"88",	--1458
		x"00",	--1459
		x"e4",	--1460
		x"2f",	--1461
		x"1f",	--1462
		x"87",	--1463
		x"00",	--1464
		x"2f",	--1465
		x"de",	--1466
		x"8a",	--1467
		x"00",	--1468
		x"db",	--1469
		x"b2",	--1470
		x"fe",	--1471
		x"60",	--1472
		x"37",	--1473
		x"38",	--1474
		x"39",	--1475
		x"3a",	--1476
		x"3b",	--1477
		x"3c",	--1478
		x"3d",	--1479
		x"3e",	--1480
		x"3f",	--1481
		x"00",	--1482
		x"8f",	--1483
		x"00",	--1484
		x"0f",	--1485
		x"30",	--1486
		x"2f",	--1487
		x"2e",	--1488
		x"1f",	--1489
		x"02",	--1490
		x"30",	--1491
		x"8f",	--1492
		x"00",	--1493
		x"30",	--1494
		x"8f",	--1495
		x"00",	--1496
		x"3f",	--1497
		x"a8",	--1498
		x"b0",	--1499
		x"7e",	--1500
		x"82",	--1501
		x"0a",	--1502
		x"0f",	--1503
		x"30",	--1504
		x"0c",	--1505
		x"2f",	--1506
		x"8f",	--1507
		x"00",	--1508
		x"1d",	--1509
		x"0e",	--1510
		x"1f",	--1511
		x"0a",	--1512
		x"b0",	--1513
		x"c2",	--1514
		x"30",	--1515
		x"5e",	--1516
		x"81",	--1517
		x"3e",	--1518
		x"fc",	--1519
		x"c2",	--1520
		x"84",	--1521
		x"0f",	--1522
		x"30",	--1523
		x"3f",	--1524
		x"0f",	--1525
		x"5f",	--1526
		x"72",	--1527
		x"8f",	--1528
		x"b0",	--1529
		x"d8",	--1530
		x"30",	--1531
		x"0b",	--1532
		x"0b",	--1533
		x"0e",	--1534
		x"0e",	--1535
		x"0e",	--1536
		x"0e",	--1537
		x"0e",	--1538
		x"0f",	--1539
		x"b0",	--1540
		x"e8",	--1541
		x"0f",	--1542
		x"b0",	--1543
		x"e8",	--1544
		x"3b",	--1545
		x"30",	--1546
		x"0b",	--1547
		x"0a",	--1548
		x"0a",	--1549
		x"3b",	--1550
		x"07",	--1551
		x"0e",	--1552
		x"4d",	--1553
		x"7d",	--1554
		x"0f",	--1555
		x"03",	--1556
		x"0e",	--1557
		x"7d",	--1558
		x"fd",	--1559
		x"1e",	--1560
		x"0a",	--1561
		x"3f",	--1562
		x"31",	--1563
		x"b0",	--1564
		x"d8",	--1565
		x"3b",	--1566
		x"3b",	--1567
		x"ef",	--1568
		x"3a",	--1569
		x"3b",	--1570
		x"30",	--1571
		x"3f",	--1572
		x"30",	--1573
		x"f5",	--1574
		x"0b",	--1575
		x"0b",	--1576
		x"0e",	--1577
		x"8e",	--1578
		x"8e",	--1579
		x"0f",	--1580
		x"b0",	--1581
		x"f8",	--1582
		x"0f",	--1583
		x"b0",	--1584
		x"f8",	--1585
		x"3b",	--1586
		x"30",	--1587
		x"0b",	--1588
		x"0a",	--1589
		x"0a",	--1590
		x"0b",	--1591
		x"0d",	--1592
		x"8d",	--1593
		x"8d",	--1594
		x"0f",	--1595
		x"b0",	--1596
		x"f8",	--1597
		x"0f",	--1598
		x"b0",	--1599
		x"f8",	--1600
		x"0c",	--1601
		x"0d",	--1602
		x"8d",	--1603
		x"8c",	--1604
		x"4d",	--1605
		x"0d",	--1606
		x"0f",	--1607
		x"b0",	--1608
		x"f8",	--1609
		x"0f",	--1610
		x"b0",	--1611
		x"f8",	--1612
		x"3a",	--1613
		x"3b",	--1614
		x"30",	--1615
		x"0b",	--1616
		x"0a",	--1617
		x"09",	--1618
		x"0a",	--1619
		x"0e",	--1620
		x"19",	--1621
		x"09",	--1622
		x"39",	--1623
		x"0b",	--1624
		x"0d",	--1625
		x"0d",	--1626
		x"6f",	--1627
		x"8f",	--1628
		x"b0",	--1629
		x"f8",	--1630
		x"0b",	--1631
		x"0e",	--1632
		x"1b",	--1633
		x"3b",	--1634
		x"07",	--1635
		x"05",	--1636
		x"3f",	--1637
		x"20",	--1638
		x"b0",	--1639
		x"d8",	--1640
		x"ef",	--1641
		x"3f",	--1642
		x"3a",	--1643
		x"b0",	--1644
		x"d8",	--1645
		x"ea",	--1646
		x"39",	--1647
		x"3a",	--1648
		x"3b",	--1649
		x"30",	--1650
		x"0b",	--1651
		x"0a",	--1652
		x"09",	--1653
		x"0a",	--1654
		x"0e",	--1655
		x"17",	--1656
		x"09",	--1657
		x"39",	--1658
		x"0b",	--1659
		x"6f",	--1660
		x"8f",	--1661
		x"b0",	--1662
		x"e8",	--1663
		x"0b",	--1664
		x"0e",	--1665
		x"1b",	--1666
		x"3b",	--1667
		x"07",	--1668
		x"f6",	--1669
		x"3f",	--1670
		x"20",	--1671
		x"b0",	--1672
		x"d8",	--1673
		x"6f",	--1674
		x"8f",	--1675
		x"b0",	--1676
		x"e8",	--1677
		x"0b",	--1678
		x"f2",	--1679
		x"39",	--1680
		x"3a",	--1681
		x"3b",	--1682
		x"30",	--1683
		x"0b",	--1684
		x"0a",	--1685
		x"09",	--1686
		x"31",	--1687
		x"ec",	--1688
		x"0b",	--1689
		x"0f",	--1690
		x"34",	--1691
		x"3b",	--1692
		x"0a",	--1693
		x"38",	--1694
		x"09",	--1695
		x"0a",	--1696
		x"0a",	--1697
		x"3e",	--1698
		x"0a",	--1699
		x"0f",	--1700
		x"b0",	--1701
		x"46",	--1702
		x"7f",	--1703
		x"30",	--1704
		x"ca",	--1705
		x"00",	--1706
		x"19",	--1707
		x"3e",	--1708
		x"0a",	--1709
		x"0f",	--1710
		x"b0",	--1711
		x"14",	--1712
		x"0b",	--1713
		x"3f",	--1714
		x"0a",	--1715
		x"eb",	--1716
		x"0a",	--1717
		x"1a",	--1718
		x"09",	--1719
		x"3e",	--1720
		x"0a",	--1721
		x"0f",	--1722
		x"b0",	--1723
		x"46",	--1724
		x"7f",	--1725
		x"30",	--1726
		x"c9",	--1727
		x"00",	--1728
		x"3a",	--1729
		x"0f",	--1730
		x"0f",	--1731
		x"6f",	--1732
		x"8f",	--1733
		x"b0",	--1734
		x"d8",	--1735
		x"0a",	--1736
		x"f7",	--1737
		x"31",	--1738
		x"14",	--1739
		x"39",	--1740
		x"3a",	--1741
		x"3b",	--1742
		x"30",	--1743
		x"3f",	--1744
		x"2d",	--1745
		x"b0",	--1746
		x"d8",	--1747
		x"3b",	--1748
		x"1b",	--1749
		x"c5",	--1750
		x"1a",	--1751
		x"09",	--1752
		x"dd",	--1753
		x"0b",	--1754
		x"0a",	--1755
		x"09",	--1756
		x"0b",	--1757
		x"3b",	--1758
		x"39",	--1759
		x"6f",	--1760
		x"4f",	--1761
		x"0b",	--1762
		x"1a",	--1763
		x"8f",	--1764
		x"b0",	--1765
		x"d8",	--1766
		x"0a",	--1767
		x"09",	--1768
		x"19",	--1769
		x"5f",	--1770
		x"01",	--1771
		x"4f",	--1772
		x"10",	--1773
		x"7f",	--1774
		x"25",	--1775
		x"f3",	--1776
		x"0a",	--1777
		x"1a",	--1778
		x"5f",	--1779
		x"01",	--1780
		x"7f",	--1781
		x"db",	--1782
		x"7f",	--1783
		x"54",	--1784
		x"ee",	--1785
		x"4f",	--1786
		x"0f",	--1787
		x"10",	--1788
		x"ca",	--1789
		x"39",	--1790
		x"3a",	--1791
		x"3b",	--1792
		x"30",	--1793
		x"09",	--1794
		x"29",	--1795
		x"1e",	--1796
		x"02",	--1797
		x"2f",	--1798
		x"b0",	--1799
		x"a0",	--1800
		x"0b",	--1801
		x"dd",	--1802
		x"09",	--1803
		x"29",	--1804
		x"2f",	--1805
		x"b0",	--1806
		x"4e",	--1807
		x"0b",	--1808
		x"d6",	--1809
		x"0f",	--1810
		x"2b",	--1811
		x"29",	--1812
		x"6f",	--1813
		x"4f",	--1814
		x"d0",	--1815
		x"19",	--1816
		x"8f",	--1817
		x"b0",	--1818
		x"d8",	--1819
		x"7f",	--1820
		x"4f",	--1821
		x"fa",	--1822
		x"c8",	--1823
		x"09",	--1824
		x"29",	--1825
		x"1e",	--1826
		x"02",	--1827
		x"2f",	--1828
		x"b0",	--1829
		x"e6",	--1830
		x"0b",	--1831
		x"bf",	--1832
		x"09",	--1833
		x"29",	--1834
		x"2e",	--1835
		x"0f",	--1836
		x"8f",	--1837
		x"8f",	--1838
		x"8f",	--1839
		x"8f",	--1840
		x"b0",	--1841
		x"68",	--1842
		x"0b",	--1843
		x"b3",	--1844
		x"09",	--1845
		x"29",	--1846
		x"2f",	--1847
		x"b0",	--1848
		x"28",	--1849
		x"0b",	--1850
		x"ac",	--1851
		x"09",	--1852
		x"29",	--1853
		x"2f",	--1854
		x"b0",	--1855
		x"d8",	--1856
		x"0b",	--1857
		x"a5",	--1858
		x"09",	--1859
		x"29",	--1860
		x"2f",	--1861
		x"b0",	--1862
		x"f8",	--1863
		x"0b",	--1864
		x"9e",	--1865
		x"09",	--1866
		x"29",	--1867
		x"2f",	--1868
		x"b0",	--1869
		x"16",	--1870
		x"0b",	--1871
		x"97",	--1872
		x"3f",	--1873
		x"25",	--1874
		x"b0",	--1875
		x"d8",	--1876
		x"92",	--1877
		x"0f",	--1878
		x"0e",	--1879
		x"1f",	--1880
		x"16",	--1881
		x"df",	--1882
		x"85",	--1883
		x"e8",	--1884
		x"1f",	--1885
		x"16",	--1886
		x"3f",	--1887
		x"3f",	--1888
		x"13",	--1889
		x"92",	--1890
		x"16",	--1891
		x"1e",	--1892
		x"16",	--1893
		x"1f",	--1894
		x"18",	--1895
		x"0e",	--1896
		x"02",	--1897
		x"92",	--1898
		x"18",	--1899
		x"f2",	--1900
		x"10",	--1901
		x"81",	--1902
		x"3e",	--1903
		x"3f",	--1904
		x"b1",	--1905
		x"f0",	--1906
		x"00",	--1907
		x"00",	--1908
		x"82",	--1909
		x"16",	--1910
		x"ec",	--1911
		x"0c",	--1912
		x"0d",	--1913
		x"3e",	--1914
		x"00",	--1915
		x"3f",	--1916
		x"6e",	--1917
		x"b0",	--1918
		x"4e",	--1919
		x"3e",	--1920
		x"82",	--1921
		x"82",	--1922
		x"f2",	--1923
		x"11",	--1924
		x"80",	--1925
		x"30",	--1926
		x"1e",	--1927
		x"16",	--1928
		x"1f",	--1929
		x"18",	--1930
		x"0e",	--1931
		x"05",	--1932
		x"1f",	--1933
		x"16",	--1934
		x"1f",	--1935
		x"18",	--1936
		x"30",	--1937
		x"1d",	--1938
		x"16",	--1939
		x"1e",	--1940
		x"18",	--1941
		x"3f",	--1942
		x"40",	--1943
		x"0f",	--1944
		x"0f",	--1945
		x"30",	--1946
		x"1f",	--1947
		x"18",	--1948
		x"5f",	--1949
		x"e8",	--1950
		x"1d",	--1951
		x"18",	--1952
		x"1e",	--1953
		x"16",	--1954
		x"0d",	--1955
		x"0b",	--1956
		x"1e",	--1957
		x"18",	--1958
		x"3e",	--1959
		x"3f",	--1960
		x"03",	--1961
		x"82",	--1962
		x"18",	--1963
		x"30",	--1964
		x"92",	--1965
		x"18",	--1966
		x"30",	--1967
		x"4f",	--1968
		x"30",	--1969
		x"0b",	--1970
		x"0a",	--1971
		x"0a",	--1972
		x"0b",	--1973
		x"0c",	--1974
		x"3d",	--1975
		x"00",	--1976
		x"b0",	--1977
		x"48",	--1978
		x"0f",	--1979
		x"07",	--1980
		x"0e",	--1981
		x"0f",	--1982
		x"b0",	--1983
		x"98",	--1984
		x"3a",	--1985
		x"3b",	--1986
		x"30",	--1987
		x"0c",	--1988
		x"3d",	--1989
		x"00",	--1990
		x"0e",	--1991
		x"0f",	--1992
		x"b0",	--1993
		x"84",	--1994
		x"b0",	--1995
		x"98",	--1996
		x"0e",	--1997
		x"3f",	--1998
		x"00",	--1999
		x"3a",	--2000
		x"3b",	--2001
		x"30",	--2002
		x"0b",	--2003
		x"0a",	--2004
		x"09",	--2005
		x"08",	--2006
		x"07",	--2007
		x"06",	--2008
		x"05",	--2009
		x"04",	--2010
		x"31",	--2011
		x"fa",	--2012
		x"08",	--2013
		x"6b",	--2014
		x"6b",	--2015
		x"67",	--2016
		x"6c",	--2017
		x"6c",	--2018
		x"e9",	--2019
		x"6b",	--2020
		x"02",	--2021
		x"30",	--2022
		x"26",	--2023
		x"6c",	--2024
		x"e3",	--2025
		x"6c",	--2026
		x"bb",	--2027
		x"6b",	--2028
		x"df",	--2029
		x"91",	--2030
		x"02",	--2031
		x"00",	--2032
		x"1b",	--2033
		x"02",	--2034
		x"14",	--2035
		x"04",	--2036
		x"15",	--2037
		x"06",	--2038
		x"16",	--2039
		x"04",	--2040
		x"17",	--2041
		x"06",	--2042
		x"2c",	--2043
		x"0c",	--2044
		x"09",	--2045
		x"0c",	--2046
		x"bf",	--2047
		x"39",	--2048
		x"20",	--2049
		x"50",	--2050
		x"1c",	--2051
		x"d7",	--2052
		x"81",	--2053
		x"02",	--2054
		x"81",	--2055
		x"04",	--2056
		x"4c",	--2057
		x"7c",	--2058
		x"1f",	--2059
		x"0b",	--2060
		x"0a",	--2061
		x"0b",	--2062
		x"12",	--2063
		x"0b",	--2064
		x"0a",	--2065
		x"7c",	--2066
		x"fb",	--2067
		x"81",	--2068
		x"02",	--2069
		x"81",	--2070
		x"04",	--2071
		x"1c",	--2072
		x"0d",	--2073
		x"79",	--2074
		x"1f",	--2075
		x"04",	--2076
		x"0c",	--2077
		x"0d",	--2078
		x"79",	--2079
		x"fc",	--2080
		x"3c",	--2081
		x"3d",	--2082
		x"0c",	--2083
		x"0d",	--2084
		x"1a",	--2085
		x"0b",	--2086
		x"0c",	--2087
		x"02",	--2088
		x"0d",	--2089
		x"e5",	--2090
		x"16",	--2091
		x"02",	--2092
		x"17",	--2093
		x"04",	--2094
		x"06",	--2095
		x"07",	--2096
		x"5f",	--2097
		x"01",	--2098
		x"5f",	--2099
		x"01",	--2100
		x"28",	--2101
		x"c8",	--2102
		x"01",	--2103
		x"a8",	--2104
		x"02",	--2105
		x"0e",	--2106
		x"0f",	--2107
		x"0e",	--2108
		x"0f",	--2109
		x"88",	--2110
		x"04",	--2111
		x"88",	--2112
		x"06",	--2113
		x"f8",	--2114
		x"03",	--2115
		x"00",	--2116
		x"0f",	--2117
		x"4d",	--2118
		x"0f",	--2119
		x"31",	--2120
		x"06",	--2121
		x"34",	--2122
		x"35",	--2123
		x"36",	--2124
		x"37",	--2125
		x"38",	--2126
		x"39",	--2127
		x"3a",	--2128
		x"3b",	--2129
		x"30",	--2130
		x"2b",	--2131
		x"67",	--2132
		x"81",	--2133
		x"00",	--2134
		x"04",	--2135
		x"05",	--2136
		x"5f",	--2137
		x"01",	--2138
		x"5f",	--2139
		x"01",	--2140
		x"d8",	--2141
		x"4f",	--2142
		x"68",	--2143
		x"0e",	--2144
		x"0f",	--2145
		x"0e",	--2146
		x"0f",	--2147
		x"0f",	--2148
		x"69",	--2149
		x"c8",	--2150
		x"01",	--2151
		x"a8",	--2152
		x"02",	--2153
		x"88",	--2154
		x"04",	--2155
		x"88",	--2156
		x"06",	--2157
		x"0c",	--2158
		x"0d",	--2159
		x"3c",	--2160
		x"3d",	--2161
		x"3d",	--2162
		x"ff",	--2163
		x"05",	--2164
		x"3d",	--2165
		x"00",	--2166
		x"17",	--2167
		x"3c",	--2168
		x"15",	--2169
		x"1b",	--2170
		x"02",	--2171
		x"3b",	--2172
		x"0e",	--2173
		x"0f",	--2174
		x"0a",	--2175
		x"3b",	--2176
		x"0c",	--2177
		x"0d",	--2178
		x"3c",	--2179
		x"3d",	--2180
		x"3d",	--2181
		x"ff",	--2182
		x"f5",	--2183
		x"3c",	--2184
		x"88",	--2185
		x"04",	--2186
		x"88",	--2187
		x"06",	--2188
		x"88",	--2189
		x"02",	--2190
		x"f8",	--2191
		x"03",	--2192
		x"00",	--2193
		x"0f",	--2194
		x"b3",	--2195
		x"0c",	--2196
		x"0d",	--2197
		x"1c",	--2198
		x"0d",	--2199
		x"12",	--2200
		x"0f",	--2201
		x"0e",	--2202
		x"0a",	--2203
		x"0b",	--2204
		x"0a",	--2205
		x"0b",	--2206
		x"88",	--2207
		x"04",	--2208
		x"88",	--2209
		x"06",	--2210
		x"98",	--2211
		x"02",	--2212
		x"0f",	--2213
		x"a1",	--2214
		x"6b",	--2215
		x"9f",	--2216
		x"ad",	--2217
		x"00",	--2218
		x"9d",	--2219
		x"02",	--2220
		x"02",	--2221
		x"9d",	--2222
		x"04",	--2223
		x"04",	--2224
		x"9d",	--2225
		x"06",	--2226
		x"06",	--2227
		x"5e",	--2228
		x"01",	--2229
		x"5e",	--2230
		x"01",	--2231
		x"cd",	--2232
		x"01",	--2233
		x"0f",	--2234
		x"8c",	--2235
		x"06",	--2236
		x"07",	--2237
		x"9a",	--2238
		x"39",	--2239
		x"19",	--2240
		x"39",	--2241
		x"20",	--2242
		x"8f",	--2243
		x"3e",	--2244
		x"3c",	--2245
		x"b6",	--2246
		x"c1",	--2247
		x"0e",	--2248
		x"0f",	--2249
		x"0e",	--2250
		x"0f",	--2251
		x"97",	--2252
		x"0f",	--2253
		x"79",	--2254
		x"d8",	--2255
		x"01",	--2256
		x"a8",	--2257
		x"02",	--2258
		x"3e",	--2259
		x"3f",	--2260
		x"1e",	--2261
		x"0f",	--2262
		x"88",	--2263
		x"04",	--2264
		x"88",	--2265
		x"06",	--2266
		x"92",	--2267
		x"0c",	--2268
		x"7b",	--2269
		x"81",	--2270
		x"00",	--2271
		x"81",	--2272
		x"02",	--2273
		x"81",	--2274
		x"04",	--2275
		x"4d",	--2276
		x"7d",	--2277
		x"1f",	--2278
		x"0c",	--2279
		x"4b",	--2280
		x"0c",	--2281
		x"0d",	--2282
		x"12",	--2283
		x"0d",	--2284
		x"0c",	--2285
		x"7b",	--2286
		x"fb",	--2287
		x"81",	--2288
		x"02",	--2289
		x"81",	--2290
		x"04",	--2291
		x"1c",	--2292
		x"0d",	--2293
		x"79",	--2294
		x"1f",	--2295
		x"04",	--2296
		x"0c",	--2297
		x"0d",	--2298
		x"79",	--2299
		x"fc",	--2300
		x"3c",	--2301
		x"3d",	--2302
		x"0c",	--2303
		x"0d",	--2304
		x"1a",	--2305
		x"0b",	--2306
		x"0c",	--2307
		x"04",	--2308
		x"0d",	--2309
		x"02",	--2310
		x"0a",	--2311
		x"0b",	--2312
		x"14",	--2313
		x"02",	--2314
		x"15",	--2315
		x"04",	--2316
		x"04",	--2317
		x"05",	--2318
		x"49",	--2319
		x"0a",	--2320
		x"0b",	--2321
		x"18",	--2322
		x"6c",	--2323
		x"33",	--2324
		x"df",	--2325
		x"01",	--2326
		x"01",	--2327
		x"2f",	--2328
		x"3f",	--2329
		x"84",	--2330
		x"2c",	--2331
		x"31",	--2332
		x"e0",	--2333
		x"81",	--2334
		x"04",	--2335
		x"81",	--2336
		x"06",	--2337
		x"81",	--2338
		x"00",	--2339
		x"81",	--2340
		x"02",	--2341
		x"0e",	--2342
		x"3e",	--2343
		x"18",	--2344
		x"0f",	--2345
		x"2f",	--2346
		x"b0",	--2347
		x"5a",	--2348
		x"0e",	--2349
		x"3e",	--2350
		x"10",	--2351
		x"0f",	--2352
		x"b0",	--2353
		x"5a",	--2354
		x"0d",	--2355
		x"3d",	--2356
		x"0e",	--2357
		x"3e",	--2358
		x"10",	--2359
		x"0f",	--2360
		x"3f",	--2361
		x"18",	--2362
		x"b0",	--2363
		x"a6",	--2364
		x"b0",	--2365
		x"7c",	--2366
		x"31",	--2367
		x"20",	--2368
		x"30",	--2369
		x"31",	--2370
		x"e0",	--2371
		x"81",	--2372
		x"04",	--2373
		x"81",	--2374
		x"06",	--2375
		x"81",	--2376
		x"00",	--2377
		x"81",	--2378
		x"02",	--2379
		x"0e",	--2380
		x"3e",	--2381
		x"18",	--2382
		x"0f",	--2383
		x"2f",	--2384
		x"b0",	--2385
		x"5a",	--2386
		x"0e",	--2387
		x"3e",	--2388
		x"10",	--2389
		x"0f",	--2390
		x"b0",	--2391
		x"5a",	--2392
		x"d1",	--2393
		x"11",	--2394
		x"0d",	--2395
		x"3d",	--2396
		x"0e",	--2397
		x"3e",	--2398
		x"10",	--2399
		x"0f",	--2400
		x"3f",	--2401
		x"18",	--2402
		x"b0",	--2403
		x"a6",	--2404
		x"b0",	--2405
		x"7c",	--2406
		x"31",	--2407
		x"20",	--2408
		x"30",	--2409
		x"0b",	--2410
		x"0a",	--2411
		x"09",	--2412
		x"08",	--2413
		x"07",	--2414
		x"06",	--2415
		x"05",	--2416
		x"04",	--2417
		x"31",	--2418
		x"dc",	--2419
		x"81",	--2420
		x"04",	--2421
		x"81",	--2422
		x"06",	--2423
		x"81",	--2424
		x"00",	--2425
		x"81",	--2426
		x"02",	--2427
		x"0e",	--2428
		x"3e",	--2429
		x"18",	--2430
		x"0f",	--2431
		x"2f",	--2432
		x"b0",	--2433
		x"5a",	--2434
		x"0e",	--2435
		x"3e",	--2436
		x"10",	--2437
		x"0f",	--2438
		x"b0",	--2439
		x"5a",	--2440
		x"5f",	--2441
		x"18",	--2442
		x"6f",	--2443
		x"b6",	--2444
		x"5e",	--2445
		x"10",	--2446
		x"6e",	--2447
		x"d9",	--2448
		x"6f",	--2449
		x"ae",	--2450
		x"6e",	--2451
		x"e2",	--2452
		x"6f",	--2453
		x"ac",	--2454
		x"6e",	--2455
		x"d1",	--2456
		x"14",	--2457
		x"1c",	--2458
		x"15",	--2459
		x"1e",	--2460
		x"18",	--2461
		x"14",	--2462
		x"19",	--2463
		x"16",	--2464
		x"3c",	--2465
		x"20",	--2466
		x"0e",	--2467
		x"0f",	--2468
		x"06",	--2469
		x"07",	--2470
		x"81",	--2471
		x"20",	--2472
		x"81",	--2473
		x"22",	--2474
		x"0a",	--2475
		x"0b",	--2476
		x"81",	--2477
		x"20",	--2478
		x"08",	--2479
		x"08",	--2480
		x"09",	--2481
		x"12",	--2482
		x"05",	--2483
		x"04",	--2484
		x"b1",	--2485
		x"20",	--2486
		x"19",	--2487
		x"14",	--2488
		x"0d",	--2489
		x"0a",	--2490
		x"0b",	--2491
		x"0e",	--2492
		x"0f",	--2493
		x"1c",	--2494
		x"0d",	--2495
		x"0b",	--2496
		x"03",	--2497
		x"0b",	--2498
		x"0c",	--2499
		x"0d",	--2500
		x"0e",	--2501
		x"0f",	--2502
		x"06",	--2503
		x"07",	--2504
		x"09",	--2505
		x"e5",	--2506
		x"16",	--2507
		x"07",	--2508
		x"e2",	--2509
		x"0a",	--2510
		x"f5",	--2511
		x"f2",	--2512
		x"81",	--2513
		x"20",	--2514
		x"81",	--2515
		x"22",	--2516
		x"0c",	--2517
		x"1a",	--2518
		x"1a",	--2519
		x"1a",	--2520
		x"12",	--2521
		x"06",	--2522
		x"26",	--2523
		x"81",	--2524
		x"0a",	--2525
		x"5d",	--2526
		x"d1",	--2527
		x"11",	--2528
		x"19",	--2529
		x"83",	--2530
		x"c1",	--2531
		x"09",	--2532
		x"0c",	--2533
		x"3c",	--2534
		x"3f",	--2535
		x"00",	--2536
		x"18",	--2537
		x"1d",	--2538
		x"0a",	--2539
		x"3d",	--2540
		x"1a",	--2541
		x"20",	--2542
		x"1b",	--2543
		x"22",	--2544
		x"0c",	--2545
		x"0e",	--2546
		x"0f",	--2547
		x"0b",	--2548
		x"2a",	--2549
		x"0a",	--2550
		x"0b",	--2551
		x"3d",	--2552
		x"3f",	--2553
		x"00",	--2554
		x"f5",	--2555
		x"81",	--2556
		x"20",	--2557
		x"81",	--2558
		x"22",	--2559
		x"81",	--2560
		x"0a",	--2561
		x"0c",	--2562
		x"0d",	--2563
		x"3c",	--2564
		x"7f",	--2565
		x"0d",	--2566
		x"3c",	--2567
		x"40",	--2568
		x"44",	--2569
		x"81",	--2570
		x"0c",	--2571
		x"81",	--2572
		x"0e",	--2573
		x"f1",	--2574
		x"03",	--2575
		x"08",	--2576
		x"0f",	--2577
		x"3f",	--2578
		x"b0",	--2579
		x"7c",	--2580
		x"31",	--2581
		x"24",	--2582
		x"34",	--2583
		x"35",	--2584
		x"36",	--2585
		x"37",	--2586
		x"38",	--2587
		x"39",	--2588
		x"3a",	--2589
		x"3b",	--2590
		x"30",	--2591
		x"1e",	--2592
		x"0f",	--2593
		x"d3",	--2594
		x"3a",	--2595
		x"03",	--2596
		x"08",	--2597
		x"1e",	--2598
		x"10",	--2599
		x"1c",	--2600
		x"20",	--2601
		x"1d",	--2602
		x"22",	--2603
		x"12",	--2604
		x"0d",	--2605
		x"0c",	--2606
		x"06",	--2607
		x"07",	--2608
		x"06",	--2609
		x"37",	--2610
		x"00",	--2611
		x"81",	--2612
		x"20",	--2613
		x"81",	--2614
		x"22",	--2615
		x"12",	--2616
		x"0f",	--2617
		x"0e",	--2618
		x"1a",	--2619
		x"0f",	--2620
		x"e7",	--2621
		x"81",	--2622
		x"0a",	--2623
		x"a6",	--2624
		x"6e",	--2625
		x"36",	--2626
		x"5f",	--2627
		x"d1",	--2628
		x"11",	--2629
		x"19",	--2630
		x"20",	--2631
		x"c1",	--2632
		x"19",	--2633
		x"0f",	--2634
		x"3f",	--2635
		x"18",	--2636
		x"c5",	--2637
		x"0d",	--2638
		x"ba",	--2639
		x"0c",	--2640
		x"0d",	--2641
		x"3c",	--2642
		x"80",	--2643
		x"0d",	--2644
		x"0c",	--2645
		x"b3",	--2646
		x"0d",	--2647
		x"b1",	--2648
		x"81",	--2649
		x"20",	--2650
		x"03",	--2651
		x"81",	--2652
		x"22",	--2653
		x"ab",	--2654
		x"3e",	--2655
		x"40",	--2656
		x"0f",	--2657
		x"3e",	--2658
		x"80",	--2659
		x"3f",	--2660
		x"a4",	--2661
		x"4d",	--2662
		x"7b",	--2663
		x"4f",	--2664
		x"de",	--2665
		x"5f",	--2666
		x"d1",	--2667
		x"11",	--2668
		x"19",	--2669
		x"06",	--2670
		x"c1",	--2671
		x"11",	--2672
		x"0f",	--2673
		x"3f",	--2674
		x"10",	--2675
		x"9e",	--2676
		x"4f",	--2677
		x"f8",	--2678
		x"6f",	--2679
		x"f1",	--2680
		x"3f",	--2681
		x"84",	--2682
		x"97",	--2683
		x"0b",	--2684
		x"0a",	--2685
		x"09",	--2686
		x"08",	--2687
		x"07",	--2688
		x"31",	--2689
		x"e8",	--2690
		x"81",	--2691
		x"04",	--2692
		x"81",	--2693
		x"06",	--2694
		x"81",	--2695
		x"00",	--2696
		x"81",	--2697
		x"02",	--2698
		x"0e",	--2699
		x"3e",	--2700
		x"10",	--2701
		x"0f",	--2702
		x"2f",	--2703
		x"b0",	--2704
		x"5a",	--2705
		x"0e",	--2706
		x"3e",	--2707
		x"0f",	--2708
		x"b0",	--2709
		x"5a",	--2710
		x"5f",	--2711
		x"10",	--2712
		x"6f",	--2713
		x"5d",	--2714
		x"5e",	--2715
		x"08",	--2716
		x"6e",	--2717
		x"82",	--2718
		x"d1",	--2719
		x"09",	--2720
		x"11",	--2721
		x"6f",	--2722
		x"58",	--2723
		x"6f",	--2724
		x"56",	--2725
		x"6e",	--2726
		x"6f",	--2727
		x"6e",	--2728
		x"4c",	--2729
		x"1d",	--2730
		x"12",	--2731
		x"1d",	--2732
		x"0a",	--2733
		x"81",	--2734
		x"12",	--2735
		x"1e",	--2736
		x"14",	--2737
		x"1f",	--2738
		x"16",	--2739
		x"18",	--2740
		x"0c",	--2741
		x"19",	--2742
		x"0e",	--2743
		x"0f",	--2744
		x"1e",	--2745
		x"0e",	--2746
		x"0f",	--2747
		x"3d",	--2748
		x"81",	--2749
		x"12",	--2750
		x"37",	--2751
		x"1f",	--2752
		x"0c",	--2753
		x"3d",	--2754
		x"00",	--2755
		x"0a",	--2756
		x"0b",	--2757
		x"0b",	--2758
		x"0a",	--2759
		x"0b",	--2760
		x"0e",	--2761
		x"0f",	--2762
		x"12",	--2763
		x"0d",	--2764
		x"0c",	--2765
		x"0e",	--2766
		x"0f",	--2767
		x"37",	--2768
		x"0b",	--2769
		x"0f",	--2770
		x"f7",	--2771
		x"f2",	--2772
		x"0e",	--2773
		x"f4",	--2774
		x"ef",	--2775
		x"09",	--2776
		x"e5",	--2777
		x"0e",	--2778
		x"e3",	--2779
		x"dd",	--2780
		x"0c",	--2781
		x"0d",	--2782
		x"3c",	--2783
		x"7f",	--2784
		x"0d",	--2785
		x"3c",	--2786
		x"40",	--2787
		x"1c",	--2788
		x"81",	--2789
		x"14",	--2790
		x"81",	--2791
		x"16",	--2792
		x"0f",	--2793
		x"3f",	--2794
		x"10",	--2795
		x"b0",	--2796
		x"7c",	--2797
		x"31",	--2798
		x"18",	--2799
		x"37",	--2800
		x"38",	--2801
		x"39",	--2802
		x"3a",	--2803
		x"3b",	--2804
		x"30",	--2805
		x"e1",	--2806
		x"10",	--2807
		x"0f",	--2808
		x"3f",	--2809
		x"10",	--2810
		x"f0",	--2811
		x"4f",	--2812
		x"fa",	--2813
		x"3f",	--2814
		x"84",	--2815
		x"eb",	--2816
		x"0d",	--2817
		x"e2",	--2818
		x"0c",	--2819
		x"0d",	--2820
		x"3c",	--2821
		x"80",	--2822
		x"0d",	--2823
		x"0c",	--2824
		x"db",	--2825
		x"0d",	--2826
		x"d9",	--2827
		x"0e",	--2828
		x"02",	--2829
		x"0f",	--2830
		x"d5",	--2831
		x"3a",	--2832
		x"40",	--2833
		x"0b",	--2834
		x"3a",	--2835
		x"80",	--2836
		x"3b",	--2837
		x"ce",	--2838
		x"81",	--2839
		x"14",	--2840
		x"81",	--2841
		x"16",	--2842
		x"81",	--2843
		x"12",	--2844
		x"0f",	--2845
		x"3f",	--2846
		x"10",	--2847
		x"cb",	--2848
		x"0f",	--2849
		x"3f",	--2850
		x"c8",	--2851
		x"31",	--2852
		x"e8",	--2853
		x"81",	--2854
		x"04",	--2855
		x"81",	--2856
		x"06",	--2857
		x"81",	--2858
		x"00",	--2859
		x"81",	--2860
		x"02",	--2861
		x"0e",	--2862
		x"3e",	--2863
		x"10",	--2864
		x"0f",	--2865
		x"2f",	--2866
		x"b0",	--2867
		x"5a",	--2868
		x"0e",	--2869
		x"3e",	--2870
		x"0f",	--2871
		x"b0",	--2872
		x"5a",	--2873
		x"e1",	--2874
		x"10",	--2875
		x"0d",	--2876
		x"e1",	--2877
		x"08",	--2878
		x"0a",	--2879
		x"0e",	--2880
		x"3e",	--2881
		x"0f",	--2882
		x"3f",	--2883
		x"10",	--2884
		x"b0",	--2885
		x"7e",	--2886
		x"31",	--2887
		x"18",	--2888
		x"30",	--2889
		x"3f",	--2890
		x"fb",	--2891
		x"31",	--2892
		x"f4",	--2893
		x"81",	--2894
		x"00",	--2895
		x"81",	--2896
		x"02",	--2897
		x"0e",	--2898
		x"2e",	--2899
		x"0f",	--2900
		x"b0",	--2901
		x"5a",	--2902
		x"5f",	--2903
		x"04",	--2904
		x"6f",	--2905
		x"28",	--2906
		x"27",	--2907
		x"6f",	--2908
		x"07",	--2909
		x"1d",	--2910
		x"06",	--2911
		x"0d",	--2912
		x"21",	--2913
		x"3d",	--2914
		x"1f",	--2915
		x"09",	--2916
		x"c1",	--2917
		x"05",	--2918
		x"26",	--2919
		x"3e",	--2920
		x"3f",	--2921
		x"ff",	--2922
		x"31",	--2923
		x"0c",	--2924
		x"30",	--2925
		x"1e",	--2926
		x"08",	--2927
		x"1f",	--2928
		x"0a",	--2929
		x"3c",	--2930
		x"1e",	--2931
		x"4c",	--2932
		x"4d",	--2933
		x"7d",	--2934
		x"1f",	--2935
		x"0f",	--2936
		x"c1",	--2937
		x"05",	--2938
		x"ef",	--2939
		x"3e",	--2940
		x"3f",	--2941
		x"1e",	--2942
		x"0f",	--2943
		x"31",	--2944
		x"0c",	--2945
		x"30",	--2946
		x"0e",	--2947
		x"0f",	--2948
		x"31",	--2949
		x"0c",	--2950
		x"30",	--2951
		x"12",	--2952
		x"0f",	--2953
		x"0e",	--2954
		x"7d",	--2955
		x"fb",	--2956
		x"eb",	--2957
		x"0e",	--2958
		x"3f",	--2959
		x"00",	--2960
		x"31",	--2961
		x"0c",	--2962
		x"30",	--2963
		x"0b",	--2964
		x"0a",	--2965
		x"09",	--2966
		x"08",	--2967
		x"31",	--2968
		x"0a",	--2969
		x"0b",	--2970
		x"c1",	--2971
		x"01",	--2972
		x"0e",	--2973
		x"0d",	--2974
		x"0b",	--2975
		x"0b",	--2976
		x"e1",	--2977
		x"00",	--2978
		x"0f",	--2979
		x"b0",	--2980
		x"7c",	--2981
		x"31",	--2982
		x"38",	--2983
		x"39",	--2984
		x"3a",	--2985
		x"3b",	--2986
		x"30",	--2987
		x"f1",	--2988
		x"03",	--2989
		x"00",	--2990
		x"b1",	--2991
		x"1e",	--2992
		x"02",	--2993
		x"81",	--2994
		x"04",	--2995
		x"81",	--2996
		x"06",	--2997
		x"0e",	--2998
		x"0f",	--2999
		x"b0",	--3000
		x"0a",	--3001
		x"3f",	--3002
		x"0f",	--3003
		x"18",	--3004
		x"e5",	--3005
		x"81",	--3006
		x"04",	--3007
		x"81",	--3008
		x"06",	--3009
		x"4e",	--3010
		x"7e",	--3011
		x"1f",	--3012
		x"06",	--3013
		x"3e",	--3014
		x"1e",	--3015
		x"0e",	--3016
		x"81",	--3017
		x"02",	--3018
		x"d7",	--3019
		x"91",	--3020
		x"04",	--3021
		x"04",	--3022
		x"91",	--3023
		x"06",	--3024
		x"06",	--3025
		x"7e",	--3026
		x"f8",	--3027
		x"f1",	--3028
		x"0e",	--3029
		x"3e",	--3030
		x"1e",	--3031
		x"1c",	--3032
		x"0d",	--3033
		x"48",	--3034
		x"78",	--3035
		x"1f",	--3036
		x"04",	--3037
		x"0c",	--3038
		x"0d",	--3039
		x"78",	--3040
		x"fc",	--3041
		x"3c",	--3042
		x"3d",	--3043
		x"0c",	--3044
		x"0d",	--3045
		x"18",	--3046
		x"09",	--3047
		x"0c",	--3048
		x"04",	--3049
		x"0d",	--3050
		x"02",	--3051
		x"08",	--3052
		x"09",	--3053
		x"7e",	--3054
		x"1f",	--3055
		x"0e",	--3056
		x"0d",	--3057
		x"0e",	--3058
		x"0d",	--3059
		x"0e",	--3060
		x"81",	--3061
		x"04",	--3062
		x"81",	--3063
		x"06",	--3064
		x"3e",	--3065
		x"1e",	--3066
		x"0e",	--3067
		x"81",	--3068
		x"02",	--3069
		x"a4",	--3070
		x"12",	--3071
		x"0b",	--3072
		x"0a",	--3073
		x"7e",	--3074
		x"fb",	--3075
		x"ec",	--3076
		x"0b",	--3077
		x"0a",	--3078
		x"09",	--3079
		x"1f",	--3080
		x"17",	--3081
		x"3e",	--3082
		x"00",	--3083
		x"2c",	--3084
		x"3a",	--3085
		x"18",	--3086
		x"0b",	--3087
		x"39",	--3088
		x"0c",	--3089
		x"0d",	--3090
		x"4f",	--3091
		x"4f",	--3092
		x"17",	--3093
		x"3c",	--3094
		x"8c",	--3095
		x"6e",	--3096
		x"0f",	--3097
		x"0a",	--3098
		x"0b",	--3099
		x"0f",	--3100
		x"39",	--3101
		x"3a",	--3102
		x"3b",	--3103
		x"30",	--3104
		x"3f",	--3105
		x"00",	--3106
		x"0f",	--3107
		x"3a",	--3108
		x"0b",	--3109
		x"39",	--3110
		x"18",	--3111
		x"0c",	--3112
		x"0d",	--3113
		x"4f",	--3114
		x"4f",	--3115
		x"e9",	--3116
		x"12",	--3117
		x"0d",	--3118
		x"0c",	--3119
		x"7f",	--3120
		x"fb",	--3121
		x"e3",	--3122
		x"3a",	--3123
		x"10",	--3124
		x"0b",	--3125
		x"39",	--3126
		x"10",	--3127
		x"ef",	--3128
		x"3a",	--3129
		x"20",	--3130
		x"0b",	--3131
		x"09",	--3132
		x"ea",	--3133
		x"0b",	--3134
		x"0a",	--3135
		x"09",	--3136
		x"08",	--3137
		x"07",	--3138
		x"0d",	--3139
		x"1e",	--3140
		x"04",	--3141
		x"1f",	--3142
		x"06",	--3143
		x"5a",	--3144
		x"01",	--3145
		x"6c",	--3146
		x"6c",	--3147
		x"70",	--3148
		x"6c",	--3149
		x"6a",	--3150
		x"6c",	--3151
		x"36",	--3152
		x"0e",	--3153
		x"32",	--3154
		x"1b",	--3155
		x"02",	--3156
		x"3b",	--3157
		x"82",	--3158
		x"6d",	--3159
		x"3b",	--3160
		x"80",	--3161
		x"5e",	--3162
		x"0c",	--3163
		x"0d",	--3164
		x"3c",	--3165
		x"7f",	--3166
		x"0d",	--3167
		x"3c",	--3168
		x"40",	--3169
		x"40",	--3170
		x"3e",	--3171
		x"3f",	--3172
		x"0f",	--3173
		x"0f",	--3174
		x"4a",	--3175
		x"0d",	--3176
		x"3d",	--3177
		x"7f",	--3178
		x"12",	--3179
		x"0f",	--3180
		x"0e",	--3181
		x"12",	--3182
		x"0f",	--3183
		x"0e",	--3184
		x"12",	--3185
		x"0f",	--3186
		x"0e",	--3187
		x"12",	--3188
		x"0f",	--3189
		x"0e",	--3190
		x"12",	--3191
		x"0f",	--3192
		x"0e",	--3193
		x"12",	--3194
		x"0f",	--3195
		x"0e",	--3196
		x"12",	--3197
		x"0f",	--3198
		x"0e",	--3199
		x"3e",	--3200
		x"3f",	--3201
		x"7f",	--3202
		x"4d",	--3203
		x"05",	--3204
		x"0f",	--3205
		x"cc",	--3206
		x"4d",	--3207
		x"0e",	--3208
		x"0f",	--3209
		x"4d",	--3210
		x"0d",	--3211
		x"0d",	--3212
		x"0d",	--3213
		x"0d",	--3214
		x"0d",	--3215
		x"0d",	--3216
		x"0d",	--3217
		x"0c",	--3218
		x"3c",	--3219
		x"7f",	--3220
		x"0c",	--3221
		x"4f",	--3222
		x"0f",	--3223
		x"0f",	--3224
		x"0f",	--3225
		x"0d",	--3226
		x"0d",	--3227
		x"0f",	--3228
		x"37",	--3229
		x"38",	--3230
		x"39",	--3231
		x"3a",	--3232
		x"3b",	--3233
		x"30",	--3234
		x"0d",	--3235
		x"be",	--3236
		x"0c",	--3237
		x"0d",	--3238
		x"3c",	--3239
		x"80",	--3240
		x"0d",	--3241
		x"0c",	--3242
		x"02",	--3243
		x"0d",	--3244
		x"b8",	--3245
		x"3e",	--3246
		x"40",	--3247
		x"0f",	--3248
		x"b4",	--3249
		x"12",	--3250
		x"0f",	--3251
		x"0e",	--3252
		x"0d",	--3253
		x"3d",	--3254
		x"80",	--3255
		x"b2",	--3256
		x"7d",	--3257
		x"0e",	--3258
		x"0f",	--3259
		x"cd",	--3260
		x"0e",	--3261
		x"3f",	--3262
		x"10",	--3263
		x"3e",	--3264
		x"3f",	--3265
		x"7f",	--3266
		x"7d",	--3267
		x"c5",	--3268
		x"37",	--3269
		x"82",	--3270
		x"07",	--3271
		x"37",	--3272
		x"1a",	--3273
		x"4f",	--3274
		x"0c",	--3275
		x"0d",	--3276
		x"4b",	--3277
		x"7b",	--3278
		x"1f",	--3279
		x"05",	--3280
		x"12",	--3281
		x"0d",	--3282
		x"0c",	--3283
		x"7b",	--3284
		x"fb",	--3285
		x"18",	--3286
		x"09",	--3287
		x"77",	--3288
		x"1f",	--3289
		x"04",	--3290
		x"08",	--3291
		x"09",	--3292
		x"77",	--3293
		x"fc",	--3294
		x"38",	--3295
		x"39",	--3296
		x"08",	--3297
		x"09",	--3298
		x"1e",	--3299
		x"0f",	--3300
		x"08",	--3301
		x"04",	--3302
		x"09",	--3303
		x"02",	--3304
		x"0e",	--3305
		x"0f",	--3306
		x"08",	--3307
		x"09",	--3308
		x"08",	--3309
		x"09",	--3310
		x"0e",	--3311
		x"0f",	--3312
		x"3e",	--3313
		x"7f",	--3314
		x"0f",	--3315
		x"3e",	--3316
		x"40",	--3317
		x"26",	--3318
		x"38",	--3319
		x"3f",	--3320
		x"09",	--3321
		x"0e",	--3322
		x"0f",	--3323
		x"12",	--3324
		x"0f",	--3325
		x"0e",	--3326
		x"12",	--3327
		x"0f",	--3328
		x"0e",	--3329
		x"12",	--3330
		x"0f",	--3331
		x"0e",	--3332
		x"12",	--3333
		x"0f",	--3334
		x"0e",	--3335
		x"12",	--3336
		x"0f",	--3337
		x"0e",	--3338
		x"12",	--3339
		x"0f",	--3340
		x"0e",	--3341
		x"12",	--3342
		x"0f",	--3343
		x"0e",	--3344
		x"3e",	--3345
		x"3f",	--3346
		x"7f",	--3347
		x"5d",	--3348
		x"39",	--3349
		x"00",	--3350
		x"72",	--3351
		x"4d",	--3352
		x"70",	--3353
		x"08",	--3354
		x"09",	--3355
		x"da",	--3356
		x"0f",	--3357
		x"d8",	--3358
		x"0e",	--3359
		x"0f",	--3360
		x"3e",	--3361
		x"80",	--3362
		x"0f",	--3363
		x"0e",	--3364
		x"04",	--3365
		x"38",	--3366
		x"40",	--3367
		x"09",	--3368
		x"d0",	--3369
		x"0f",	--3370
		x"ce",	--3371
		x"f9",	--3372
		x"0b",	--3373
		x"0a",	--3374
		x"2a",	--3375
		x"5b",	--3376
		x"02",	--3377
		x"3b",	--3378
		x"7f",	--3379
		x"1d",	--3380
		x"02",	--3381
		x"12",	--3382
		x"0d",	--3383
		x"12",	--3384
		x"0d",	--3385
		x"12",	--3386
		x"0d",	--3387
		x"12",	--3388
		x"0d",	--3389
		x"12",	--3390
		x"0d",	--3391
		x"12",	--3392
		x"0d",	--3393
		x"12",	--3394
		x"0d",	--3395
		x"4d",	--3396
		x"5f",	--3397
		x"03",	--3398
		x"3f",	--3399
		x"80",	--3400
		x"0f",	--3401
		x"0f",	--3402
		x"ce",	--3403
		x"01",	--3404
		x"0d",	--3405
		x"2d",	--3406
		x"0a",	--3407
		x"51",	--3408
		x"be",	--3409
		x"82",	--3410
		x"02",	--3411
		x"0c",	--3412
		x"0d",	--3413
		x"0c",	--3414
		x"0d",	--3415
		x"0c",	--3416
		x"0d",	--3417
		x"0c",	--3418
		x"0d",	--3419
		x"0c",	--3420
		x"0d",	--3421
		x"0c",	--3422
		x"0d",	--3423
		x"0c",	--3424
		x"0d",	--3425
		x"0c",	--3426
		x"0d",	--3427
		x"fe",	--3428
		x"03",	--3429
		x"00",	--3430
		x"3d",	--3431
		x"00",	--3432
		x"0b",	--3433
		x"3f",	--3434
		x"81",	--3435
		x"0c",	--3436
		x"0d",	--3437
		x"0a",	--3438
		x"3f",	--3439
		x"3d",	--3440
		x"00",	--3441
		x"f9",	--3442
		x"8e",	--3443
		x"02",	--3444
		x"8e",	--3445
		x"04",	--3446
		x"8e",	--3447
		x"06",	--3448
		x"3a",	--3449
		x"3b",	--3450
		x"30",	--3451
		x"3d",	--3452
		x"ff",	--3453
		x"2a",	--3454
		x"3d",	--3455
		x"81",	--3456
		x"8e",	--3457
		x"02",	--3458
		x"fe",	--3459
		x"03",	--3460
		x"00",	--3461
		x"0c",	--3462
		x"0d",	--3463
		x"0c",	--3464
		x"0d",	--3465
		x"0c",	--3466
		x"0d",	--3467
		x"0c",	--3468
		x"0d",	--3469
		x"0c",	--3470
		x"0d",	--3471
		x"0c",	--3472
		x"0d",	--3473
		x"0c",	--3474
		x"0d",	--3475
		x"0c",	--3476
		x"0d",	--3477
		x"0a",	--3478
		x"0b",	--3479
		x"0a",	--3480
		x"3b",	--3481
		x"00",	--3482
		x"8e",	--3483
		x"04",	--3484
		x"8e",	--3485
		x"06",	--3486
		x"3a",	--3487
		x"3b",	--3488
		x"30",	--3489
		x"0b",	--3490
		x"ad",	--3491
		x"ee",	--3492
		x"00",	--3493
		x"3a",	--3494
		x"3b",	--3495
		x"30",	--3496
		x"0a",	--3497
		x"0c",	--3498
		x"0c",	--3499
		x"0d",	--3500
		x"0c",	--3501
		x"3d",	--3502
		x"10",	--3503
		x"0c",	--3504
		x"02",	--3505
		x"0d",	--3506
		x"08",	--3507
		x"de",	--3508
		x"00",	--3509
		x"e4",	--3510
		x"0b",	--3511
		x"f2",	--3512
		x"ee",	--3513
		x"00",	--3514
		x"e3",	--3515
		x"ce",	--3516
		x"00",	--3517
		x"dc",	--3518
		x"0b",	--3519
		x"6d",	--3520
		x"6d",	--3521
		x"12",	--3522
		x"6c",	--3523
		x"6c",	--3524
		x"0f",	--3525
		x"6d",	--3526
		x"41",	--3527
		x"6c",	--3528
		x"11",	--3529
		x"6d",	--3530
		x"0d",	--3531
		x"6c",	--3532
		x"14",	--3533
		x"5d",	--3534
		x"01",	--3535
		x"5d",	--3536
		x"01",	--3537
		x"14",	--3538
		x"4d",	--3539
		x"09",	--3540
		x"1e",	--3541
		x"0f",	--3542
		x"3b",	--3543
		x"30",	--3544
		x"6c",	--3545
		x"28",	--3546
		x"ce",	--3547
		x"01",	--3548
		x"f7",	--3549
		x"3e",	--3550
		x"0f",	--3551
		x"3b",	--3552
		x"30",	--3553
		x"cf",	--3554
		x"01",	--3555
		x"f0",	--3556
		x"3e",	--3557
		x"f8",	--3558
		x"1b",	--3559
		x"02",	--3560
		x"1c",	--3561
		x"02",	--3562
		x"0c",	--3563
		x"e6",	--3564
		x"0b",	--3565
		x"16",	--3566
		x"1b",	--3567
		x"04",	--3568
		x"1f",	--3569
		x"06",	--3570
		x"1c",	--3571
		x"04",	--3572
		x"1e",	--3573
		x"06",	--3574
		x"0e",	--3575
		x"da",	--3576
		x"0f",	--3577
		x"02",	--3578
		x"0c",	--3579
		x"d6",	--3580
		x"0f",	--3581
		x"06",	--3582
		x"0e",	--3583
		x"02",	--3584
		x"0b",	--3585
		x"02",	--3586
		x"0e",	--3587
		x"d1",	--3588
		x"4d",	--3589
		x"ce",	--3590
		x"3e",	--3591
		x"d6",	--3592
		x"6c",	--3593
		x"d7",	--3594
		x"5e",	--3595
		x"01",	--3596
		x"5f",	--3597
		x"01",	--3598
		x"0e",	--3599
		x"c5",	--3600
		x"1e",	--3601
		x"1c",	--3602
		x"1e",	--3603
		x"0b",	--3604
		x"1d",	--3605
		x"1a",	--3606
		x"cd",	--3607
		x"00",	--3608
		x"1d",	--3609
		x"82",	--3610
		x"1a",	--3611
		x"3e",	--3612
		x"82",	--3613
		x"1c",	--3614
		x"30",	--3615
		x"3f",	--3616
		x"30",	--3617
		x"0b",	--3618
		x"0a",	--3619
		x"21",	--3620
		x"81",	--3621
		x"00",	--3622
		x"1a",	--3623
		x"1a",	--3624
		x"1b",	--3625
		x"1c",	--3626
		x"0d",	--3627
		x"0e",	--3628
		x"3f",	--3629
		x"22",	--3630
		x"b0",	--3631
		x"76",	--3632
		x"0f",	--3633
		x"05",	--3634
		x"0e",	--3635
		x"0e",	--3636
		x"ce",	--3637
		x"ff",	--3638
		x"04",	--3639
		x"1e",	--3640
		x"1a",	--3641
		x"ce",	--3642
		x"00",	--3643
		x"21",	--3644
		x"3a",	--3645
		x"3b",	--3646
		x"30",	--3647
		x"92",	--3648
		x"02",	--3649
		x"1a",	--3650
		x"b2",	--3651
		x"ff",	--3652
		x"1c",	--3653
		x"0e",	--3654
		x"3e",	--3655
		x"06",	--3656
		x"1f",	--3657
		x"04",	--3658
		x"b0",	--3659
		x"44",	--3660
		x"30",	--3661
		x"92",	--3662
		x"02",	--3663
		x"1a",	--3664
		x"92",	--3665
		x"04",	--3666
		x"1c",	--3667
		x"0e",	--3668
		x"3e",	--3669
		x"1f",	--3670
		x"06",	--3671
		x"b0",	--3672
		x"44",	--3673
		x"30",	--3674
		x"0c",	--3675
		x"82",	--3676
		x"1a",	--3677
		x"b2",	--3678
		x"ff",	--3679
		x"1c",	--3680
		x"0e",	--3681
		x"0f",	--3682
		x"b0",	--3683
		x"44",	--3684
		x"30",	--3685
		x"82",	--3686
		x"1a",	--3687
		x"82",	--3688
		x"1c",	--3689
		x"0e",	--3690
		x"0f",	--3691
		x"b0",	--3692
		x"44",	--3693
		x"30",	--3694
		x"0b",	--3695
		x"0a",	--3696
		x"09",	--3697
		x"08",	--3698
		x"07",	--3699
		x"06",	--3700
		x"05",	--3701
		x"04",	--3702
		x"31",	--3703
		x"08",	--3704
		x"81",	--3705
		x"04",	--3706
		x"09",	--3707
		x"1f",	--3708
		x"1a",	--3709
		x"1d",	--3710
		x"1c",	--3711
		x"4c",	--3712
		x"04",	--3713
		x"84",	--3714
		x"45",	--3715
		x"4e",	--3716
		x"7e",	--3717
		x"40",	--3718
		x"11",	--3719
		x"f1",	--3720
		x"30",	--3721
		x"00",	--3722
		x"0e",	--3723
		x"8e",	--3724
		x"5e",	--3725
		x"03",	--3726
		x"7e",	--3727
		x"58",	--3728
		x"02",	--3729
		x"7e",	--3730
		x"78",	--3731
		x"c1",	--3732
		x"01",	--3733
		x"0c",	--3734
		x"2c",	--3735
		x"0f",	--3736
		x"7e",	--3737
		x"20",	--3738
		x"04",	--3739
		x"f1",	--3740
		x"30",	--3741
		x"00",	--3742
		x"04",	--3743
		x"4c",	--3744
		x"05",	--3745
		x"c1",	--3746
		x"00",	--3747
		x"0c",	--3748
		x"1c",	--3749
		x"01",	--3750
		x"0c",	--3751
		x"0a",	--3752
		x"8c",	--3753
		x"8c",	--3754
		x"8c",	--3755
		x"8c",	--3756
		x"0b",	--3757
		x"06",	--3758
		x"0c",	--3759
		x"8c",	--3760
		x"8c",	--3761
		x"8c",	--3762
		x"8c",	--3763
		x"07",	--3764
		x"0a",	--3765
		x"0b",	--3766
		x"0e",	--3767
		x"8e",	--3768
		x"c1",	--3769
		x"02",	--3770
		x"6e",	--3771
		x"02",	--3772
		x"07",	--3773
		x"01",	--3774
		x"37",	--3775
		x"4f",	--3776
		x"7f",	--3777
		x"10",	--3778
		x"3c",	--3779
		x"1d",	--3780
		x"04",	--3781
		x"3d",	--3782
		x"1d",	--3783
		x"cd",	--3784
		x"00",	--3785
		x"fc",	--3786
		x"1d",	--3787
		x"04",	--3788
		x"09",	--3789
		x"02",	--3790
		x"09",	--3791
		x"01",	--3792
		x"09",	--3793
		x"e1",	--3794
		x"02",	--3795
		x"05",	--3796
		x"09",	--3797
		x"02",	--3798
		x"09",	--3799
		x"01",	--3800
		x"09",	--3801
		x"05",	--3802
		x"07",	--3803
		x"01",	--3804
		x"05",	--3805
		x"4f",	--3806
		x"0d",	--3807
		x"f1",	--3808
		x"20",	--3809
		x"06",	--3810
		x"06",	--3811
		x"0b",	--3812
		x"0e",	--3813
		x"0f",	--3814
		x"0f",	--3815
		x"6f",	--3816
		x"8f",	--3817
		x"16",	--3818
		x"88",	--3819
		x"01",	--3820
		x"06",	--3821
		x"06",	--3822
		x"f6",	--3823
		x"0b",	--3824
		x"f1",	--3825
		x"30",	--3826
		x"06",	--3827
		x"05",	--3828
		x"05",	--3829
		x"5f",	--3830
		x"06",	--3831
		x"8f",	--3832
		x"88",	--3833
		x"1b",	--3834
		x"0f",	--3835
		x"0f",	--3836
		x"0f",	--3837
		x"f7",	--3838
		x"0a",	--3839
		x"06",	--3840
		x"0b",	--3841
		x"07",	--3842
		x"1b",	--3843
		x"0f",	--3844
		x"0f",	--3845
		x"6f",	--3846
		x"8f",	--3847
		x"16",	--3848
		x"88",	--3849
		x"06",	--3850
		x"f7",	--3851
		x"e1",	--3852
		x"02",	--3853
		x"02",	--3854
		x"4a",	--3855
		x"08",	--3856
		x"1a",	--3857
		x"04",	--3858
		x"0a",	--3859
		x"0d",	--3860
		x"3f",	--3861
		x"30",	--3862
		x"88",	--3863
		x"7a",	--3864
		x"4a",	--3865
		x"fa",	--3866
		x"44",	--3867
		x"0b",	--3868
		x"f3",	--3869
		x"37",	--3870
		x"8f",	--3871
		x"88",	--3872
		x"1b",	--3873
		x"0f",	--3874
		x"0f",	--3875
		x"6f",	--3876
		x"4f",	--3877
		x"07",	--3878
		x"07",	--3879
		x"f5",	--3880
		x"04",	--3881
		x"3f",	--3882
		x"20",	--3883
		x"88",	--3884
		x"1b",	--3885
		x"0b",	--3886
		x"fa",	--3887
		x"0f",	--3888
		x"31",	--3889
		x"34",	--3890
		x"35",	--3891
		x"36",	--3892
		x"37",	--3893
		x"38",	--3894
		x"39",	--3895
		x"3a",	--3896
		x"3b",	--3897
		x"30",	--3898
		x"0b",	--3899
		x"0a",	--3900
		x"09",	--3901
		x"08",	--3902
		x"07",	--3903
		x"06",	--3904
		x"05",	--3905
		x"04",	--3906
		x"31",	--3907
		x"b6",	--3908
		x"81",	--3909
		x"3a",	--3910
		x"06",	--3911
		x"05",	--3912
		x"81",	--3913
		x"3e",	--3914
		x"c1",	--3915
		x"2f",	--3916
		x"c1",	--3917
		x"2b",	--3918
		x"c1",	--3919
		x"2e",	--3920
		x"c1",	--3921
		x"2a",	--3922
		x"81",	--3923
		x"30",	--3924
		x"81",	--3925
		x"26",	--3926
		x"07",	--3927
		x"81",	--3928
		x"2c",	--3929
		x"0e",	--3930
		x"3e",	--3931
		x"1c",	--3932
		x"81",	--3933
		x"1c",	--3934
		x"30",	--3935
		x"f0",	--3936
		x"0f",	--3937
		x"1f",	--3938
		x"81",	--3939
		x"40",	--3940
		x"07",	--3941
		x"1e",	--3942
		x"7e",	--3943
		x"25",	--3944
		x"13",	--3945
		x"81",	--3946
		x"00",	--3947
		x"81",	--3948
		x"02",	--3949
		x"81",	--3950
		x"3e",	--3951
		x"c1",	--3952
		x"2f",	--3953
		x"c1",	--3954
		x"2b",	--3955
		x"c1",	--3956
		x"2e",	--3957
		x"c1",	--3958
		x"2a",	--3959
		x"81",	--3960
		x"30",	--3961
		x"30",	--3962
		x"e6",	--3963
		x"05",	--3964
		x"8e",	--3965
		x"0f",	--3966
		x"91",	--3967
		x"3c",	--3968
		x"91",	--3969
		x"2c",	--3970
		x"30",	--3971
		x"cc",	--3972
		x"7e",	--3973
		x"63",	--3974
		x"c5",	--3975
		x"7e",	--3976
		x"64",	--3977
		x"27",	--3978
		x"7e",	--3979
		x"30",	--3980
		x"94",	--3981
		x"7e",	--3982
		x"31",	--3983
		x"1a",	--3984
		x"7e",	--3985
		x"2a",	--3986
		x"77",	--3987
		x"7e",	--3988
		x"2b",	--3989
		x"0a",	--3990
		x"7e",	--3991
		x"23",	--3992
		x"42",	--3993
		x"7e",	--3994
		x"25",	--3995
		x"e0",	--3996
		x"7e",	--3997
		x"20",	--3998
		x"32",	--3999
		x"56",	--4000
		x"7e",	--4001
		x"2d",	--4002
		x"49",	--4003
		x"7e",	--4004
		x"2e",	--4005
		x"5b",	--4006
		x"7e",	--4007
		x"2b",	--4008
		x"28",	--4009
		x"47",	--4010
		x"7e",	--4011
		x"3a",	--4012
		x"8c",	--4013
		x"7e",	--4014
		x"58",	--4015
		x"21",	--4016
		x"e9",	--4017
		x"7e",	--4018
		x"6f",	--4019
		x"24",	--4020
		x"7e",	--4021
		x"70",	--4022
		x"0a",	--4023
		x"7e",	--4024
		x"69",	--4025
		x"e3",	--4026
		x"7e",	--4027
		x"6c",	--4028
		x"22",	--4029
		x"7e",	--4030
		x"64",	--4031
		x"11",	--4032
		x"dc",	--4033
		x"7e",	--4034
		x"73",	--4035
		x"98",	--4036
		x"7e",	--4037
		x"74",	--4038
		x"04",	--4039
		x"7e",	--4040
		x"70",	--4041
		x"07",	--4042
		x"b8",	--4043
		x"7e",	--4044
		x"75",	--4045
		x"d1",	--4046
		x"7e",	--4047
		x"78",	--4048
		x"d2",	--4049
		x"19",	--4050
		x"3e",	--4051
		x"18",	--4052
		x"2c",	--4053
		x"08",	--4054
		x"30",	--4055
		x"ba",	--4056
		x"b1",	--4057
		x"28",	--4058
		x"cb",	--4059
		x"f1",	--4060
		x"00",	--4061
		x"30",	--4062
		x"ea",	--4063
		x"69",	--4064
		x"59",	--4065
		x"6e",	--4066
		x"04",	--4067
		x"7e",	--4068
		x"fe",	--4069
		x"6e",	--4070
		x"01",	--4071
		x"5e",	--4072
		x"c1",	--4073
		x"00",	--4074
		x"30",	--4075
		x"ea",	--4076
		x"f1",	--4077
		x"10",	--4078
		x"00",	--4079
		x"30",	--4080
		x"ea",	--4081
		x"f1",	--4082
		x"2b",	--4083
		x"02",	--4084
		x"30",	--4085
		x"ea",	--4086
		x"f1",	--4087
		x"2b",	--4088
		x"02",	--4089
		x"02",	--4090
		x"30",	--4091
		x"ea",	--4092
		x"f1",	--4093
		x"20",	--4094
		x"02",	--4095
		x"30",	--4096
		x"ea",	--4097
		x"c1",	--4098
		x"2a",	--4099
		x"02",	--4100
		x"30",	--4101
		x"d0",	--4102
		x"d1",	--4103
		x"2e",	--4104
		x"30",	--4105
		x"ea",	--4106
		x"0e",	--4107
		x"2e",	--4108
		x"2a",	--4109
		x"0a",	--4110
		x"03",	--4111
		x"81",	--4112
		x"26",	--4113
		x"0d",	--4114
		x"c1",	--4115
		x"2e",	--4116
		x"02",	--4117
		x"30",	--4118
		x"e0",	--4119
		x"f1",	--4120
		x"10",	--4121
		x"00",	--4122
		x"3a",	--4123
		x"81",	--4124
		x"26",	--4125
		x"91",	--4126
		x"26",	--4127
		x"05",	--4128
		x"27",	--4129
		x"81",	--4130
		x"26",	--4131
		x"15",	--4132
		x"c1",	--4133
		x"2e",	--4134
		x"12",	--4135
		x"69",	--4136
		x"79",	--4137
		x"10",	--4138
		x"5e",	--4139
		x"01",	--4140
		x"4e",	--4141
		x"4e",	--4142
		x"0e",	--4143
		x"0e",	--4144
		x"4e",	--4145
		x"6a",	--4146
		x"7a",	--4147
		x"7f",	--4148
		x"4a",	--4149
		x"c1",	--4150
		x"00",	--4151
		x"30",	--4152
		x"ea",	--4153
		x"1a",	--4154
		x"26",	--4155
		x"0a",	--4156
		x"0c",	--4157
		x"0c",	--4158
		x"0c",	--4159
		x"0a",	--4160
		x"81",	--4161
		x"26",	--4162
		x"b1",	--4163
		x"d0",	--4164
		x"26",	--4165
		x"8e",	--4166
		x"81",	--4167
		x"26",	--4168
		x"d1",	--4169
		x"2a",	--4170
		x"30",	--4171
		x"ea",	--4172
		x"07",	--4173
		x"27",	--4174
		x"6e",	--4175
		x"c1",	--4176
		x"2e",	--4177
		x"03",	--4178
		x"c1",	--4179
		x"2a",	--4180
		x"26",	--4181
		x"c1",	--4182
		x"04",	--4183
		x"c1",	--4184
		x"05",	--4185
		x"0e",	--4186
		x"2e",	--4187
		x"03",	--4188
		x"07",	--4189
		x"27",	--4190
		x"2e",	--4191
		x"c1",	--4192
		x"2e",	--4193
		x"07",	--4194
		x"e1",	--4195
		x"01",	--4196
		x"1f",	--4197
		x"26",	--4198
		x"c1",	--4199
		x"03",	--4200
		x"06",	--4201
		x"c1",	--4202
		x"2a",	--4203
		x"03",	--4204
		x"91",	--4205
		x"26",	--4206
		x"30",	--4207
		x"0e",	--4208
		x"02",	--4209
		x"3e",	--4210
		x"8c",	--4211
		x"11",	--4212
		x"04",	--4213
		x"11",	--4214
		x"04",	--4215
		x"1d",	--4216
		x"34",	--4217
		x"1f",	--4218
		x"3e",	--4219
		x"b0",	--4220
		x"de",	--4221
		x"21",	--4222
		x"81",	--4223
		x"2c",	--4224
		x"05",	--4225
		x"30",	--4226
		x"cc",	--4227
		x"07",	--4228
		x"27",	--4229
		x"29",	--4230
		x"81",	--4231
		x"1e",	--4232
		x"5e",	--4233
		x"09",	--4234
		x"01",	--4235
		x"4e",	--4236
		x"4e",	--4237
		x"4e",	--4238
		x"4e",	--4239
		x"6a",	--4240
		x"7a",	--4241
		x"f7",	--4242
		x"4a",	--4243
		x"c1",	--4244
		x"00",	--4245
		x"05",	--4246
		x"b1",	--4247
		x"10",	--4248
		x"28",	--4249
		x"53",	--4250
		x"d1",	--4251
		x"01",	--4252
		x"06",	--4253
		x"e1",	--4254
		x"00",	--4255
		x"b1",	--4256
		x"0a",	--4257
		x"28",	--4258
		x"03",	--4259
		x"b1",	--4260
		x"10",	--4261
		x"28",	--4262
		x"6b",	--4263
		x"6b",	--4264
		x"24",	--4265
		x"0c",	--4266
		x"3c",	--4267
		x"28",	--4268
		x"17",	--4269
		x"02",	--4270
		x"16",	--4271
		x"04",	--4272
		x"1b",	--4273
		x"06",	--4274
		x"81",	--4275
		x"1e",	--4276
		x"81",	--4277
		x"20",	--4278
		x"81",	--4279
		x"22",	--4280
		x"81",	--4281
		x"24",	--4282
		x"d1",	--4283
		x"2b",	--4284
		x"08",	--4285
		x"06",	--4286
		x"07",	--4287
		x"04",	--4288
		x"06",	--4289
		x"02",	--4290
		x"0b",	--4291
		x"02",	--4292
		x"c1",	--4293
		x"2b",	--4294
		x"0b",	--4295
		x"0b",	--4296
		x"0b",	--4297
		x"c1",	--4298
		x"2f",	--4299
		x"05",	--4300
		x"20",	--4301
		x"5b",	--4302
		x"07",	--4303
		x"0d",	--4304
		x"27",	--4305
		x"28",	--4306
		x"1b",	--4307
		x"02",	--4308
		x"81",	--4309
		x"1e",	--4310
		x"81",	--4311
		x"20",	--4312
		x"d1",	--4313
		x"2b",	--4314
		x"08",	--4315
		x"09",	--4316
		x"06",	--4317
		x"27",	--4318
		x"2b",	--4319
		x"81",	--4320
		x"1e",	--4321
		x"d1",	--4322
		x"2b",	--4323
		x"0b",	--4324
		x"02",	--4325
		x"c1",	--4326
		x"2b",	--4327
		x"0b",	--4328
		x"0b",	--4329
		x"0b",	--4330
		x"c1",	--4331
		x"2f",	--4332
		x"05",	--4333
		x"f1",	--4334
		x"00",	--4335
		x"12",	--4336
		x"c1",	--4337
		x"2b",	--4338
		x"0f",	--4339
		x"68",	--4340
		x"b1",	--4341
		x"10",	--4342
		x"28",	--4343
		x"03",	--4344
		x"78",	--4345
		x"40",	--4346
		x"05",	--4347
		x"b1",	--4348
		x"28",	--4349
		x"04",	--4350
		x"78",	--4351
		x"20",	--4352
		x"c1",	--4353
		x"00",	--4354
		x"68",	--4355
		x"68",	--4356
		x"30",	--4357
		x"c1",	--4358
		x"2f",	--4359
		x"2d",	--4360
		x"f1",	--4361
		x"2d",	--4362
		x"02",	--4363
		x"68",	--4364
		x"11",	--4365
		x"b1",	--4366
		x"1e",	--4367
		x"b1",	--4368
		x"20",	--4369
		x"b1",	--4370
		x"22",	--4371
		x"b1",	--4372
		x"24",	--4373
		x"91",	--4374
		x"1e",	--4375
		x"81",	--4376
		x"20",	--4377
		x"81",	--4378
		x"22",	--4379
		x"81",	--4380
		x"24",	--4381
		x"17",	--4382
		x"58",	--4383
		x"0f",	--4384
		x"1a",	--4385
		x"1e",	--4386
		x"1b",	--4387
		x"20",	--4388
		x"3a",	--4389
		x"3b",	--4390
		x"0e",	--4391
		x"0f",	--4392
		x"1e",	--4393
		x"0f",	--4394
		x"81",	--4395
		x"1e",	--4396
		x"81",	--4397
		x"20",	--4398
		x"06",	--4399
		x"1a",	--4400
		x"1e",	--4401
		x"3a",	--4402
		x"1a",	--4403
		x"81",	--4404
		x"1e",	--4405
		x"c1",	--4406
		x"1b",	--4407
		x"68",	--4408
		x"6a",	--4409
		x"16",	--4410
		x"1e",	--4411
		x"91",	--4412
		x"20",	--4413
		x"3c",	--4414
		x"18",	--4415
		x"22",	--4416
		x"14",	--4417
		x"24",	--4418
		x"07",	--4419
		x"37",	--4420
		x"1a",	--4421
		x"09",	--4422
		x"91",	--4423
		x"28",	--4424
		x"32",	--4425
		x"1b",	--4426
		x"28",	--4427
		x"8b",	--4428
		x"8b",	--4429
		x"8b",	--4430
		x"8b",	--4431
		x"81",	--4432
		x"34",	--4433
		x"81",	--4434
		x"36",	--4435
		x"81",	--4436
		x"38",	--4437
		x"11",	--4438
		x"3a",	--4439
		x"11",	--4440
		x"3a",	--4441
		x"11",	--4442
		x"3a",	--4443
		x"11",	--4444
		x"3a",	--4445
		x"0c",	--4446
		x"1d",	--4447
		x"44",	--4448
		x"0e",	--4449
		x"0f",	--4450
		x"b0",	--4451
		x"80",	--4452
		x"31",	--4453
		x"0b",	--4454
		x"3c",	--4455
		x"0a",	--4456
		x"05",	--4457
		x"7b",	--4458
		x"30",	--4459
		x"c7",	--4460
		x"00",	--4461
		x"0c",	--4462
		x"4b",	--4463
		x"d1",	--4464
		x"01",	--4465
		x"03",	--4466
		x"7a",	--4467
		x"37",	--4468
		x"02",	--4469
		x"7a",	--4470
		x"57",	--4471
		x"4a",	--4472
		x"c7",	--4473
		x"00",	--4474
		x"06",	--4475
		x"36",	--4476
		x"11",	--4477
		x"3a",	--4478
		x"11",	--4479
		x"3a",	--4480
		x"11",	--4481
		x"3a",	--4482
		x"11",	--4483
		x"3a",	--4484
		x"0c",	--4485
		x"1d",	--4486
		x"44",	--4487
		x"0e",	--4488
		x"0f",	--4489
		x"b0",	--4490
		x"5a",	--4491
		x"31",	--4492
		x"09",	--4493
		x"81",	--4494
		x"3c",	--4495
		x"08",	--4496
		x"04",	--4497
		x"37",	--4498
		x"0c",	--4499
		x"b2",	--4500
		x"0d",	--4501
		x"b0",	--4502
		x"0e",	--4503
		x"ae",	--4504
		x"0f",	--4505
		x"ac",	--4506
		x"81",	--4507
		x"1e",	--4508
		x"81",	--4509
		x"20",	--4510
		x"81",	--4511
		x"22",	--4512
		x"81",	--4513
		x"24",	--4514
		x"6c",	--4515
		x"58",	--4516
		x"3e",	--4517
		x"14",	--4518
		x"1e",	--4519
		x"17",	--4520
		x"20",	--4521
		x"08",	--4522
		x"38",	--4523
		x"1a",	--4524
		x"19",	--4525
		x"28",	--4526
		x"89",	--4527
		x"89",	--4528
		x"89",	--4529
		x"89",	--4530
		x"1c",	--4531
		x"28",	--4532
		x"0d",	--4533
		x"0e",	--4534
		x"0f",	--4535
		x"b0",	--4536
		x"84",	--4537
		x"0b",	--4538
		x"3e",	--4539
		x"0a",	--4540
		x"05",	--4541
		x"7b",	--4542
		x"30",	--4543
		x"c8",	--4544
		x"00",	--4545
		x"0c",	--4546
		x"4b",	--4547
		x"d1",	--4548
		x"01",	--4549
		x"03",	--4550
		x"7a",	--4551
		x"37",	--4552
		x"02",	--4553
		x"7a",	--4554
		x"57",	--4555
		x"4a",	--4556
		x"c8",	--4557
		x"00",	--4558
		x"06",	--4559
		x"36",	--4560
		x"1c",	--4561
		x"28",	--4562
		x"0d",	--4563
		x"0e",	--4564
		x"0f",	--4565
		x"b0",	--4566
		x"4e",	--4567
		x"04",	--4568
		x"07",	--4569
		x"38",	--4570
		x"0e",	--4571
		x"d0",	--4572
		x"0f",	--4573
		x"ce",	--4574
		x"81",	--4575
		x"1e",	--4576
		x"81",	--4577
		x"20",	--4578
		x"2c",	--4579
		x"17",	--4580
		x"1e",	--4581
		x"08",	--4582
		x"38",	--4583
		x"1a",	--4584
		x"1e",	--4585
		x"28",	--4586
		x"0f",	--4587
		x"b0",	--4588
		x"f4",	--4589
		x"0d",	--4590
		x"3f",	--4591
		x"0a",	--4592
		x"05",	--4593
		x"7d",	--4594
		x"30",	--4595
		x"c8",	--4596
		x"00",	--4597
		x"0c",	--4598
		x"4d",	--4599
		x"d1",	--4600
		x"01",	--4601
		x"03",	--4602
		x"7c",	--4603
		x"37",	--4604
		x"02",	--4605
		x"7c",	--4606
		x"57",	--4607
		x"4c",	--4608
		x"c8",	--4609
		x"00",	--4610
		x"06",	--4611
		x"36",	--4612
		x"1e",	--4613
		x"28",	--4614
		x"0f",	--4615
		x"b0",	--4616
		x"da",	--4617
		x"07",	--4618
		x"38",	--4619
		x"0f",	--4620
		x"db",	--4621
		x"81",	--4622
		x"1e",	--4623
		x"b1",	--4624
		x"0a",	--4625
		x"28",	--4626
		x"02",	--4627
		x"c1",	--4628
		x"02",	--4629
		x"c1",	--4630
		x"2e",	--4631
		x"2a",	--4632
		x"0f",	--4633
		x"3f",	--4634
		x"1c",	--4635
		x"81",	--4636
		x"42",	--4637
		x"1a",	--4638
		x"1c",	--4639
		x"8a",	--4640
		x"8a",	--4641
		x"8a",	--4642
		x"8a",	--4643
		x"81",	--4644
		x"44",	--4645
		x"81",	--4646
		x"46",	--4647
		x"0a",	--4648
		x"8a",	--4649
		x"8a",	--4650
		x"8a",	--4651
		x"8a",	--4652
		x"81",	--4653
		x"48",	--4654
		x"1c",	--4655
		x"42",	--4656
		x"1d",	--4657
		x"44",	--4658
		x"1c",	--4659
		x"46",	--4660
		x"1d",	--4661
		x"48",	--4662
		x"2c",	--4663
		x"1c",	--4664
		x"26",	--4665
		x"0e",	--4666
		x"e1",	--4667
		x"01",	--4668
		x"5e",	--4669
		x"26",	--4670
		x"4e",	--4671
		x"c1",	--4672
		x"03",	--4673
		x"06",	--4674
		x"c1",	--4675
		x"2a",	--4676
		x"03",	--4677
		x"91",	--4678
		x"26",	--4679
		x"30",	--4680
		x"11",	--4681
		x"04",	--4682
		x"11",	--4683
		x"04",	--4684
		x"1d",	--4685
		x"34",	--4686
		x"0e",	--4687
		x"1e",	--4688
		x"1f",	--4689
		x"3e",	--4690
		x"b0",	--4691
		x"de",	--4692
		x"21",	--4693
		x"81",	--4694
		x"2c",	--4695
		x"0d",	--4696
		x"7f",	--4697
		x"8f",	--4698
		x"91",	--4699
		x"3c",	--4700
		x"0e",	--4701
		x"0e",	--4702
		x"19",	--4703
		x"40",	--4704
		x"f7",	--4705
		x"81",	--4706
		x"3e",	--4707
		x"81",	--4708
		x"2c",	--4709
		x"07",	--4710
		x"0e",	--4711
		x"91",	--4712
		x"26",	--4713
		x"30",	--4714
		x"d1",	--4715
		x"2e",	--4716
		x"c1",	--4717
		x"2a",	--4718
		x"03",	--4719
		x"05",	--4720
		x"d1",	--4721
		x"2a",	--4722
		x"81",	--4723
		x"26",	--4724
		x"17",	--4725
		x"16",	--4726
		x"40",	--4727
		x"6e",	--4728
		x"4e",	--4729
		x"02",	--4730
		x"30",	--4731
		x"c2",	--4732
		x"1f",	--4733
		x"2c",	--4734
		x"31",	--4735
		x"4a",	--4736
		x"34",	--4737
		x"35",	--4738
		x"36",	--4739
		x"37",	--4740
		x"38",	--4741
		x"39",	--4742
		x"3a",	--4743
		x"3b",	--4744
		x"30",	--4745
		x"0d",	--4746
		x"0f",	--4747
		x"04",	--4748
		x"3d",	--4749
		x"03",	--4750
		x"3f",	--4751
		x"1f",	--4752
		x"0e",	--4753
		x"03",	--4754
		x"5d",	--4755
		x"3e",	--4756
		x"1e",	--4757
		x"0d",	--4758
		x"b0",	--4759
		x"da",	--4760
		x"3d",	--4761
		x"6d",	--4762
		x"02",	--4763
		x"3e",	--4764
		x"1e",	--4765
		x"5d",	--4766
		x"02",	--4767
		x"3f",	--4768
		x"1f",	--4769
		x"30",	--4770
		x"b0",	--4771
		x"14",	--4772
		x"0f",	--4773
		x"30",	--4774
		x"0b",	--4775
		x"0a",	--4776
		x"09",	--4777
		x"79",	--4778
		x"20",	--4779
		x"0a",	--4780
		x"0b",	--4781
		x"0c",	--4782
		x"0d",	--4783
		x"0e",	--4784
		x"0f",	--4785
		x"0c",	--4786
		x"0d",	--4787
		x"0d",	--4788
		x"06",	--4789
		x"02",	--4790
		x"0c",	--4791
		x"03",	--4792
		x"0c",	--4793
		x"0d",	--4794
		x"1e",	--4795
		x"19",	--4796
		x"f2",	--4797
		x"39",	--4798
		x"3a",	--4799
		x"3b",	--4800
		x"30",	--4801
		x"b0",	--4802
		x"4e",	--4803
		x"0e",	--4804
		x"0f",	--4805
		x"30",	--4806
		x"0b",	--4807
		x"0b",	--4808
		x"0f",	--4809
		x"06",	--4810
		x"3b",	--4811
		x"03",	--4812
		x"3e",	--4813
		x"3f",	--4814
		x"1e",	--4815
		x"0f",	--4816
		x"0d",	--4817
		x"05",	--4818
		x"5b",	--4819
		x"3c",	--4820
		x"3d",	--4821
		x"1c",	--4822
		x"0d",	--4823
		x"b0",	--4824
		x"4e",	--4825
		x"6b",	--4826
		x"04",	--4827
		x"3c",	--4828
		x"3d",	--4829
		x"1c",	--4830
		x"0d",	--4831
		x"5b",	--4832
		x"04",	--4833
		x"3e",	--4834
		x"3f",	--4835
		x"1e",	--4836
		x"0f",	--4837
		x"3b",	--4838
		x"30",	--4839
		x"b0",	--4840
		x"8e",	--4841
		x"0e",	--4842
		x"0f",	--4843
		x"30",	--4844
		x"7c",	--4845
		x"10",	--4846
		x"0d",	--4847
		x"0e",	--4848
		x"0f",	--4849
		x"0e",	--4850
		x"0e",	--4851
		x"02",	--4852
		x"0e",	--4853
		x"1f",	--4854
		x"1c",	--4855
		x"f8",	--4856
		x"30",	--4857
		x"b0",	--4858
		x"da",	--4859
		x"0f",	--4860
		x"30",	--4861
		x"07",	--4862
		x"06",	--4863
		x"05",	--4864
		x"04",	--4865
		x"30",	--4866
		x"40",	--4867
		x"04",	--4868
		x"05",	--4869
		x"06",	--4870
		x"07",	--4871
		x"08",	--4872
		x"09",	--4873
		x"0a",	--4874
		x"0b",	--4875
		x"0c",	--4876
		x"0d",	--4877
		x"0e",	--4878
		x"0f",	--4879
		x"08",	--4880
		x"09",	--4881
		x"0a",	--4882
		x"0b",	--4883
		x"0b",	--4884
		x"0e",	--4885
		x"08",	--4886
		x"0a",	--4887
		x"0b",	--4888
		x"05",	--4889
		x"09",	--4890
		x"08",	--4891
		x"02",	--4892
		x"08",	--4893
		x"05",	--4894
		x"08",	--4895
		x"09",	--4896
		x"0a",	--4897
		x"0b",	--4898
		x"1c",	--4899
		x"91",	--4900
		x"00",	--4901
		x"e5",	--4902
		x"21",	--4903
		x"34",	--4904
		x"35",	--4905
		x"36",	--4906
		x"37",	--4907
		x"30",	--4908
		x"0b",	--4909
		x"0a",	--4910
		x"09",	--4911
		x"08",	--4912
		x"18",	--4913
		x"0a",	--4914
		x"19",	--4915
		x"0c",	--4916
		x"1a",	--4917
		x"0e",	--4918
		x"1b",	--4919
		x"10",	--4920
		x"b0",	--4921
		x"fc",	--4922
		x"38",	--4923
		x"39",	--4924
		x"3a",	--4925
		x"3b",	--4926
		x"30",	--4927
		x"0b",	--4928
		x"0a",	--4929
		x"09",	--4930
		x"08",	--4931
		x"18",	--4932
		x"0a",	--4933
		x"19",	--4934
		x"0c",	--4935
		x"1a",	--4936
		x"0e",	--4937
		x"1b",	--4938
		x"10",	--4939
		x"b0",	--4940
		x"fc",	--4941
		x"0c",	--4942
		x"0d",	--4943
		x"0e",	--4944
		x"0f",	--4945
		x"38",	--4946
		x"39",	--4947
		x"3a",	--4948
		x"3b",	--4949
		x"30",	--4950
		x"0b",	--4951
		x"0a",	--4952
		x"09",	--4953
		x"08",	--4954
		x"07",	--4955
		x"18",	--4956
		x"0c",	--4957
		x"19",	--4958
		x"0e",	--4959
		x"1a",	--4960
		x"10",	--4961
		x"1b",	--4962
		x"12",	--4963
		x"b0",	--4964
		x"fc",	--4965
		x"17",	--4966
		x"14",	--4967
		x"87",	--4968
		x"00",	--4969
		x"87",	--4970
		x"02",	--4971
		x"87",	--4972
		x"04",	--4973
		x"87",	--4974
		x"06",	--4975
		x"37",	--4976
		x"38",	--4977
		x"39",	--4978
		x"3a",	--4979
		x"3b",	--4980
		x"30",	--4981
		x"00",	--4982
		x"32",	--4983
		x"f0",	--4984
		x"fd",	--4985
		x"57",	--4986
		x"69",	--4987
		x"69",	--4988
		x"67",	--4989
		x"66",	--4990
		x"72",	--4991
		x"61",	--4992
		x"6e",	--4993
		x"77",	--4994
		x"2e",	--4995
		x"69",	--4996
		x"20",	--4997
		x"69",	--4998
		x"65",	--4999
		x"0a",	--5000
		x"57",	--5001
		x"20",	--5002
		x"68",	--5003
		x"75",	--5004
		x"64",	--5005
		x"6e",	--5006
		x"74",	--5007
		x"73",	--5008
		x"65",	--5009
		x"74",	--5010
		x"61",	--5011
		x"0d",	--5012
		x"00",	--5013
		x"74",	--5014
		x"70",	--5015
		x"0a",	--5016
		x"65",	--5017
		x"72",	--5018
		x"72",	--5019
		x"20",	--5020
		x"69",	--5021
		x"73",	--5022
		x"6e",	--5023
		x"20",	--5024
		x"72",	--5025
		x"75",	--5026
		x"65",	--5027
		x"74",	--5028
		x"0a",	--5029
		x"63",	--5030
		x"72",	--5031
		x"65",	--5032
		x"74",	--5033
		x"75",	--5034
		x"61",	--5035
		x"65",	--5036
		x"0d",	--5037
		x"00",	--5038
		x"25",	--5039
		x"20",	--5040
		x"45",	--5041
		x"54",	--5042
		x"52",	--5043
		x"47",	--5044
		x"54",	--5045
		x"3c",	--5046
		x"49",	--5047
		x"45",	--5048
		x"55",	--5049
		x"3e",	--5050
		x"0a",	--5051
		x"25",	--5052
		x"20",	--5053
		x"64",	--5054
		x"0a",	--5055
		x"25",	--5056
		x"64",	--5057
		x"25",	--5058
		x"64",	--5059
		x"25",	--5060
		x"0d",	--5061
		x"00",	--5062
		x"64",	--5063
		x"25",	--5064
		x"0d",	--5065
		x"00",	--5066
		x"ba",	--5067
		x"e2",	--5068
		x"e8",	--5069
		x"f0",	--5070
		x"f8",	--5071
		x"00",	--5072
		x"d2",	--5073
		x"da",	--5074
		x"0d",	--5075
		x"3d",	--5076
		x"3d",	--5077
		x"3d",	--5078
		x"20",	--5079
		x"61",	--5080
		x"63",	--5081
		x"6c",	--5082
		x"4d",	--5083
		x"55",	--5084
		x"3d",	--5085
		x"3d",	--5086
		x"3d",	--5087
		x"0d",	--5088
		x"00",	--5089
		x"6e",	--5090
		x"65",	--5091
		x"61",	--5092
		x"74",	--5093
		x"76",	--5094
		x"20",	--5095
		x"6f",	--5096
		x"65",	--5097
		x"77",	--5098
		x"69",	--5099
		x"65",	--5100
		x"72",	--5101
		x"61",	--5102
		x"00",	--5103
		x"75",	--5104
		x"7a",	--5105
		x"72",	--5106
		x"70",	--5107
		x"6d",	--5108
		x"65",	--5109
		x"63",	--5110
		x"64",	--5111
		x"72",	--5112
		x"73",	--5113
		x"65",	--5114
		x"64",	--5115
		x"63",	--5116
		x"6e",	--5117
		x"72",	--5118
		x"6c",	--5119
		x"65",	--5120
		x"00",	--5121
		x"70",	--5122
		x"65",	--5123
		x"20",	--5124
		x"6f",	--5125
		x"66",	--5126
		x"67",	--5127
		x"72",	--5128
		x"74",	--5129
		x"6f",	--5130
		x"00",	--5131
		x"6f",	--5132
		x"74",	--5133
		x"6f",	--5134
		x"64",	--5135
		x"72",	--5136
		x"0d",	--5137
		x"00",	--5138
		x"20",	--5139
		x"00",	--5140
		x"63",	--5141
		x"77",	--5142
		x"69",	--5143
		x"65",	--5144
		x"0d",	--5145
		x"65",	--5146
		x"72",	--5147
		x"72",	--5148
		x"20",	--5149
		x"69",	--5150
		x"73",	--5151
		x"6e",	--5152
		x"20",	--5153
		x"72",	--5154
		x"75",	--5155
		x"65",	--5156
		x"74",	--5157
		x"0a",	--5158
		x"63",	--5159
		x"72",	--5160
		x"65",	--5161
		x"74",	--5162
		x"75",	--5163
		x"61",	--5164
		x"65",	--5165
		x"0d",	--5166
		x"00",	--5167
		x"25",	--5168
		x"20",	--5169
		x"45",	--5170
		x"49",	--5171
		x"54",	--5172
		x"52",	--5173
		x"56",	--5174
		x"4c",	--5175
		x"45",	--5176
		x"0a",	--5177
		x"72",	--5178
		x"25",	--5179
		x"20",	--5180
		x"3d",	--5181
		x"64",	--5182
		x"0a",	--5183
		x"09",	--5184
		x"73",	--5185
		x"52",	--5186
		x"47",	--5187
		x"53",	--5188
		x"45",	--5189
		x"0d",	--5190
		x"00",	--5191
		x"65",	--5192
		x"64",	--5193
		x"0d",	--5194
		x"25",	--5195
		x"20",	--5196
		x"73",	--5197
		x"6e",	--5198
		x"74",	--5199
		x"61",	--5200
		x"6e",	--5201
		x"6d",	--5202
		x"65",	--5203
		x"0d",	--5204
		x"00",	--5205
		x"63",	--5206
		x"25",	--5207
		x"0d",	--5208
		x"00",	--5209
		x"63",	--5210
		x"20",	--5211
		x"6f",	--5212
		x"73",	--5213
		x"63",	--5214
		x"20",	--5215
		x"6f",	--5216
		x"6d",	--5217
		x"6e",	--5218
		x"0d",	--5219
		x"00",	--5220
		x"a2",	--5221
		x"d0",	--5222
		x"d0",	--5223
		x"d0",	--5224
		x"d0",	--5225
		x"d0",	--5226
		x"d0",	--5227
		x"d0",	--5228
		x"d0",	--5229
		x"d0",	--5230
		x"d0",	--5231
		x"d0",	--5232
		x"d0",	--5233
		x"d0",	--5234
		x"d0",	--5235
		x"d0",	--5236
		x"d0",	--5237
		x"d0",	--5238
		x"d0",	--5239
		x"d0",	--5240
		x"d0",	--5241
		x"d0",	--5242
		x"d0",	--5243
		x"d0",	--5244
		x"d0",	--5245
		x"d0",	--5246
		x"d0",	--5247
		x"d0",	--5248
		x"d0",	--5249
		x"94",	--5250
		x"d0",	--5251
		x"d0",	--5252
		x"d0",	--5253
		x"d0",	--5254
		x"d0",	--5255
		x"d0",	--5256
		x"d0",	--5257
		x"d0",	--5258
		x"d0",	--5259
		x"d0",	--5260
		x"d0",	--5261
		x"d0",	--5262
		x"d0",	--5263
		x"d0",	--5264
		x"d0",	--5265
		x"d0",	--5266
		x"d0",	--5267
		x"d0",	--5268
		x"d0",	--5269
		x"d0",	--5270
		x"d0",	--5271
		x"d0",	--5272
		x"d0",	--5273
		x"d0",	--5274
		x"d0",	--5275
		x"d0",	--5276
		x"d0",	--5277
		x"d0",	--5278
		x"d0",	--5279
		x"d0",	--5280
		x"d0",	--5281
		x"86",	--5282
		x"78",	--5283
		x"6a",	--5284
		x"d0",	--5285
		x"d0",	--5286
		x"d0",	--5287
		x"d0",	--5288
		x"d0",	--5289
		x"d0",	--5290
		x"d0",	--5291
		x"52",	--5292
		x"d0",	--5293
		x"40",	--5294
		x"d0",	--5295
		x"d0",	--5296
		x"d0",	--5297
		x"d0",	--5298
		x"24",	--5299
		x"d0",	--5300
		x"d0",	--5301
		x"d0",	--5302
		x"16",	--5303
		x"04",	--5304
		x"30",	--5305
		x"32",	--5306
		x"34",	--5307
		x"36",	--5308
		x"38",	--5309
		x"61",	--5310
		x"63",	--5311
		x"65",	--5312
		x"00",	--5313
		x"00",	--5314
		x"00",	--5315
		x"00",	--5316
		x"00",	--5317
		x"00",	--5318
		x"02",	--5319
		x"03",	--5320
		x"03",	--5321
		x"04",	--5322
		x"04",	--5323
		x"04",	--5324
		x"04",	--5325
		x"05",	--5326
		x"05",	--5327
		x"05",	--5328
		x"05",	--5329
		x"05",	--5330
		x"05",	--5331
		x"05",	--5332
		x"05",	--5333
		x"06",	--5334
		x"06",	--5335
		x"06",	--5336
		x"06",	--5337
		x"06",	--5338
		x"06",	--5339
		x"06",	--5340
		x"06",	--5341
		x"06",	--5342
		x"06",	--5343
		x"06",	--5344
		x"06",	--5345
		x"06",	--5346
		x"06",	--5347
		x"06",	--5348
		x"06",	--5349
		x"07",	--5350
		x"07",	--5351
		x"07",	--5352
		x"07",	--5353
		x"07",	--5354
		x"07",	--5355
		x"07",	--5356
		x"07",	--5357
		x"07",	--5358
		x"07",	--5359
		x"07",	--5360
		x"07",	--5361
		x"07",	--5362
		x"07",	--5363
		x"07",	--5364
		x"07",	--5365
		x"07",	--5366
		x"07",	--5367
		x"07",	--5368
		x"07",	--5369
		x"07",	--5370
		x"07",	--5371
		x"07",	--5372
		x"07",	--5373
		x"07",	--5374
		x"07",	--5375
		x"07",	--5376
		x"07",	--5377
		x"07",	--5378
		x"07",	--5379
		x"07",	--5380
		x"07",	--5381
		x"08",	--5382
		x"08",	--5383
		x"08",	--5384
		x"08",	--5385
		x"08",	--5386
		x"08",	--5387
		x"08",	--5388
		x"08",	--5389
		x"08",	--5390
		x"08",	--5391
		x"08",	--5392
		x"08",	--5393
		x"08",	--5394
		x"08",	--5395
		x"08",	--5396
		x"08",	--5397
		x"08",	--5398
		x"08",	--5399
		x"08",	--5400
		x"08",	--5401
		x"08",	--5402
		x"08",	--5403
		x"08",	--5404
		x"08",	--5405
		x"08",	--5406
		x"08",	--5407
		x"08",	--5408
		x"08",	--5409
		x"08",	--5410
		x"08",	--5411
		x"08",	--5412
		x"08",	--5413
		x"08",	--5414
		x"08",	--5415
		x"08",	--5416
		x"08",	--5417
		x"08",	--5418
		x"08",	--5419
		x"08",	--5420
		x"08",	--5421
		x"08",	--5422
		x"08",	--5423
		x"08",	--5424
		x"08",	--5425
		x"08",	--5426
		x"08",	--5427
		x"08",	--5428
		x"08",	--5429
		x"08",	--5430
		x"08",	--5431
		x"08",	--5432
		x"08",	--5433
		x"08",	--5434
		x"08",	--5435
		x"08",	--5436
		x"08",	--5437
		x"08",	--5438
		x"08",	--5439
		x"08",	--5440
		x"08",	--5441
		x"08",	--5442
		x"08",	--5443
		x"08",	--5444
		x"08",	--5445
		x"28",	--5446
		x"75",	--5447
		x"6c",	--5448
		x"00",	--5449
		x"ff",	--5450
		x"ff",	--5451
		x"68",	--5452
		x"6c",	--5453
		x"00",	--5454
		x"ff",	--5455
		x"ff",	--5456
		x"ff",	--5457
		x"ff",	--5458
		x"ff",	--5459
		x"ff",	--5460
		x"ff",	--5461
		x"ff",	--5462
		x"ff",	--5463
		x"ff",	--5464
		x"ff",	--5465
		x"ff",	--5466
		x"ff",	--5467
		x"ff",	--5468
		x"ff",	--5469
		x"ff",	--5470
		x"ff",	--5471
		x"ff",	--5472
		x"ff",	--5473
		x"ff",	--5474
		x"ff",	--5475
		x"ff",	--5476
		x"ff",	--5477
		x"ff",	--5478
		x"ff",	--5479
		x"ff",	--5480
		x"ff",	--5481
		x"ff",	--5482
		x"ff",	--5483
		x"ff",	--5484
		x"ff",	--5485
		x"ff",	--5486
		x"ff",	--5487
		x"ff",	--5488
		x"ff",	--5489
		x"ff",	--5490
		x"ff",	--5491
		x"ff",	--5492
		x"ff",	--5493
		x"ff",	--5494
		x"ff",	--5495
		x"ff",	--5496
		x"ff",	--5497
		x"ff",	--5498
		x"ff",	--5499
		x"ff",	--5500
		x"ff",	--5501
		x"ff",	--5502
		x"ff",	--5503
		x"ff",	--5504
		x"ff",	--5505
		x"ff",	--5506
		x"ff",	--5507
		x"ff",	--5508
		x"ff",	--5509
		x"ff",	--5510
		x"ff",	--5511
		x"ff",	--5512
		x"ff",	--5513
		x"ff",	--5514
		x"ff",	--5515
		x"ff",	--5516
		x"ff",	--5517
		x"ff",	--5518
		x"ff",	--5519
		x"ff",	--5520
		x"ff",	--5521
		x"ff",	--5522
		x"ff",	--5523
		x"ff",	--5524
		x"ff",	--5525
		x"ff",	--5526
		x"ff",	--5527
		x"ff",	--5528
		x"ff",	--5529
		x"ff",	--5530
		x"ff",	--5531
		x"ff",	--5532
		x"ff",	--5533
		x"ff",	--5534
		x"ff",	--5535
		x"ff",	--5536
		x"ff",	--5537
		x"ff",	--5538
		x"ff",	--5539
		x"ff",	--5540
		x"ff",	--5541
		x"ff",	--5542
		x"ff",	--5543
		x"ff",	--5544
		x"ff",	--5545
		x"ff",	--5546
		x"ff",	--5547
		x"ff",	--5548
		x"ff",	--5549
		x"ff",	--5550
		x"ff",	--5551
		x"ff",	--5552
		x"ff",	--5553
		x"ff",	--5554
		x"ff",	--5555
		x"ff",	--5556
		x"ff",	--5557
		x"ff",	--5558
		x"ff",	--5559
		x"ff",	--5560
		x"ff",	--5561
		x"ff",	--5562
		x"ff",	--5563
		x"ff",	--5564
		x"ff",	--5565
		x"ff",	--5566
		x"ff",	--5567
		x"ff",	--5568
		x"ff",	--5569
		x"ff",	--5570
		x"ff",	--5571
		x"ff",	--5572
		x"ff",	--5573
		x"ff",	--5574
		x"ff",	--5575
		x"ff",	--5576
		x"ff",	--5577
		x"ff",	--5578
		x"ff",	--5579
		x"ff",	--5580
		x"ff",	--5581
		x"ff",	--5582
		x"ff",	--5583
		x"ff",	--5584
		x"ff",	--5585
		x"ff",	--5586
		x"ff",	--5587
		x"ff",	--5588
		x"ff",	--5589
		x"ff",	--5590
		x"ff",	--5591
		x"ff",	--5592
		x"ff",	--5593
		x"ff",	--5594
		x"ff",	--5595
		x"ff",	--5596
		x"ff",	--5597
		x"ff",	--5598
		x"ff",	--5599
		x"ff",	--5600
		x"ff",	--5601
		x"ff",	--5602
		x"ff",	--5603
		x"ff",	--5604
		x"ff",	--5605
		x"ff",	--5606
		x"ff",	--5607
		x"ff",	--5608
		x"ff",	--5609
		x"ff",	--5610
		x"ff",	--5611
		x"ff",	--5612
		x"ff",	--5613
		x"ff",	--5614
		x"ff",	--5615
		x"ff",	--5616
		x"ff",	--5617
		x"ff",	--5618
		x"ff",	--5619
		x"ff",	--5620
		x"ff",	--5621
		x"ff",	--5622
		x"ff",	--5623
		x"ff",	--5624
		x"ff",	--5625
		x"ff",	--5626
		x"ff",	--5627
		x"ff",	--5628
		x"ff",	--5629
		x"ff",	--5630
		x"ff",	--5631
		x"ff",	--5632
		x"ff",	--5633
		x"ff",	--5634
		x"ff",	--5635
		x"ff",	--5636
		x"ff",	--5637
		x"ff",	--5638
		x"ff",	--5639
		x"ff",	--5640
		x"ff",	--5641
		x"ff",	--5642
		x"ff",	--5643
		x"ff",	--5644
		x"ff",	--5645
		x"ff",	--5646
		x"ff",	--5647
		x"ff",	--5648
		x"ff",	--5649
		x"ff",	--5650
		x"ff",	--5651
		x"ff",	--5652
		x"ff",	--5653
		x"ff",	--5654
		x"ff",	--5655
		x"ff",	--5656
		x"ff",	--5657
		x"ff",	--5658
		x"ff",	--5659
		x"ff",	--5660
		x"ff",	--5661
		x"ff",	--5662
		x"ff",	--5663
		x"ff",	--5664
		x"ff",	--5665
		x"ff",	--5666
		x"ff",	--5667
		x"ff",	--5668
		x"ff",	--5669
		x"ff",	--5670
		x"ff",	--5671
		x"ff",	--5672
		x"ff",	--5673
		x"ff",	--5674
		x"ff",	--5675
		x"ff",	--5676
		x"ff",	--5677
		x"ff",	--5678
		x"ff",	--5679
		x"ff",	--5680
		x"ff",	--5681
		x"ff",	--5682
		x"ff",	--5683
		x"ff",	--5684
		x"ff",	--5685
		x"ff",	--5686
		x"ff",	--5687
		x"ff",	--5688
		x"ff",	--5689
		x"ff",	--5690
		x"ff",	--5691
		x"ff",	--5692
		x"ff",	--5693
		x"ff",	--5694
		x"ff",	--5695
		x"ff",	--5696
		x"ff",	--5697
		x"ff",	--5698
		x"ff",	--5699
		x"ff",	--5700
		x"ff",	--5701
		x"ff",	--5702
		x"ff",	--5703
		x"ff",	--5704
		x"ff",	--5705
		x"ff",	--5706
		x"ff",	--5707
		x"ff",	--5708
		x"ff",	--5709
		x"ff",	--5710
		x"ff",	--5711
		x"ff",	--5712
		x"ff",	--5713
		x"ff",	--5714
		x"ff",	--5715
		x"ff",	--5716
		x"ff",	--5717
		x"ff",	--5718
		x"ff",	--5719
		x"ff",	--5720
		x"ff",	--5721
		x"ff",	--5722
		x"ff",	--5723
		x"ff",	--5724
		x"ff",	--5725
		x"ff",	--5726
		x"ff",	--5727
		x"ff",	--5728
		x"ff",	--5729
		x"ff",	--5730
		x"ff",	--5731
		x"ff",	--5732
		x"ff",	--5733
		x"ff",	--5734
		x"ff",	--5735
		x"ff",	--5736
		x"ff",	--5737
		x"ff",	--5738
		x"ff",	--5739
		x"ff",	--5740
		x"ff",	--5741
		x"ff",	--5742
		x"ff",	--5743
		x"ff",	--5744
		x"ff",	--5745
		x"ff",	--5746
		x"ff",	--5747
		x"ff",	--5748
		x"ff",	--5749
		x"ff",	--5750
		x"ff",	--5751
		x"ff",	--5752
		x"ff",	--5753
		x"ff",	--5754
		x"ff",	--5755
		x"ff",	--5756
		x"ff",	--5757
		x"ff",	--5758
		x"ff",	--5759
		x"ff",	--5760
		x"ff",	--5761
		x"ff",	--5762
		x"ff",	--5763
		x"ff",	--5764
		x"ff",	--5765
		x"ff",	--5766
		x"ff",	--5767
		x"ff",	--5768
		x"ff",	--5769
		x"ff",	--5770
		x"ff",	--5771
		x"ff",	--5772
		x"ff",	--5773
		x"ff",	--5774
		x"ff",	--5775
		x"ff",	--5776
		x"ff",	--5777
		x"ff",	--5778
		x"ff",	--5779
		x"ff",	--5780
		x"ff",	--5781
		x"ff",	--5782
		x"ff",	--5783
		x"ff",	--5784
		x"ff",	--5785
		x"ff",	--5786
		x"ff",	--5787
		x"ff",	--5788
		x"ff",	--5789
		x"ff",	--5790
		x"ff",	--5791
		x"ff",	--5792
		x"ff",	--5793
		x"ff",	--5794
		x"ff",	--5795
		x"ff",	--5796
		x"ff",	--5797
		x"ff",	--5798
		x"ff",	--5799
		x"ff",	--5800
		x"ff",	--5801
		x"ff",	--5802
		x"ff",	--5803
		x"ff",	--5804
		x"ff",	--5805
		x"ff",	--5806
		x"ff",	--5807
		x"ff",	--5808
		x"ff",	--5809
		x"ff",	--5810
		x"ff",	--5811
		x"ff",	--5812
		x"ff",	--5813
		x"ff",	--5814
		x"ff",	--5815
		x"ff",	--5816
		x"ff",	--5817
		x"ff",	--5818
		x"ff",	--5819
		x"ff",	--5820
		x"ff",	--5821
		x"ff",	--5822
		x"ff",	--5823
		x"ff",	--5824
		x"ff",	--5825
		x"ff",	--5826
		x"ff",	--5827
		x"ff",	--5828
		x"ff",	--5829
		x"ff",	--5830
		x"ff",	--5831
		x"ff",	--5832
		x"ff",	--5833
		x"ff",	--5834
		x"ff",	--5835
		x"ff",	--5836
		x"ff",	--5837
		x"ff",	--5838
		x"ff",	--5839
		x"ff",	--5840
		x"ff",	--5841
		x"ff",	--5842
		x"ff",	--5843
		x"ff",	--5844
		x"ff",	--5845
		x"ff",	--5846
		x"ff",	--5847
		x"ff",	--5848
		x"ff",	--5849
		x"ff",	--5850
		x"ff",	--5851
		x"ff",	--5852
		x"ff",	--5853
		x"ff",	--5854
		x"ff",	--5855
		x"ff",	--5856
		x"ff",	--5857
		x"ff",	--5858
		x"ff",	--5859
		x"ff",	--5860
		x"ff",	--5861
		x"ff",	--5862
		x"ff",	--5863
		x"ff",	--5864
		x"ff",	--5865
		x"ff",	--5866
		x"ff",	--5867
		x"ff",	--5868
		x"ff",	--5869
		x"ff",	--5870
		x"ff",	--5871
		x"ff",	--5872
		x"ff",	--5873
		x"ff",	--5874
		x"ff",	--5875
		x"ff",	--5876
		x"ff",	--5877
		x"ff",	--5878
		x"ff",	--5879
		x"ff",	--5880
		x"ff",	--5881
		x"ff",	--5882
		x"ff",	--5883
		x"ff",	--5884
		x"ff",	--5885
		x"ff",	--5886
		x"ff",	--5887
		x"ff",	--5888
		x"ff",	--5889
		x"ff",	--5890
		x"ff",	--5891
		x"ff",	--5892
		x"ff",	--5893
		x"ff",	--5894
		x"ff",	--5895
		x"ff",	--5896
		x"ff",	--5897
		x"ff",	--5898
		x"ff",	--5899
		x"ff",	--5900
		x"ff",	--5901
		x"ff",	--5902
		x"ff",	--5903
		x"ff",	--5904
		x"ff",	--5905
		x"ff",	--5906
		x"ff",	--5907
		x"ff",	--5908
		x"ff",	--5909
		x"ff",	--5910
		x"ff",	--5911
		x"ff",	--5912
		x"ff",	--5913
		x"ff",	--5914
		x"ff",	--5915
		x"ff",	--5916
		x"ff",	--5917
		x"ff",	--5918
		x"ff",	--5919
		x"ff",	--5920
		x"ff",	--5921
		x"ff",	--5922
		x"ff",	--5923
		x"ff",	--5924
		x"ff",	--5925
		x"ff",	--5926
		x"ff",	--5927
		x"ff",	--5928
		x"ff",	--5929
		x"ff",	--5930
		x"ff",	--5931
		x"ff",	--5932
		x"ff",	--5933
		x"ff",	--5934
		x"ff",	--5935
		x"ff",	--5936
		x"ff",	--5937
		x"ff",	--5938
		x"ff",	--5939
		x"ff",	--5940
		x"ff",	--5941
		x"ff",	--5942
		x"ff",	--5943
		x"ff",	--5944
		x"ff",	--5945
		x"ff",	--5946
		x"ff",	--5947
		x"ff",	--5948
		x"ff",	--5949
		x"ff",	--5950
		x"ff",	--5951
		x"ff",	--5952
		x"ff",	--5953
		x"ff",	--5954
		x"ff",	--5955
		x"ff",	--5956
		x"ff",	--5957
		x"ff",	--5958
		x"ff",	--5959
		x"ff",	--5960
		x"ff",	--5961
		x"ff",	--5962
		x"ff",	--5963
		x"ff",	--5964
		x"ff",	--5965
		x"ff",	--5966
		x"ff",	--5967
		x"ff",	--5968
		x"ff",	--5969
		x"ff",	--5970
		x"ff",	--5971
		x"ff",	--5972
		x"ff",	--5973
		x"ff",	--5974
		x"ff",	--5975
		x"ff",	--5976
		x"ff",	--5977
		x"ff",	--5978
		x"ff",	--5979
		x"ff",	--5980
		x"ff",	--5981
		x"ff",	--5982
		x"ff",	--5983
		x"ff",	--5984
		x"ff",	--5985
		x"ff",	--5986
		x"ff",	--5987
		x"ff",	--5988
		x"ff",	--5989
		x"ff",	--5990
		x"ff",	--5991
		x"ff",	--5992
		x"ff",	--5993
		x"ff",	--5994
		x"ff",	--5995
		x"ff",	--5996
		x"ff",	--5997
		x"ff",	--5998
		x"ff",	--5999
		x"ff",	--6000
		x"ff",	--6001
		x"ff",	--6002
		x"ff",	--6003
		x"ff",	--6004
		x"ff",	--6005
		x"ff",	--6006
		x"ff",	--6007
		x"ff",	--6008
		x"ff",	--6009
		x"ff",	--6010
		x"ff",	--6011
		x"ff",	--6012
		x"ff",	--6013
		x"ff",	--6014
		x"ff",	--6015
		x"ff",	--6016
		x"ff",	--6017
		x"ff",	--6018
		x"ff",	--6019
		x"ff",	--6020
		x"ff",	--6021
		x"ff",	--6022
		x"ff",	--6023
		x"ff",	--6024
		x"ff",	--6025
		x"ff",	--6026
		x"ff",	--6027
		x"ff",	--6028
		x"ff",	--6029
		x"ff",	--6030
		x"ff",	--6031
		x"ff",	--6032
		x"ff",	--6033
		x"ff",	--6034
		x"ff",	--6035
		x"ff",	--6036
		x"ff",	--6037
		x"ff",	--6038
		x"ff",	--6039
		x"ff",	--6040
		x"ff",	--6041
		x"ff",	--6042
		x"ff",	--6043
		x"ff",	--6044
		x"ff",	--6045
		x"ff",	--6046
		x"ff",	--6047
		x"ff",	--6048
		x"ff",	--6049
		x"ff",	--6050
		x"ff",	--6051
		x"ff",	--6052
		x"ff",	--6053
		x"ff",	--6054
		x"ff",	--6055
		x"ff",	--6056
		x"ff",	--6057
		x"ff",	--6058
		x"ff",	--6059
		x"ff",	--6060
		x"ff",	--6061
		x"ff",	--6062
		x"ff",	--6063
		x"ff",	--6064
		x"ff",	--6065
		x"ff",	--6066
		x"ff",	--6067
		x"ff",	--6068
		x"ff",	--6069
		x"ff",	--6070
		x"ff",	--6071
		x"ff",	--6072
		x"ff",	--6073
		x"ff",	--6074
		x"ff",	--6075
		x"ff",	--6076
		x"ff",	--6077
		x"ff",	--6078
		x"ff",	--6079
		x"ff",	--6080
		x"ff",	--6081
		x"ff",	--6082
		x"ff",	--6083
		x"ff",	--6084
		x"ff",	--6085
		x"ff",	--6086
		x"ff",	--6087
		x"ff",	--6088
		x"ff",	--6089
		x"ff",	--6090
		x"ff",	--6091
		x"ff",	--6092
		x"ff",	--6093
		x"ff",	--6094
		x"ff",	--6095
		x"ff",	--6096
		x"ff",	--6097
		x"ff",	--6098
		x"ff",	--6099
		x"ff",	--6100
		x"ff",	--6101
		x"ff",	--6102
		x"ff",	--6103
		x"ff",	--6104
		x"ff",	--6105
		x"ff",	--6106
		x"ff",	--6107
		x"ff",	--6108
		x"ff",	--6109
		x"ff",	--6110
		x"ff",	--6111
		x"ff",	--6112
		x"ff",	--6113
		x"ff",	--6114
		x"ff",	--6115
		x"ff",	--6116
		x"ff",	--6117
		x"ff",	--6118
		x"ff",	--6119
		x"ff",	--6120
		x"ff",	--6121
		x"ff",	--6122
		x"ff",	--6123
		x"ff",	--6124
		x"ff",	--6125
		x"ff",	--6126
		x"ff",	--6127
		x"ff",	--6128
		x"ff",	--6129
		x"ff",	--6130
		x"ff",	--6131
		x"ff",	--6132
		x"ff",	--6133
		x"ff",	--6134
		x"ff",	--6135
		x"ff",	--6136
		x"ff",	--6137
		x"ff",	--6138
		x"ff",	--6139
		x"ff",	--6140
		x"ff",	--6141
		x"ff",	--6142
		x"ff",	--6143
		x"ff",	--6144
		x"ff",	--6145
		x"ff",	--6146
		x"ff",	--6147
		x"ff",	--6148
		x"ff",	--6149
		x"ff",	--6150
		x"ff",	--6151
		x"ff",	--6152
		x"ff",	--6153
		x"ff",	--6154
		x"ff",	--6155
		x"ff",	--6156
		x"ff",	--6157
		x"ff",	--6158
		x"ff",	--6159
		x"ff",	--6160
		x"ff",	--6161
		x"ff",	--6162
		x"ff",	--6163
		x"ff",	--6164
		x"ff",	--6165
		x"ff",	--6166
		x"ff",	--6167
		x"ff",	--6168
		x"ff",	--6169
		x"ff",	--6170
		x"ff",	--6171
		x"ff",	--6172
		x"ff",	--6173
		x"ff",	--6174
		x"ff",	--6175
		x"ff",	--6176
		x"ff",	--6177
		x"ff",	--6178
		x"ff",	--6179
		x"ff",	--6180
		x"ff",	--6181
		x"ff",	--6182
		x"ff",	--6183
		x"ff",	--6184
		x"ff",	--6185
		x"ff",	--6186
		x"ff",	--6187
		x"ff",	--6188
		x"ff",	--6189
		x"ff",	--6190
		x"ff",	--6191
		x"ff",	--6192
		x"ff",	--6193
		x"ff",	--6194
		x"ff",	--6195
		x"ff",	--6196
		x"ff",	--6197
		x"ff",	--6198
		x"ff",	--6199
		x"ff",	--6200
		x"ff",	--6201
		x"ff",	--6202
		x"ff",	--6203
		x"ff",	--6204
		x"ff",	--6205
		x"ff",	--6206
		x"ff",	--6207
		x"ff",	--6208
		x"ff",	--6209
		x"ff",	--6210
		x"ff",	--6211
		x"ff",	--6212
		x"ff",	--6213
		x"ff",	--6214
		x"ff",	--6215
		x"ff",	--6216
		x"ff",	--6217
		x"ff",	--6218
		x"ff",	--6219
		x"ff",	--6220
		x"ff",	--6221
		x"ff",	--6222
		x"ff",	--6223
		x"ff",	--6224
		x"ff",	--6225
		x"ff",	--6226
		x"ff",	--6227
		x"ff",	--6228
		x"ff",	--6229
		x"ff",	--6230
		x"ff",	--6231
		x"ff",	--6232
		x"ff",	--6233
		x"ff",	--6234
		x"ff",	--6235
		x"ff",	--6236
		x"ff",	--6237
		x"ff",	--6238
		x"ff",	--6239
		x"ff",	--6240
		x"ff",	--6241
		x"ff",	--6242
		x"ff",	--6243
		x"ff",	--6244
		x"ff",	--6245
		x"ff",	--6246
		x"ff",	--6247
		x"ff",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"ff",	--6252
		x"ff",	--6253
		x"ff",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"60",	--8176
		x"60",	--8177
		x"60",	--8178
		x"60",	--8179
		x"60",	--8180
		x"60",	--8181
		x"60",	--8182
		x"ac",	--8183
		x"fe",	--8184
		x"60",	--8185
		x"60",	--8186
		x"60",	--8187
		x"60",	--8188
		x"60",	--8189
		x"60",	--8190
		x"00");	--8191
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"ea",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"ce",	--44
		x"12",	--45
		x"c9",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"e7",	--50
		x"12",	--51
		x"cd",	--52
		x"53",	--53
		x"40",	--54
		x"e7",	--55
		x"40",	--56
		x"c5",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"c9",	--61
		x"40",	--62
		x"e7",	--63
		x"40",	--64
		x"c6",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"c9",	--69
		x"40",	--70
		x"e7",	--71
		x"40",	--72
		x"c7",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"c9",	--77
		x"40",	--78
		x"e7",	--79
		x"40",	--80
		x"c2",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"c9",	--85
		x"40",	--86
		x"e7",	--87
		x"40",	--88
		x"c3",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"c9",	--93
		x"40",	--94
		x"e7",	--95
		x"40",	--96
		x"c4",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"c9",	--101
		x"40",	--102
		x"e7",	--103
		x"40",	--104
		x"c2",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"c9",	--109
		x"40",	--110
		x"e8",	--111
		x"40",	--112
		x"c2",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"c9",	--117
		x"40",	--118
		x"e8",	--119
		x"40",	--120
		x"c2",	--121
		x"40",	--122
		x"00",	--123
		x"12",	--124
		x"c9",	--125
		x"43",	--126
		x"43",	--127
		x"12",	--128
		x"c9",	--129
		x"43",	--130
		x"40",	--131
		x"4e",	--132
		x"40",	--133
		x"01",	--134
		x"41",	--135
		x"50",	--136
		x"00",	--137
		x"12",	--138
		x"c8",	--139
		x"41",	--140
		x"50",	--141
		x"00",	--142
		x"12",	--143
		x"c8",	--144
		x"43",	--145
		x"40",	--146
		x"4e",	--147
		x"40",	--148
		x"01",	--149
		x"41",	--150
		x"50",	--151
		x"00",	--152
		x"12",	--153
		x"c8",	--154
		x"41",	--155
		x"50",	--156
		x"00",	--157
		x"12",	--158
		x"c8",	--159
		x"41",	--160
		x"50",	--161
		x"00",	--162
		x"41",	--163
		x"50",	--164
		x"00",	--165
		x"12",	--166
		x"c3",	--167
		x"40",	--168
		x"01",	--169
		x"41",	--170
		x"52",	--171
		x"12",	--172
		x"cb",	--173
		x"40",	--174
		x"01",	--175
		x"41",	--176
		x"53",	--177
		x"12",	--178
		x"cb",	--179
		x"41",	--180
		x"53",	--181
		x"41",	--182
		x"52",	--183
		x"12",	--184
		x"c4",	--185
		x"41",	--186
		x"50",	--187
		x"00",	--188
		x"41",	--189
		x"50",	--190
		x"00",	--191
		x"12",	--192
		x"c4",	--193
		x"12",	--194
		x"ca",	--195
		x"40",	--196
		x"01",	--197
		x"41",	--198
		x"12",	--199
		x"cb",	--200
		x"41",	--201
		x"12",	--202
		x"c2",	--203
		x"40",	--204
		x"00",	--205
		x"40",	--206
		x"17",	--207
		x"41",	--208
		x"12",	--209
		x"cb",	--210
		x"43",	--211
		x"43",	--212
		x"43",	--213
		x"41",	--214
		x"50",	--215
		x"00",	--216
		x"12",	--217
		x"c2",	--218
		x"43",	--219
		x"43",	--220
		x"43",	--221
		x"41",	--222
		x"50",	--223
		x"00",	--224
		x"12",	--225
		x"c2",	--226
		x"41",	--227
		x"50",	--228
		x"00",	--229
		x"41",	--230
		x"50",	--231
		x"00",	--232
		x"12",	--233
		x"c2",	--234
		x"40",	--235
		x"ff",	--236
		x"00",	--237
		x"d2",	--238
		x"43",	--239
		x"12",	--240
		x"cf",	--241
		x"93",	--242
		x"27",	--243
		x"12",	--244
		x"cf",	--245
		x"92",	--246
		x"24",	--247
		x"90",	--248
		x"00",	--249
		x"20",	--250
		x"12",	--251
		x"e8",	--252
		x"12",	--253
		x"cd",	--254
		x"53",	--255
		x"40",	--256
		x"00",	--257
		x"51",	--258
		x"5f",	--259
		x"43",	--260
		x"00",	--261
		x"4f",	--262
		x"41",	--263
		x"00",	--264
		x"12",	--265
		x"c9",	--266
		x"43",	--267
		x"3f",	--268
		x"93",	--269
		x"27",	--270
		x"53",	--271
		x"12",	--272
		x"e8",	--273
		x"12",	--274
		x"cd",	--275
		x"53",	--276
		x"3f",	--277
		x"90",	--278
		x"00",	--279
		x"2f",	--280
		x"93",	--281
		x"02",	--282
		x"24",	--283
		x"4f",	--284
		x"11",	--285
		x"12",	--286
		x"12",	--287
		x"e8",	--288
		x"4f",	--289
		x"00",	--290
		x"12",	--291
		x"cd",	--292
		x"52",	--293
		x"41",	--294
		x"00",	--295
		x"40",	--296
		x"00",	--297
		x"51",	--298
		x"5b",	--299
		x"4f",	--300
		x"00",	--301
		x"53",	--302
		x"3f",	--303
		x"40",	--304
		x"e6",	--305
		x"4f",	--306
		x"02",	--307
		x"41",	--308
		x"12",	--309
		x"12",	--310
		x"82",	--311
		x"4f",	--312
		x"4e",	--313
		x"93",	--314
		x"38",	--315
		x"41",	--316
		x"4b",	--317
		x"00",	--318
		x"12",	--319
		x"c7",	--320
		x"4f",	--321
		x"93",	--322
		x"24",	--323
		x"41",	--324
		x"4b",	--325
		x"00",	--326
		x"4d",	--327
		x"00",	--328
		x"12",	--329
		x"c7",	--330
		x"4f",	--331
		x"41",	--332
		x"00",	--333
		x"42",	--334
		x"02",	--335
		x"12",	--336
		x"cb",	--337
		x"43",	--338
		x"52",	--339
		x"41",	--340
		x"41",	--341
		x"41",	--342
		x"40",	--343
		x"00",	--344
		x"40",	--345
		x"17",	--346
		x"3f",	--347
		x"40",	--348
		x"17",	--349
		x"3f",	--350
		x"41",	--351
		x"43",	--352
		x"41",	--353
		x"43",	--354
		x"41",	--355
		x"40",	--356
		x"c0",	--357
		x"01",	--358
		x"40",	--359
		x"00",	--360
		x"01",	--361
		x"40",	--362
		x"02",	--363
		x"01",	--364
		x"12",	--365
		x"e6",	--366
		x"12",	--367
		x"cd",	--368
		x"43",	--369
		x"01",	--370
		x"40",	--371
		x"e7",	--372
		x"00",	--373
		x"12",	--374
		x"cd",	--375
		x"53",	--376
		x"43",	--377
		x"41",	--378
		x"12",	--379
		x"c6",	--380
		x"41",	--381
		x"12",	--382
		x"12",	--383
		x"43",	--384
		x"40",	--385
		x"3f",	--386
		x"4a",	--387
		x"4b",	--388
		x"42",	--389
		x"02",	--390
		x"12",	--391
		x"c8",	--392
		x"4a",	--393
		x"4b",	--394
		x"42",	--395
		x"02",	--396
		x"12",	--397
		x"c8",	--398
		x"12",	--399
		x"e7",	--400
		x"12",	--401
		x"cd",	--402
		x"53",	--403
		x"41",	--404
		x"41",	--405
		x"41",	--406
		x"4f",	--407
		x"02",	--408
		x"4e",	--409
		x"02",	--410
		x"41",	--411
		x"12",	--412
		x"12",	--413
		x"83",	--414
		x"4f",	--415
		x"4e",	--416
		x"93",	--417
		x"02",	--418
		x"24",	--419
		x"90",	--420
		x"00",	--421
		x"38",	--422
		x"20",	--423
		x"41",	--424
		x"4b",	--425
		x"00",	--426
		x"12",	--427
		x"c7",	--428
		x"4f",	--429
		x"41",	--430
		x"4b",	--431
		x"00",	--432
		x"12",	--433
		x"c7",	--434
		x"4f",	--435
		x"12",	--436
		x"12",	--437
		x"12",	--438
		x"e7",	--439
		x"12",	--440
		x"cd",	--441
		x"50",	--442
		x"00",	--443
		x"4a",	--444
		x"43",	--445
		x"12",	--446
		x"d7",	--447
		x"43",	--448
		x"40",	--449
		x"42",	--450
		x"12",	--451
		x"d4",	--452
		x"4e",	--453
		x"4f",	--454
		x"43",	--455
		x"40",	--456
		x"3f",	--457
		x"12",	--458
		x"d2",	--459
		x"4e",	--460
		x"4f",	--461
		x"42",	--462
		x"02",	--463
		x"12",	--464
		x"c8",	--465
		x"4b",	--466
		x"43",	--467
		x"12",	--468
		x"d7",	--469
		x"43",	--470
		x"40",	--471
		x"42",	--472
		x"12",	--473
		x"d4",	--474
		x"4e",	--475
		x"4f",	--476
		x"42",	--477
		x"02",	--478
		x"12",	--479
		x"c8",	--480
		x"43",	--481
		x"53",	--482
		x"41",	--483
		x"41",	--484
		x"41",	--485
		x"41",	--486
		x"4b",	--487
		x"00",	--488
		x"12",	--489
		x"c7",	--490
		x"43",	--491
		x"4f",	--492
		x"42",	--493
		x"02",	--494
		x"12",	--495
		x"ca",	--496
		x"3f",	--497
		x"43",	--498
		x"40",	--499
		x"c2",	--500
		x"12",	--501
		x"ca",	--502
		x"4f",	--503
		x"02",	--504
		x"3f",	--505
		x"12",	--506
		x"e7",	--507
		x"12",	--508
		x"cd",	--509
		x"40",	--510
		x"e7",	--511
		x"00",	--512
		x"12",	--513
		x"cd",	--514
		x"4b",	--515
		x"00",	--516
		x"12",	--517
		x"e7",	--518
		x"12",	--519
		x"cd",	--520
		x"52",	--521
		x"43",	--522
		x"3f",	--523
		x"12",	--524
		x"12",	--525
		x"42",	--526
		x"02",	--527
		x"12",	--528
		x"cb",	--529
		x"4e",	--530
		x"4f",	--531
		x"42",	--532
		x"02",	--533
		x"12",	--534
		x"cb",	--535
		x"12",	--536
		x"12",	--537
		x"e3",	--538
		x"e3",	--539
		x"53",	--540
		x"63",	--541
		x"12",	--542
		x"12",	--543
		x"12",	--544
		x"e7",	--545
		x"12",	--546
		x"02",	--547
		x"12",	--548
		x"dc",	--549
		x"50",	--550
		x"00",	--551
		x"12",	--552
		x"02",	--553
		x"12",	--554
		x"e7",	--555
		x"12",	--556
		x"cd",	--557
		x"52",	--558
		x"41",	--559
		x"41",	--560
		x"41",	--561
		x"4f",	--562
		x"02",	--563
		x"4e",	--564
		x"02",	--565
		x"41",	--566
		x"4f",	--567
		x"02",	--568
		x"4e",	--569
		x"02",	--570
		x"41",	--571
		x"12",	--572
		x"12",	--573
		x"12",	--574
		x"12",	--575
		x"83",	--576
		x"4f",	--577
		x"4e",	--578
		x"43",	--579
		x"00",	--580
		x"93",	--581
		x"24",	--582
		x"93",	--583
		x"02",	--584
		x"24",	--585
		x"43",	--586
		x"02",	--587
		x"41",	--588
		x"4b",	--589
		x"00",	--590
		x"12",	--591
		x"c7",	--592
		x"4f",	--593
		x"90",	--594
		x"00",	--595
		x"34",	--596
		x"43",	--597
		x"49",	--598
		x"48",	--599
		x"42",	--600
		x"02",	--601
		x"12",	--602
		x"ca",	--603
		x"43",	--604
		x"53",	--605
		x"41",	--606
		x"41",	--607
		x"41",	--608
		x"41",	--609
		x"41",	--610
		x"93",	--611
		x"02",	--612
		x"24",	--613
		x"43",	--614
		x"02",	--615
		x"42",	--616
		x"02",	--617
		x"12",	--618
		x"ca",	--619
		x"43",	--620
		x"53",	--621
		x"41",	--622
		x"41",	--623
		x"41",	--624
		x"41",	--625
		x"41",	--626
		x"41",	--627
		x"4b",	--628
		x"00",	--629
		x"12",	--630
		x"c7",	--631
		x"4f",	--632
		x"90",	--633
		x"00",	--634
		x"3b",	--635
		x"41",	--636
		x"4b",	--637
		x"00",	--638
		x"12",	--639
		x"c7",	--640
		x"4f",	--641
		x"41",	--642
		x"4b",	--643
		x"00",	--644
		x"12",	--645
		x"c7",	--646
		x"4f",	--647
		x"12",	--648
		x"12",	--649
		x"12",	--650
		x"e7",	--651
		x"12",	--652
		x"cd",	--653
		x"50",	--654
		x"00",	--655
		x"4a",	--656
		x"43",	--657
		x"12",	--658
		x"d7",	--659
		x"43",	--660
		x"40",	--661
		x"42",	--662
		x"12",	--663
		x"d4",	--664
		x"4e",	--665
		x"4f",	--666
		x"42",	--667
		x"02",	--668
		x"12",	--669
		x"c8",	--670
		x"4b",	--671
		x"43",	--672
		x"12",	--673
		x"d7",	--674
		x"43",	--675
		x"40",	--676
		x"42",	--677
		x"12",	--678
		x"d4",	--679
		x"4e",	--680
		x"4f",	--681
		x"42",	--682
		x"02",	--683
		x"12",	--684
		x"c8",	--685
		x"3f",	--686
		x"43",	--687
		x"12",	--688
		x"c4",	--689
		x"43",	--690
		x"53",	--691
		x"41",	--692
		x"41",	--693
		x"41",	--694
		x"41",	--695
		x"41",	--696
		x"43",	--697
		x"40",	--698
		x"c4",	--699
		x"12",	--700
		x"ca",	--701
		x"4f",	--702
		x"02",	--703
		x"3f",	--704
		x"43",	--705
		x"93",	--706
		x"02",	--707
		x"24",	--708
		x"43",	--709
		x"4f",	--710
		x"02",	--711
		x"43",	--712
		x"41",	--713
		x"42",	--714
		x"00",	--715
		x"4e",	--716
		x"be",	--717
		x"20",	--718
		x"df",	--719
		x"00",	--720
		x"41",	--721
		x"cf",	--722
		x"00",	--723
		x"41",	--724
		x"42",	--725
		x"02",	--726
		x"92",	--727
		x"2c",	--728
		x"4e",	--729
		x"5f",	--730
		x"4f",	--731
		x"e7",	--732
		x"43",	--733
		x"00",	--734
		x"90",	--735
		x"00",	--736
		x"38",	--737
		x"43",	--738
		x"02",	--739
		x"41",	--740
		x"53",	--741
		x"4e",	--742
		x"02",	--743
		x"41",	--744
		x"40",	--745
		x"00",	--746
		x"00",	--747
		x"3f",	--748
		x"40",	--749
		x"00",	--750
		x"00",	--751
		x"3f",	--752
		x"42",	--753
		x"00",	--754
		x"3f",	--755
		x"40",	--756
		x"00",	--757
		x"00",	--758
		x"3f",	--759
		x"40",	--760
		x"00",	--761
		x"00",	--762
		x"3f",	--763
		x"40",	--764
		x"00",	--765
		x"00",	--766
		x"3f",	--767
		x"40",	--768
		x"00",	--769
		x"00",	--770
		x"3f",	--771
		x"4e",	--772
		x"00",	--773
		x"4d",	--774
		x"00",	--775
		x"4c",	--776
		x"00",	--777
		x"43",	--778
		x"00",	--779
		x"43",	--780
		x"00",	--781
		x"43",	--782
		x"00",	--783
		x"41",	--784
		x"43",	--785
		x"00",	--786
		x"43",	--787
		x"00",	--788
		x"43",	--789
		x"00",	--790
		x"41",	--791
		x"4e",	--792
		x"00",	--793
		x"41",	--794
		x"4e",	--795
		x"00",	--796
		x"41",	--797
		x"4e",	--798
		x"00",	--799
		x"41",	--800
		x"4e",	--801
		x"00",	--802
		x"41",	--803
		x"4f",	--804
		x"00",	--805
		x"8e",	--806
		x"4d",	--807
		x"5f",	--808
		x"00",	--809
		x"4d",	--810
		x"00",	--811
		x"12",	--812
		x"c2",	--813
		x"43",	--814
		x"4e",	--815
		x"01",	--816
		x"4f",	--817
		x"01",	--818
		x"42",	--819
		x"01",	--820
		x"41",	--821
		x"12",	--822
		x"c2",	--823
		x"43",	--824
		x"4d",	--825
		x"01",	--826
		x"4f",	--827
		x"00",	--828
		x"01",	--829
		x"42",	--830
		x"01",	--831
		x"41",	--832
		x"5c",	--833
		x"8f",	--834
		x"00",	--835
		x"12",	--836
		x"c2",	--837
		x"43",	--838
		x"4e",	--839
		x"01",	--840
		x"4f",	--841
		x"00",	--842
		x"01",	--843
		x"42",	--844
		x"01",	--845
		x"41",	--846
		x"5d",	--847
		x"41",	--848
		x"12",	--849
		x"12",	--850
		x"83",	--851
		x"4f",	--852
		x"4e",	--853
		x"12",	--854
		x"e8",	--855
		x"12",	--856
		x"cd",	--857
		x"53",	--858
		x"90",	--859
		x"00",	--860
		x"38",	--861
		x"41",	--862
		x"4b",	--863
		x"00",	--864
		x"12",	--865
		x"c7",	--866
		x"4f",	--867
		x"41",	--868
		x"4b",	--869
		x"00",	--870
		x"12",	--871
		x"c7",	--872
		x"4f",	--873
		x"12",	--874
		x"12",	--875
		x"12",	--876
		x"e8",	--877
		x"12",	--878
		x"cd",	--879
		x"50",	--880
		x"00",	--881
		x"4b",	--882
		x"00",	--883
		x"43",	--884
		x"53",	--885
		x"41",	--886
		x"41",	--887
		x"41",	--888
		x"12",	--889
		x"e8",	--890
		x"12",	--891
		x"cd",	--892
		x"40",	--893
		x"e8",	--894
		x"00",	--895
		x"12",	--896
		x"cd",	--897
		x"4b",	--898
		x"00",	--899
		x"12",	--900
		x"e8",	--901
		x"12",	--902
		x"cd",	--903
		x"52",	--904
		x"43",	--905
		x"3f",	--906
		x"12",	--907
		x"83",	--908
		x"4e",	--909
		x"93",	--910
		x"24",	--911
		x"38",	--912
		x"12",	--913
		x"e8",	--914
		x"12",	--915
		x"cd",	--916
		x"53",	--917
		x"41",	--918
		x"4b",	--919
		x"00",	--920
		x"12",	--921
		x"c7",	--922
		x"12",	--923
		x"12",	--924
		x"12",	--925
		x"e8",	--926
		x"12",	--927
		x"cd",	--928
		x"50",	--929
		x"00",	--930
		x"43",	--931
		x"53",	--932
		x"41",	--933
		x"41",	--934
		x"12",	--935
		x"e8",	--936
		x"12",	--937
		x"cd",	--938
		x"40",	--939
		x"e8",	--940
		x"00",	--941
		x"12",	--942
		x"cd",	--943
		x"4b",	--944
		x"00",	--945
		x"12",	--946
		x"e8",	--947
		x"12",	--948
		x"cd",	--949
		x"52",	--950
		x"43",	--951
		x"3f",	--952
		x"12",	--953
		x"12",	--954
		x"43",	--955
		x"00",	--956
		x"4f",	--957
		x"93",	--958
		x"24",	--959
		x"53",	--960
		x"43",	--961
		x"43",	--962
		x"3c",	--963
		x"90",	--964
		x"00",	--965
		x"2c",	--966
		x"5c",	--967
		x"5c",	--968
		x"5c",	--969
		x"5c",	--970
		x"11",	--971
		x"5d",	--972
		x"50",	--973
		x"ff",	--974
		x"43",	--975
		x"4f",	--976
		x"93",	--977
		x"24",	--978
		x"90",	--979
		x"00",	--980
		x"24",	--981
		x"4d",	--982
		x"50",	--983
		x"ff",	--984
		x"93",	--985
		x"23",	--986
		x"90",	--987
		x"00",	--988
		x"2c",	--989
		x"5c",	--990
		x"4c",	--991
		x"5b",	--992
		x"5b",	--993
		x"5b",	--994
		x"11",	--995
		x"5d",	--996
		x"50",	--997
		x"ff",	--998
		x"4f",	--999
		x"93",	--1000
		x"23",	--1001
		x"43",	--1002
		x"00",	--1003
		x"4c",	--1004
		x"41",	--1005
		x"41",	--1006
		x"41",	--1007
		x"43",	--1008
		x"3f",	--1009
		x"4d",	--1010
		x"50",	--1011
		x"ff",	--1012
		x"90",	--1013
		x"00",	--1014
		x"2c",	--1015
		x"5c",	--1016
		x"5c",	--1017
		x"5c",	--1018
		x"5c",	--1019
		x"11",	--1020
		x"5d",	--1021
		x"50",	--1022
		x"ff",	--1023
		x"43",	--1024
		x"3f",	--1025
		x"4d",	--1026
		x"50",	--1027
		x"ff",	--1028
		x"90",	--1029
		x"00",	--1030
		x"2c",	--1031
		x"5c",	--1032
		x"5c",	--1033
		x"5c",	--1034
		x"5c",	--1035
		x"11",	--1036
		x"5d",	--1037
		x"50",	--1038
		x"ff",	--1039
		x"43",	--1040
		x"3f",	--1041
		x"11",	--1042
		x"12",	--1043
		x"12",	--1044
		x"e8",	--1045
		x"12",	--1046
		x"cd",	--1047
		x"52",	--1048
		x"43",	--1049
		x"4c",	--1050
		x"41",	--1051
		x"41",	--1052
		x"41",	--1053
		x"43",	--1054
		x"3f",	--1055
		x"12",	--1056
		x"12",	--1057
		x"4e",	--1058
		x"4c",	--1059
		x"4e",	--1060
		x"00",	--1061
		x"4d",	--1062
		x"00",	--1063
		x"4c",	--1064
		x"00",	--1065
		x"4d",	--1066
		x"43",	--1067
		x"40",	--1068
		x"36",	--1069
		x"40",	--1070
		x"01",	--1071
		x"12",	--1072
		x"e5",	--1073
		x"4e",	--1074
		x"00",	--1075
		x"12",	--1076
		x"c2",	--1077
		x"43",	--1078
		x"4a",	--1079
		x"01",	--1080
		x"40",	--1081
		x"00",	--1082
		x"01",	--1083
		x"42",	--1084
		x"01",	--1085
		x"00",	--1086
		x"41",	--1087
		x"43",	--1088
		x"41",	--1089
		x"41",	--1090
		x"41",	--1091
		x"12",	--1092
		x"12",	--1093
		x"12",	--1094
		x"43",	--1095
		x"00",	--1096
		x"40",	--1097
		x"3f",	--1098
		x"00",	--1099
		x"4f",	--1100
		x"4b",	--1101
		x"00",	--1102
		x"43",	--1103
		x"12",	--1104
		x"d7",	--1105
		x"43",	--1106
		x"40",	--1107
		x"3f",	--1108
		x"12",	--1109
		x"d2",	--1110
		x"4e",	--1111
		x"4f",	--1112
		x"4b",	--1113
		x"00",	--1114
		x"43",	--1115
		x"12",	--1116
		x"d7",	--1117
		x"4e",	--1118
		x"4f",	--1119
		x"48",	--1120
		x"49",	--1121
		x"12",	--1122
		x"d2",	--1123
		x"12",	--1124
		x"cf",	--1125
		x"4e",	--1126
		x"00",	--1127
		x"43",	--1128
		x"00",	--1129
		x"41",	--1130
		x"41",	--1131
		x"41",	--1132
		x"41",	--1133
		x"12",	--1134
		x"12",	--1135
		x"12",	--1136
		x"4d",	--1137
		x"4e",	--1138
		x"4d",	--1139
		x"00",	--1140
		x"4e",	--1141
		x"00",	--1142
		x"4f",	--1143
		x"49",	--1144
		x"00",	--1145
		x"43",	--1146
		x"12",	--1147
		x"d7",	--1148
		x"4e",	--1149
		x"4f",	--1150
		x"4a",	--1151
		x"4b",	--1152
		x"12",	--1153
		x"d2",	--1154
		x"4e",	--1155
		x"4f",	--1156
		x"49",	--1157
		x"00",	--1158
		x"43",	--1159
		x"12",	--1160
		x"d7",	--1161
		x"4e",	--1162
		x"4f",	--1163
		x"4a",	--1164
		x"4b",	--1165
		x"12",	--1166
		x"d2",	--1167
		x"12",	--1168
		x"cf",	--1169
		x"4e",	--1170
		x"00",	--1171
		x"41",	--1172
		x"41",	--1173
		x"41",	--1174
		x"41",	--1175
		x"4f",	--1176
		x"4e",	--1177
		x"00",	--1178
		x"41",	--1179
		x"12",	--1180
		x"12",	--1181
		x"93",	--1182
		x"02",	--1183
		x"38",	--1184
		x"40",	--1185
		x"02",	--1186
		x"43",	--1187
		x"12",	--1188
		x"4b",	--1189
		x"ff",	--1190
		x"11",	--1191
		x"12",	--1192
		x"12",	--1193
		x"e8",	--1194
		x"12",	--1195
		x"cd",	--1196
		x"50",	--1197
		x"00",	--1198
		x"53",	--1199
		x"50",	--1200
		x"00",	--1201
		x"92",	--1202
		x"02",	--1203
		x"3b",	--1204
		x"43",	--1205
		x"41",	--1206
		x"41",	--1207
		x"41",	--1208
		x"42",	--1209
		x"02",	--1210
		x"90",	--1211
		x"00",	--1212
		x"34",	--1213
		x"4e",	--1214
		x"5f",	--1215
		x"5e",	--1216
		x"5f",	--1217
		x"50",	--1218
		x"02",	--1219
		x"40",	--1220
		x"00",	--1221
		x"00",	--1222
		x"40",	--1223
		x"c9",	--1224
		x"00",	--1225
		x"40",	--1226
		x"02",	--1227
		x"00",	--1228
		x"53",	--1229
		x"4e",	--1230
		x"02",	--1231
		x"41",	--1232
		x"12",	--1233
		x"42",	--1234
		x"02",	--1235
		x"90",	--1236
		x"00",	--1237
		x"34",	--1238
		x"4b",	--1239
		x"5c",	--1240
		x"5b",	--1241
		x"5c",	--1242
		x"50",	--1243
		x"02",	--1244
		x"4f",	--1245
		x"00",	--1246
		x"4e",	--1247
		x"00",	--1248
		x"4d",	--1249
		x"00",	--1250
		x"53",	--1251
		x"4b",	--1252
		x"02",	--1253
		x"43",	--1254
		x"41",	--1255
		x"41",	--1256
		x"43",	--1257
		x"3f",	--1258
		x"12",	--1259
		x"50",	--1260
		x"ff",	--1261
		x"42",	--1262
		x"02",	--1263
		x"93",	--1264
		x"38",	--1265
		x"92",	--1266
		x"02",	--1267
		x"24",	--1268
		x"40",	--1269
		x"02",	--1270
		x"43",	--1271
		x"3c",	--1272
		x"50",	--1273
		x"00",	--1274
		x"9f",	--1275
		x"ff",	--1276
		x"24",	--1277
		x"53",	--1278
		x"9b",	--1279
		x"23",	--1280
		x"12",	--1281
		x"e8",	--1282
		x"12",	--1283
		x"cd",	--1284
		x"53",	--1285
		x"43",	--1286
		x"50",	--1287
		x"00",	--1288
		x"41",	--1289
		x"41",	--1290
		x"43",	--1291
		x"4e",	--1292
		x"00",	--1293
		x"4e",	--1294
		x"93",	--1295
		x"24",	--1296
		x"53",	--1297
		x"43",	--1298
		x"3c",	--1299
		x"4e",	--1300
		x"93",	--1301
		x"24",	--1302
		x"53",	--1303
		x"92",	--1304
		x"34",	--1305
		x"90",	--1306
		x"00",	--1307
		x"23",	--1308
		x"43",	--1309
		x"ff",	--1310
		x"4f",	--1311
		x"5d",	--1312
		x"51",	--1313
		x"4e",	--1314
		x"00",	--1315
		x"53",	--1316
		x"4e",	--1317
		x"93",	--1318
		x"23",	--1319
		x"4c",	--1320
		x"5e",	--1321
		x"5e",	--1322
		x"5c",	--1323
		x"50",	--1324
		x"02",	--1325
		x"41",	--1326
		x"12",	--1327
		x"00",	--1328
		x"50",	--1329
		x"00",	--1330
		x"41",	--1331
		x"41",	--1332
		x"43",	--1333
		x"3f",	--1334
		x"d0",	--1335
		x"02",	--1336
		x"01",	--1337
		x"40",	--1338
		x"0b",	--1339
		x"01",	--1340
		x"43",	--1341
		x"41",	--1342
		x"12",	--1343
		x"4f",	--1344
		x"42",	--1345
		x"02",	--1346
		x"90",	--1347
		x"00",	--1348
		x"34",	--1349
		x"4f",	--1350
		x"5c",	--1351
		x"4c",	--1352
		x"5d",	--1353
		x"5d",	--1354
		x"5d",	--1355
		x"8c",	--1356
		x"50",	--1357
		x"03",	--1358
		x"43",	--1359
		x"00",	--1360
		x"43",	--1361
		x"00",	--1362
		x"43",	--1363
		x"00",	--1364
		x"4b",	--1365
		x"00",	--1366
		x"4e",	--1367
		x"00",	--1368
		x"4f",	--1369
		x"53",	--1370
		x"4e",	--1371
		x"02",	--1372
		x"41",	--1373
		x"41",	--1374
		x"43",	--1375
		x"3f",	--1376
		x"5f",	--1377
		x"4f",	--1378
		x"5c",	--1379
		x"5c",	--1380
		x"5c",	--1381
		x"8f",	--1382
		x"50",	--1383
		x"03",	--1384
		x"43",	--1385
		x"00",	--1386
		x"4e",	--1387
		x"00",	--1388
		x"43",	--1389
		x"00",	--1390
		x"4d",	--1391
		x"00",	--1392
		x"43",	--1393
		x"00",	--1394
		x"43",	--1395
		x"41",	--1396
		x"5f",	--1397
		x"4f",	--1398
		x"5e",	--1399
		x"5e",	--1400
		x"5e",	--1401
		x"8f",	--1402
		x"43",	--1403
		x"03",	--1404
		x"43",	--1405
		x"41",	--1406
		x"12",	--1407
		x"12",	--1408
		x"12",	--1409
		x"12",	--1410
		x"12",	--1411
		x"12",	--1412
		x"12",	--1413
		x"12",	--1414
		x"12",	--1415
		x"93",	--1416
		x"02",	--1417
		x"38",	--1418
		x"40",	--1419
		x"03",	--1420
		x"4a",	--1421
		x"53",	--1422
		x"4a",	--1423
		x"52",	--1424
		x"4a",	--1425
		x"50",	--1426
		x"00",	--1427
		x"43",	--1428
		x"3c",	--1429
		x"53",	--1430
		x"4f",	--1431
		x"00",	--1432
		x"53",	--1433
		x"50",	--1434
		x"00",	--1435
		x"50",	--1436
		x"00",	--1437
		x"50",	--1438
		x"00",	--1439
		x"50",	--1440
		x"00",	--1441
		x"92",	--1442
		x"02",	--1443
		x"34",	--1444
		x"93",	--1445
		x"00",	--1446
		x"27",	--1447
		x"4b",	--1448
		x"9b",	--1449
		x"00",	--1450
		x"2b",	--1451
		x"43",	--1452
		x"00",	--1453
		x"4b",	--1454
		x"00",	--1455
		x"12",	--1456
		x"00",	--1457
		x"93",	--1458
		x"00",	--1459
		x"27",	--1460
		x"47",	--1461
		x"53",	--1462
		x"4f",	--1463
		x"00",	--1464
		x"98",	--1465
		x"2b",	--1466
		x"43",	--1467
		x"00",	--1468
		x"3f",	--1469
		x"f0",	--1470
		x"ff",	--1471
		x"01",	--1472
		x"41",	--1473
		x"41",	--1474
		x"41",	--1475
		x"41",	--1476
		x"41",	--1477
		x"41",	--1478
		x"41",	--1479
		x"41",	--1480
		x"41",	--1481
		x"13",	--1482
		x"4e",	--1483
		x"00",	--1484
		x"43",	--1485
		x"41",	--1486
		x"4f",	--1487
		x"4f",	--1488
		x"4f",	--1489
		x"00",	--1490
		x"41",	--1491
		x"43",	--1492
		x"00",	--1493
		x"41",	--1494
		x"4e",	--1495
		x"00",	--1496
		x"40",	--1497
		x"cb",	--1498
		x"12",	--1499
		x"ca",	--1500
		x"4f",	--1501
		x"02",	--1502
		x"43",	--1503
		x"41",	--1504
		x"4d",	--1505
		x"4f",	--1506
		x"4e",	--1507
		x"00",	--1508
		x"43",	--1509
		x"4c",	--1510
		x"42",	--1511
		x"02",	--1512
		x"12",	--1513
		x"ca",	--1514
		x"41",	--1515
		x"42",	--1516
		x"00",	--1517
		x"f2",	--1518
		x"23",	--1519
		x"4f",	--1520
		x"00",	--1521
		x"43",	--1522
		x"41",	--1523
		x"f0",	--1524
		x"00",	--1525
		x"4f",	--1526
		x"e9",	--1527
		x"11",	--1528
		x"12",	--1529
		x"cb",	--1530
		x"41",	--1531
		x"12",	--1532
		x"4f",	--1533
		x"4f",	--1534
		x"11",	--1535
		x"11",	--1536
		x"11",	--1537
		x"11",	--1538
		x"4e",	--1539
		x"12",	--1540
		x"cb",	--1541
		x"4b",	--1542
		x"12",	--1543
		x"cb",	--1544
		x"41",	--1545
		x"41",	--1546
		x"12",	--1547
		x"12",	--1548
		x"4f",	--1549
		x"40",	--1550
		x"00",	--1551
		x"4a",	--1552
		x"4b",	--1553
		x"f0",	--1554
		x"00",	--1555
		x"24",	--1556
		x"11",	--1557
		x"53",	--1558
		x"23",	--1559
		x"f3",	--1560
		x"24",	--1561
		x"40",	--1562
		x"00",	--1563
		x"12",	--1564
		x"cb",	--1565
		x"53",	--1566
		x"93",	--1567
		x"23",	--1568
		x"41",	--1569
		x"41",	--1570
		x"41",	--1571
		x"40",	--1572
		x"00",	--1573
		x"3f",	--1574
		x"12",	--1575
		x"4f",	--1576
		x"4f",	--1577
		x"10",	--1578
		x"11",	--1579
		x"4e",	--1580
		x"12",	--1581
		x"cb",	--1582
		x"4b",	--1583
		x"12",	--1584
		x"cb",	--1585
		x"41",	--1586
		x"41",	--1587
		x"12",	--1588
		x"12",	--1589
		x"4e",	--1590
		x"4f",	--1591
		x"4f",	--1592
		x"10",	--1593
		x"11",	--1594
		x"4d",	--1595
		x"12",	--1596
		x"cb",	--1597
		x"4b",	--1598
		x"12",	--1599
		x"cb",	--1600
		x"4b",	--1601
		x"4a",	--1602
		x"10",	--1603
		x"10",	--1604
		x"ec",	--1605
		x"ec",	--1606
		x"4d",	--1607
		x"12",	--1608
		x"cb",	--1609
		x"4a",	--1610
		x"12",	--1611
		x"cb",	--1612
		x"41",	--1613
		x"41",	--1614
		x"41",	--1615
		x"12",	--1616
		x"12",	--1617
		x"12",	--1618
		x"4f",	--1619
		x"93",	--1620
		x"24",	--1621
		x"4e",	--1622
		x"53",	--1623
		x"43",	--1624
		x"4a",	--1625
		x"5b",	--1626
		x"4d",	--1627
		x"11",	--1628
		x"12",	--1629
		x"cb",	--1630
		x"99",	--1631
		x"24",	--1632
		x"53",	--1633
		x"b0",	--1634
		x"00",	--1635
		x"20",	--1636
		x"40",	--1637
		x"00",	--1638
		x"12",	--1639
		x"cb",	--1640
		x"3f",	--1641
		x"40",	--1642
		x"00",	--1643
		x"12",	--1644
		x"cb",	--1645
		x"3f",	--1646
		x"41",	--1647
		x"41",	--1648
		x"41",	--1649
		x"41",	--1650
		x"12",	--1651
		x"12",	--1652
		x"12",	--1653
		x"4f",	--1654
		x"93",	--1655
		x"24",	--1656
		x"4e",	--1657
		x"53",	--1658
		x"43",	--1659
		x"4a",	--1660
		x"11",	--1661
		x"12",	--1662
		x"cb",	--1663
		x"99",	--1664
		x"24",	--1665
		x"53",	--1666
		x"b0",	--1667
		x"00",	--1668
		x"23",	--1669
		x"40",	--1670
		x"00",	--1671
		x"12",	--1672
		x"cb",	--1673
		x"4a",	--1674
		x"11",	--1675
		x"12",	--1676
		x"cb",	--1677
		x"99",	--1678
		x"23",	--1679
		x"41",	--1680
		x"41",	--1681
		x"41",	--1682
		x"41",	--1683
		x"12",	--1684
		x"12",	--1685
		x"12",	--1686
		x"50",	--1687
		x"ff",	--1688
		x"4f",	--1689
		x"93",	--1690
		x"38",	--1691
		x"90",	--1692
		x"00",	--1693
		x"38",	--1694
		x"43",	--1695
		x"41",	--1696
		x"59",	--1697
		x"40",	--1698
		x"00",	--1699
		x"4b",	--1700
		x"12",	--1701
		x"e5",	--1702
		x"50",	--1703
		x"00",	--1704
		x"4f",	--1705
		x"00",	--1706
		x"53",	--1707
		x"40",	--1708
		x"00",	--1709
		x"4b",	--1710
		x"12",	--1711
		x"e5",	--1712
		x"4f",	--1713
		x"90",	--1714
		x"00",	--1715
		x"37",	--1716
		x"49",	--1717
		x"53",	--1718
		x"51",	--1719
		x"40",	--1720
		x"00",	--1721
		x"4b",	--1722
		x"12",	--1723
		x"e5",	--1724
		x"50",	--1725
		x"00",	--1726
		x"4f",	--1727
		x"00",	--1728
		x"53",	--1729
		x"41",	--1730
		x"5a",	--1731
		x"4f",	--1732
		x"11",	--1733
		x"12",	--1734
		x"cb",	--1735
		x"93",	--1736
		x"23",	--1737
		x"50",	--1738
		x"00",	--1739
		x"41",	--1740
		x"41",	--1741
		x"41",	--1742
		x"41",	--1743
		x"40",	--1744
		x"00",	--1745
		x"12",	--1746
		x"cb",	--1747
		x"e3",	--1748
		x"53",	--1749
		x"3f",	--1750
		x"43",	--1751
		x"43",	--1752
		x"3f",	--1753
		x"12",	--1754
		x"12",	--1755
		x"12",	--1756
		x"41",	--1757
		x"52",	--1758
		x"4b",	--1759
		x"49",	--1760
		x"93",	--1761
		x"20",	--1762
		x"3c",	--1763
		x"11",	--1764
		x"12",	--1765
		x"cb",	--1766
		x"49",	--1767
		x"4a",	--1768
		x"53",	--1769
		x"4a",	--1770
		x"00",	--1771
		x"93",	--1772
		x"24",	--1773
		x"90",	--1774
		x"00",	--1775
		x"23",	--1776
		x"49",	--1777
		x"53",	--1778
		x"49",	--1779
		x"00",	--1780
		x"50",	--1781
		x"ff",	--1782
		x"90",	--1783
		x"00",	--1784
		x"2f",	--1785
		x"4f",	--1786
		x"5f",	--1787
		x"4f",	--1788
		x"e8",	--1789
		x"41",	--1790
		x"41",	--1791
		x"41",	--1792
		x"41",	--1793
		x"4b",	--1794
		x"52",	--1795
		x"4b",	--1796
		x"00",	--1797
		x"4b",	--1798
		x"12",	--1799
		x"cc",	--1800
		x"49",	--1801
		x"3f",	--1802
		x"4b",	--1803
		x"53",	--1804
		x"4b",	--1805
		x"12",	--1806
		x"cc",	--1807
		x"49",	--1808
		x"3f",	--1809
		x"4b",	--1810
		x"53",	--1811
		x"4f",	--1812
		x"49",	--1813
		x"93",	--1814
		x"27",	--1815
		x"53",	--1816
		x"11",	--1817
		x"12",	--1818
		x"cb",	--1819
		x"49",	--1820
		x"93",	--1821
		x"23",	--1822
		x"3f",	--1823
		x"4b",	--1824
		x"52",	--1825
		x"4b",	--1826
		x"00",	--1827
		x"4b",	--1828
		x"12",	--1829
		x"cc",	--1830
		x"49",	--1831
		x"3f",	--1832
		x"4b",	--1833
		x"53",	--1834
		x"4b",	--1835
		x"4e",	--1836
		x"10",	--1837
		x"11",	--1838
		x"10",	--1839
		x"11",	--1840
		x"12",	--1841
		x"cc",	--1842
		x"49",	--1843
		x"3f",	--1844
		x"4b",	--1845
		x"53",	--1846
		x"4b",	--1847
		x"12",	--1848
		x"cd",	--1849
		x"49",	--1850
		x"3f",	--1851
		x"4b",	--1852
		x"53",	--1853
		x"4b",	--1854
		x"12",	--1855
		x"cb",	--1856
		x"49",	--1857
		x"3f",	--1858
		x"4b",	--1859
		x"53",	--1860
		x"4b",	--1861
		x"12",	--1862
		x"cb",	--1863
		x"49",	--1864
		x"3f",	--1865
		x"4b",	--1866
		x"53",	--1867
		x"4b",	--1868
		x"12",	--1869
		x"cc",	--1870
		x"49",	--1871
		x"3f",	--1872
		x"40",	--1873
		x"00",	--1874
		x"12",	--1875
		x"cb",	--1876
		x"3f",	--1877
		x"12",	--1878
		x"12",	--1879
		x"42",	--1880
		x"02",	--1881
		x"42",	--1882
		x"00",	--1883
		x"04",	--1884
		x"42",	--1885
		x"02",	--1886
		x"90",	--1887
		x"00",	--1888
		x"34",	--1889
		x"53",	--1890
		x"02",	--1891
		x"42",	--1892
		x"02",	--1893
		x"42",	--1894
		x"02",	--1895
		x"9f",	--1896
		x"20",	--1897
		x"53",	--1898
		x"02",	--1899
		x"40",	--1900
		x"00",	--1901
		x"00",	--1902
		x"41",	--1903
		x"41",	--1904
		x"c0",	--1905
		x"00",	--1906
		x"00",	--1907
		x"13",	--1908
		x"43",	--1909
		x"02",	--1910
		x"3f",	--1911
		x"4e",	--1912
		x"4f",	--1913
		x"40",	--1914
		x"36",	--1915
		x"40",	--1916
		x"01",	--1917
		x"12",	--1918
		x"e5",	--1919
		x"53",	--1920
		x"4e",	--1921
		x"00",	--1922
		x"40",	--1923
		x"00",	--1924
		x"00",	--1925
		x"41",	--1926
		x"42",	--1927
		x"02",	--1928
		x"42",	--1929
		x"02",	--1930
		x"9f",	--1931
		x"38",	--1932
		x"42",	--1933
		x"02",	--1934
		x"82",	--1935
		x"02",	--1936
		x"41",	--1937
		x"42",	--1938
		x"02",	--1939
		x"42",	--1940
		x"02",	--1941
		x"40",	--1942
		x"00",	--1943
		x"8d",	--1944
		x"8e",	--1945
		x"41",	--1946
		x"42",	--1947
		x"02",	--1948
		x"4f",	--1949
		x"04",	--1950
		x"42",	--1951
		x"02",	--1952
		x"42",	--1953
		x"02",	--1954
		x"9e",	--1955
		x"24",	--1956
		x"42",	--1957
		x"02",	--1958
		x"90",	--1959
		x"00",	--1960
		x"38",	--1961
		x"43",	--1962
		x"02",	--1963
		x"41",	--1964
		x"53",	--1965
		x"02",	--1966
		x"41",	--1967
		x"43",	--1968
		x"41",	--1969
		x"12",	--1970
		x"12",	--1971
		x"4e",	--1972
		x"4f",	--1973
		x"43",	--1974
		x"40",	--1975
		x"4f",	--1976
		x"12",	--1977
		x"d6",	--1978
		x"93",	--1979
		x"34",	--1980
		x"4a",	--1981
		x"4b",	--1982
		x"12",	--1983
		x"d6",	--1984
		x"41",	--1985
		x"41",	--1986
		x"41",	--1987
		x"43",	--1988
		x"40",	--1989
		x"4f",	--1990
		x"4a",	--1991
		x"4b",	--1992
		x"12",	--1993
		x"d2",	--1994
		x"12",	--1995
		x"d6",	--1996
		x"53",	--1997
		x"60",	--1998
		x"80",	--1999
		x"41",	--2000
		x"41",	--2001
		x"41",	--2002
		x"12",	--2003
		x"12",	--2004
		x"12",	--2005
		x"12",	--2006
		x"12",	--2007
		x"12",	--2008
		x"12",	--2009
		x"12",	--2010
		x"50",	--2011
		x"ff",	--2012
		x"4d",	--2013
		x"4f",	--2014
		x"93",	--2015
		x"28",	--2016
		x"4e",	--2017
		x"93",	--2018
		x"28",	--2019
		x"92",	--2020
		x"20",	--2021
		x"40",	--2022
		x"d2",	--2023
		x"92",	--2024
		x"24",	--2025
		x"93",	--2026
		x"24",	--2027
		x"93",	--2028
		x"24",	--2029
		x"4f",	--2030
		x"00",	--2031
		x"00",	--2032
		x"4e",	--2033
		x"00",	--2034
		x"4f",	--2035
		x"00",	--2036
		x"4f",	--2037
		x"00",	--2038
		x"4e",	--2039
		x"00",	--2040
		x"4e",	--2041
		x"00",	--2042
		x"41",	--2043
		x"8b",	--2044
		x"4c",	--2045
		x"93",	--2046
		x"38",	--2047
		x"90",	--2048
		x"00",	--2049
		x"34",	--2050
		x"93",	--2051
		x"38",	--2052
		x"46",	--2053
		x"00",	--2054
		x"47",	--2055
		x"00",	--2056
		x"49",	--2057
		x"f0",	--2058
		x"00",	--2059
		x"24",	--2060
		x"46",	--2061
		x"47",	--2062
		x"c3",	--2063
		x"10",	--2064
		x"10",	--2065
		x"53",	--2066
		x"23",	--2067
		x"4a",	--2068
		x"00",	--2069
		x"4b",	--2070
		x"00",	--2071
		x"43",	--2072
		x"43",	--2073
		x"f0",	--2074
		x"00",	--2075
		x"24",	--2076
		x"5c",	--2077
		x"6d",	--2078
		x"53",	--2079
		x"23",	--2080
		x"53",	--2081
		x"63",	--2082
		x"f6",	--2083
		x"f7",	--2084
		x"43",	--2085
		x"43",	--2086
		x"93",	--2087
		x"20",	--2088
		x"93",	--2089
		x"24",	--2090
		x"41",	--2091
		x"00",	--2092
		x"41",	--2093
		x"00",	--2094
		x"da",	--2095
		x"db",	--2096
		x"4f",	--2097
		x"00",	--2098
		x"9e",	--2099
		x"00",	--2100
		x"20",	--2101
		x"4f",	--2102
		x"00",	--2103
		x"41",	--2104
		x"00",	--2105
		x"46",	--2106
		x"47",	--2107
		x"54",	--2108
		x"65",	--2109
		x"4e",	--2110
		x"00",	--2111
		x"4f",	--2112
		x"00",	--2113
		x"40",	--2114
		x"00",	--2115
		x"00",	--2116
		x"93",	--2117
		x"38",	--2118
		x"48",	--2119
		x"50",	--2120
		x"00",	--2121
		x"41",	--2122
		x"41",	--2123
		x"41",	--2124
		x"41",	--2125
		x"41",	--2126
		x"41",	--2127
		x"41",	--2128
		x"41",	--2129
		x"41",	--2130
		x"91",	--2131
		x"38",	--2132
		x"4b",	--2133
		x"00",	--2134
		x"43",	--2135
		x"43",	--2136
		x"4f",	--2137
		x"00",	--2138
		x"9e",	--2139
		x"00",	--2140
		x"27",	--2141
		x"93",	--2142
		x"24",	--2143
		x"46",	--2144
		x"47",	--2145
		x"84",	--2146
		x"75",	--2147
		x"93",	--2148
		x"38",	--2149
		x"43",	--2150
		x"00",	--2151
		x"41",	--2152
		x"00",	--2153
		x"4e",	--2154
		x"00",	--2155
		x"4f",	--2156
		x"00",	--2157
		x"4e",	--2158
		x"4f",	--2159
		x"53",	--2160
		x"63",	--2161
		x"90",	--2162
		x"3f",	--2163
		x"28",	--2164
		x"90",	--2165
		x"40",	--2166
		x"2c",	--2167
		x"93",	--2168
		x"2c",	--2169
		x"48",	--2170
		x"00",	--2171
		x"53",	--2172
		x"5e",	--2173
		x"6f",	--2174
		x"4b",	--2175
		x"53",	--2176
		x"4e",	--2177
		x"4f",	--2178
		x"53",	--2179
		x"63",	--2180
		x"90",	--2181
		x"3f",	--2182
		x"2b",	--2183
		x"24",	--2184
		x"4e",	--2185
		x"00",	--2186
		x"4f",	--2187
		x"00",	--2188
		x"4a",	--2189
		x"00",	--2190
		x"40",	--2191
		x"00",	--2192
		x"00",	--2193
		x"93",	--2194
		x"37",	--2195
		x"4e",	--2196
		x"4f",	--2197
		x"f3",	--2198
		x"f3",	--2199
		x"c3",	--2200
		x"10",	--2201
		x"10",	--2202
		x"4c",	--2203
		x"4d",	--2204
		x"de",	--2205
		x"df",	--2206
		x"4a",	--2207
		x"00",	--2208
		x"4b",	--2209
		x"00",	--2210
		x"53",	--2211
		x"00",	--2212
		x"48",	--2213
		x"3f",	--2214
		x"93",	--2215
		x"23",	--2216
		x"4f",	--2217
		x"00",	--2218
		x"4f",	--2219
		x"00",	--2220
		x"00",	--2221
		x"4f",	--2222
		x"00",	--2223
		x"00",	--2224
		x"4f",	--2225
		x"00",	--2226
		x"00",	--2227
		x"4e",	--2228
		x"00",	--2229
		x"ff",	--2230
		x"00",	--2231
		x"4e",	--2232
		x"00",	--2233
		x"4d",	--2234
		x"3f",	--2235
		x"43",	--2236
		x"43",	--2237
		x"3f",	--2238
		x"e3",	--2239
		x"53",	--2240
		x"90",	--2241
		x"00",	--2242
		x"37",	--2243
		x"3f",	--2244
		x"93",	--2245
		x"2b",	--2246
		x"3f",	--2247
		x"44",	--2248
		x"45",	--2249
		x"86",	--2250
		x"77",	--2251
		x"3f",	--2252
		x"4e",	--2253
		x"3f",	--2254
		x"43",	--2255
		x"00",	--2256
		x"41",	--2257
		x"00",	--2258
		x"e3",	--2259
		x"e3",	--2260
		x"53",	--2261
		x"63",	--2262
		x"4e",	--2263
		x"00",	--2264
		x"4f",	--2265
		x"00",	--2266
		x"3f",	--2267
		x"93",	--2268
		x"27",	--2269
		x"59",	--2270
		x"00",	--2271
		x"44",	--2272
		x"00",	--2273
		x"45",	--2274
		x"00",	--2275
		x"49",	--2276
		x"f0",	--2277
		x"00",	--2278
		x"24",	--2279
		x"4d",	--2280
		x"44",	--2281
		x"45",	--2282
		x"c3",	--2283
		x"10",	--2284
		x"10",	--2285
		x"53",	--2286
		x"23",	--2287
		x"4c",	--2288
		x"00",	--2289
		x"4d",	--2290
		x"00",	--2291
		x"43",	--2292
		x"43",	--2293
		x"f0",	--2294
		x"00",	--2295
		x"24",	--2296
		x"5c",	--2297
		x"6d",	--2298
		x"53",	--2299
		x"23",	--2300
		x"53",	--2301
		x"63",	--2302
		x"f4",	--2303
		x"f5",	--2304
		x"43",	--2305
		x"43",	--2306
		x"93",	--2307
		x"20",	--2308
		x"93",	--2309
		x"20",	--2310
		x"43",	--2311
		x"43",	--2312
		x"41",	--2313
		x"00",	--2314
		x"41",	--2315
		x"00",	--2316
		x"da",	--2317
		x"db",	--2318
		x"3f",	--2319
		x"43",	--2320
		x"43",	--2321
		x"3f",	--2322
		x"92",	--2323
		x"23",	--2324
		x"9e",	--2325
		x"00",	--2326
		x"00",	--2327
		x"27",	--2328
		x"40",	--2329
		x"e9",	--2330
		x"3f",	--2331
		x"50",	--2332
		x"ff",	--2333
		x"4e",	--2334
		x"00",	--2335
		x"4f",	--2336
		x"00",	--2337
		x"4c",	--2338
		x"00",	--2339
		x"4d",	--2340
		x"00",	--2341
		x"41",	--2342
		x"50",	--2343
		x"00",	--2344
		x"41",	--2345
		x"52",	--2346
		x"12",	--2347
		x"da",	--2348
		x"41",	--2349
		x"50",	--2350
		x"00",	--2351
		x"41",	--2352
		x"12",	--2353
		x"da",	--2354
		x"41",	--2355
		x"52",	--2356
		x"41",	--2357
		x"50",	--2358
		x"00",	--2359
		x"41",	--2360
		x"50",	--2361
		x"00",	--2362
		x"12",	--2363
		x"cf",	--2364
		x"12",	--2365
		x"d8",	--2366
		x"50",	--2367
		x"00",	--2368
		x"41",	--2369
		x"50",	--2370
		x"ff",	--2371
		x"4e",	--2372
		x"00",	--2373
		x"4f",	--2374
		x"00",	--2375
		x"4c",	--2376
		x"00",	--2377
		x"4d",	--2378
		x"00",	--2379
		x"41",	--2380
		x"50",	--2381
		x"00",	--2382
		x"41",	--2383
		x"52",	--2384
		x"12",	--2385
		x"da",	--2386
		x"41",	--2387
		x"50",	--2388
		x"00",	--2389
		x"41",	--2390
		x"12",	--2391
		x"da",	--2392
		x"e3",	--2393
		x"00",	--2394
		x"41",	--2395
		x"52",	--2396
		x"41",	--2397
		x"50",	--2398
		x"00",	--2399
		x"41",	--2400
		x"50",	--2401
		x"00",	--2402
		x"12",	--2403
		x"cf",	--2404
		x"12",	--2405
		x"d8",	--2406
		x"50",	--2407
		x"00",	--2408
		x"41",	--2409
		x"12",	--2410
		x"12",	--2411
		x"12",	--2412
		x"12",	--2413
		x"12",	--2414
		x"12",	--2415
		x"12",	--2416
		x"12",	--2417
		x"50",	--2418
		x"ff",	--2419
		x"4e",	--2420
		x"00",	--2421
		x"4f",	--2422
		x"00",	--2423
		x"4c",	--2424
		x"00",	--2425
		x"4d",	--2426
		x"00",	--2427
		x"41",	--2428
		x"50",	--2429
		x"00",	--2430
		x"41",	--2431
		x"52",	--2432
		x"12",	--2433
		x"da",	--2434
		x"41",	--2435
		x"50",	--2436
		x"00",	--2437
		x"41",	--2438
		x"12",	--2439
		x"da",	--2440
		x"41",	--2441
		x"00",	--2442
		x"93",	--2443
		x"28",	--2444
		x"41",	--2445
		x"00",	--2446
		x"93",	--2447
		x"28",	--2448
		x"92",	--2449
		x"24",	--2450
		x"92",	--2451
		x"24",	--2452
		x"93",	--2453
		x"24",	--2454
		x"93",	--2455
		x"24",	--2456
		x"41",	--2457
		x"00",	--2458
		x"41",	--2459
		x"00",	--2460
		x"41",	--2461
		x"00",	--2462
		x"41",	--2463
		x"00",	--2464
		x"40",	--2465
		x"00",	--2466
		x"43",	--2467
		x"43",	--2468
		x"43",	--2469
		x"43",	--2470
		x"43",	--2471
		x"00",	--2472
		x"43",	--2473
		x"00",	--2474
		x"43",	--2475
		x"43",	--2476
		x"4c",	--2477
		x"00",	--2478
		x"3c",	--2479
		x"58",	--2480
		x"69",	--2481
		x"c3",	--2482
		x"10",	--2483
		x"10",	--2484
		x"53",	--2485
		x"00",	--2486
		x"24",	--2487
		x"b3",	--2488
		x"24",	--2489
		x"58",	--2490
		x"69",	--2491
		x"56",	--2492
		x"67",	--2493
		x"43",	--2494
		x"43",	--2495
		x"99",	--2496
		x"28",	--2497
		x"24",	--2498
		x"43",	--2499
		x"43",	--2500
		x"5c",	--2501
		x"6d",	--2502
		x"56",	--2503
		x"67",	--2504
		x"93",	--2505
		x"37",	--2506
		x"d3",	--2507
		x"d3",	--2508
		x"3f",	--2509
		x"98",	--2510
		x"2b",	--2511
		x"3f",	--2512
		x"4a",	--2513
		x"00",	--2514
		x"4b",	--2515
		x"00",	--2516
		x"4f",	--2517
		x"41",	--2518
		x"00",	--2519
		x"51",	--2520
		x"00",	--2521
		x"4a",	--2522
		x"53",	--2523
		x"46",	--2524
		x"00",	--2525
		x"43",	--2526
		x"91",	--2527
		x"00",	--2528
		x"00",	--2529
		x"24",	--2530
		x"4d",	--2531
		x"00",	--2532
		x"93",	--2533
		x"38",	--2534
		x"90",	--2535
		x"40",	--2536
		x"2c",	--2537
		x"41",	--2538
		x"00",	--2539
		x"53",	--2540
		x"41",	--2541
		x"00",	--2542
		x"41",	--2543
		x"00",	--2544
		x"4d",	--2545
		x"5e",	--2546
		x"6f",	--2547
		x"93",	--2548
		x"38",	--2549
		x"5a",	--2550
		x"6b",	--2551
		x"53",	--2552
		x"90",	--2553
		x"40",	--2554
		x"2b",	--2555
		x"4a",	--2556
		x"00",	--2557
		x"4b",	--2558
		x"00",	--2559
		x"4c",	--2560
		x"00",	--2561
		x"4e",	--2562
		x"4f",	--2563
		x"f0",	--2564
		x"00",	--2565
		x"f3",	--2566
		x"90",	--2567
		x"00",	--2568
		x"24",	--2569
		x"4e",	--2570
		x"00",	--2571
		x"4f",	--2572
		x"00",	--2573
		x"40",	--2574
		x"00",	--2575
		x"00",	--2576
		x"41",	--2577
		x"52",	--2578
		x"12",	--2579
		x"d8",	--2580
		x"50",	--2581
		x"00",	--2582
		x"41",	--2583
		x"41",	--2584
		x"41",	--2585
		x"41",	--2586
		x"41",	--2587
		x"41",	--2588
		x"41",	--2589
		x"41",	--2590
		x"41",	--2591
		x"d3",	--2592
		x"d3",	--2593
		x"3f",	--2594
		x"50",	--2595
		x"00",	--2596
		x"4a",	--2597
		x"b3",	--2598
		x"24",	--2599
		x"41",	--2600
		x"00",	--2601
		x"41",	--2602
		x"00",	--2603
		x"c3",	--2604
		x"10",	--2605
		x"10",	--2606
		x"4c",	--2607
		x"4d",	--2608
		x"d3",	--2609
		x"d0",	--2610
		x"80",	--2611
		x"46",	--2612
		x"00",	--2613
		x"47",	--2614
		x"00",	--2615
		x"c3",	--2616
		x"10",	--2617
		x"10",	--2618
		x"53",	--2619
		x"93",	--2620
		x"3b",	--2621
		x"48",	--2622
		x"00",	--2623
		x"3f",	--2624
		x"93",	--2625
		x"24",	--2626
		x"43",	--2627
		x"91",	--2628
		x"00",	--2629
		x"00",	--2630
		x"24",	--2631
		x"4f",	--2632
		x"00",	--2633
		x"41",	--2634
		x"50",	--2635
		x"00",	--2636
		x"3f",	--2637
		x"93",	--2638
		x"23",	--2639
		x"4e",	--2640
		x"4f",	--2641
		x"f0",	--2642
		x"00",	--2643
		x"f3",	--2644
		x"93",	--2645
		x"23",	--2646
		x"93",	--2647
		x"23",	--2648
		x"93",	--2649
		x"00",	--2650
		x"20",	--2651
		x"93",	--2652
		x"00",	--2653
		x"27",	--2654
		x"50",	--2655
		x"00",	--2656
		x"63",	--2657
		x"f0",	--2658
		x"ff",	--2659
		x"f3",	--2660
		x"3f",	--2661
		x"43",	--2662
		x"3f",	--2663
		x"43",	--2664
		x"3f",	--2665
		x"43",	--2666
		x"91",	--2667
		x"00",	--2668
		x"00",	--2669
		x"24",	--2670
		x"4f",	--2671
		x"00",	--2672
		x"41",	--2673
		x"50",	--2674
		x"00",	--2675
		x"3f",	--2676
		x"43",	--2677
		x"3f",	--2678
		x"93",	--2679
		x"23",	--2680
		x"40",	--2681
		x"e9",	--2682
		x"3f",	--2683
		x"12",	--2684
		x"12",	--2685
		x"12",	--2686
		x"12",	--2687
		x"12",	--2688
		x"50",	--2689
		x"ff",	--2690
		x"4e",	--2691
		x"00",	--2692
		x"4f",	--2693
		x"00",	--2694
		x"4c",	--2695
		x"00",	--2696
		x"4d",	--2697
		x"00",	--2698
		x"41",	--2699
		x"50",	--2700
		x"00",	--2701
		x"41",	--2702
		x"52",	--2703
		x"12",	--2704
		x"da",	--2705
		x"41",	--2706
		x"52",	--2707
		x"41",	--2708
		x"12",	--2709
		x"da",	--2710
		x"41",	--2711
		x"00",	--2712
		x"93",	--2713
		x"28",	--2714
		x"41",	--2715
		x"00",	--2716
		x"93",	--2717
		x"28",	--2718
		x"e1",	--2719
		x"00",	--2720
		x"00",	--2721
		x"92",	--2722
		x"24",	--2723
		x"93",	--2724
		x"24",	--2725
		x"92",	--2726
		x"24",	--2727
		x"93",	--2728
		x"24",	--2729
		x"41",	--2730
		x"00",	--2731
		x"81",	--2732
		x"00",	--2733
		x"4d",	--2734
		x"00",	--2735
		x"41",	--2736
		x"00",	--2737
		x"41",	--2738
		x"00",	--2739
		x"41",	--2740
		x"00",	--2741
		x"41",	--2742
		x"00",	--2743
		x"99",	--2744
		x"2c",	--2745
		x"5e",	--2746
		x"6f",	--2747
		x"53",	--2748
		x"4d",	--2749
		x"00",	--2750
		x"40",	--2751
		x"00",	--2752
		x"43",	--2753
		x"40",	--2754
		x"40",	--2755
		x"43",	--2756
		x"43",	--2757
		x"3c",	--2758
		x"dc",	--2759
		x"dd",	--2760
		x"88",	--2761
		x"79",	--2762
		x"c3",	--2763
		x"10",	--2764
		x"10",	--2765
		x"5e",	--2766
		x"6f",	--2767
		x"53",	--2768
		x"24",	--2769
		x"99",	--2770
		x"2b",	--2771
		x"23",	--2772
		x"98",	--2773
		x"2b",	--2774
		x"3f",	--2775
		x"9f",	--2776
		x"2b",	--2777
		x"98",	--2778
		x"2f",	--2779
		x"3f",	--2780
		x"4a",	--2781
		x"4b",	--2782
		x"f0",	--2783
		x"00",	--2784
		x"f3",	--2785
		x"90",	--2786
		x"00",	--2787
		x"24",	--2788
		x"4a",	--2789
		x"00",	--2790
		x"4b",	--2791
		x"00",	--2792
		x"41",	--2793
		x"50",	--2794
		x"00",	--2795
		x"12",	--2796
		x"d8",	--2797
		x"50",	--2798
		x"00",	--2799
		x"41",	--2800
		x"41",	--2801
		x"41",	--2802
		x"41",	--2803
		x"41",	--2804
		x"41",	--2805
		x"42",	--2806
		x"00",	--2807
		x"41",	--2808
		x"50",	--2809
		x"00",	--2810
		x"3f",	--2811
		x"9e",	--2812
		x"23",	--2813
		x"40",	--2814
		x"e9",	--2815
		x"3f",	--2816
		x"93",	--2817
		x"23",	--2818
		x"4a",	--2819
		x"4b",	--2820
		x"f0",	--2821
		x"00",	--2822
		x"f3",	--2823
		x"93",	--2824
		x"23",	--2825
		x"93",	--2826
		x"23",	--2827
		x"93",	--2828
		x"20",	--2829
		x"93",	--2830
		x"27",	--2831
		x"50",	--2832
		x"00",	--2833
		x"63",	--2834
		x"f0",	--2835
		x"ff",	--2836
		x"f3",	--2837
		x"3f",	--2838
		x"43",	--2839
		x"00",	--2840
		x"43",	--2841
		x"00",	--2842
		x"43",	--2843
		x"00",	--2844
		x"41",	--2845
		x"50",	--2846
		x"00",	--2847
		x"3f",	--2848
		x"41",	--2849
		x"52",	--2850
		x"3f",	--2851
		x"50",	--2852
		x"ff",	--2853
		x"4e",	--2854
		x"00",	--2855
		x"4f",	--2856
		x"00",	--2857
		x"4c",	--2858
		x"00",	--2859
		x"4d",	--2860
		x"00",	--2861
		x"41",	--2862
		x"50",	--2863
		x"00",	--2864
		x"41",	--2865
		x"52",	--2866
		x"12",	--2867
		x"da",	--2868
		x"41",	--2869
		x"52",	--2870
		x"41",	--2871
		x"12",	--2872
		x"da",	--2873
		x"93",	--2874
		x"00",	--2875
		x"28",	--2876
		x"93",	--2877
		x"00",	--2878
		x"28",	--2879
		x"41",	--2880
		x"52",	--2881
		x"41",	--2882
		x"50",	--2883
		x"00",	--2884
		x"12",	--2885
		x"db",	--2886
		x"50",	--2887
		x"00",	--2888
		x"41",	--2889
		x"43",	--2890
		x"3f",	--2891
		x"50",	--2892
		x"ff",	--2893
		x"4e",	--2894
		x"00",	--2895
		x"4f",	--2896
		x"00",	--2897
		x"41",	--2898
		x"52",	--2899
		x"41",	--2900
		x"12",	--2901
		x"da",	--2902
		x"41",	--2903
		x"00",	--2904
		x"93",	--2905
		x"24",	--2906
		x"28",	--2907
		x"92",	--2908
		x"24",	--2909
		x"41",	--2910
		x"00",	--2911
		x"93",	--2912
		x"38",	--2913
		x"90",	--2914
		x"00",	--2915
		x"38",	--2916
		x"93",	--2917
		x"00",	--2918
		x"20",	--2919
		x"43",	--2920
		x"40",	--2921
		x"7f",	--2922
		x"50",	--2923
		x"00",	--2924
		x"41",	--2925
		x"41",	--2926
		x"00",	--2927
		x"41",	--2928
		x"00",	--2929
		x"40",	--2930
		x"00",	--2931
		x"8d",	--2932
		x"4c",	--2933
		x"f0",	--2934
		x"00",	--2935
		x"20",	--2936
		x"93",	--2937
		x"00",	--2938
		x"27",	--2939
		x"e3",	--2940
		x"e3",	--2941
		x"53",	--2942
		x"63",	--2943
		x"50",	--2944
		x"00",	--2945
		x"41",	--2946
		x"43",	--2947
		x"43",	--2948
		x"50",	--2949
		x"00",	--2950
		x"41",	--2951
		x"c3",	--2952
		x"10",	--2953
		x"10",	--2954
		x"53",	--2955
		x"23",	--2956
		x"3f",	--2957
		x"43",	--2958
		x"40",	--2959
		x"80",	--2960
		x"50",	--2961
		x"00",	--2962
		x"41",	--2963
		x"12",	--2964
		x"12",	--2965
		x"12",	--2966
		x"12",	--2967
		x"82",	--2968
		x"4e",	--2969
		x"4f",	--2970
		x"43",	--2971
		x"00",	--2972
		x"93",	--2973
		x"20",	--2974
		x"93",	--2975
		x"20",	--2976
		x"43",	--2977
		x"00",	--2978
		x"41",	--2979
		x"12",	--2980
		x"d8",	--2981
		x"52",	--2982
		x"41",	--2983
		x"41",	--2984
		x"41",	--2985
		x"41",	--2986
		x"41",	--2987
		x"40",	--2988
		x"00",	--2989
		x"00",	--2990
		x"40",	--2991
		x"00",	--2992
		x"00",	--2993
		x"4a",	--2994
		x"00",	--2995
		x"4b",	--2996
		x"00",	--2997
		x"4a",	--2998
		x"4b",	--2999
		x"12",	--3000
		x"d8",	--3001
		x"53",	--3002
		x"93",	--3003
		x"38",	--3004
		x"27",	--3005
		x"4a",	--3006
		x"00",	--3007
		x"4b",	--3008
		x"00",	--3009
		x"4f",	--3010
		x"f0",	--3011
		x"00",	--3012
		x"20",	--3013
		x"40",	--3014
		x"00",	--3015
		x"8f",	--3016
		x"4e",	--3017
		x"00",	--3018
		x"3f",	--3019
		x"51",	--3020
		x"00",	--3021
		x"00",	--3022
		x"61",	--3023
		x"00",	--3024
		x"00",	--3025
		x"53",	--3026
		x"23",	--3027
		x"3f",	--3028
		x"4f",	--3029
		x"e3",	--3030
		x"53",	--3031
		x"43",	--3032
		x"43",	--3033
		x"4e",	--3034
		x"f0",	--3035
		x"00",	--3036
		x"24",	--3037
		x"5c",	--3038
		x"6d",	--3039
		x"53",	--3040
		x"23",	--3041
		x"53",	--3042
		x"63",	--3043
		x"fa",	--3044
		x"fb",	--3045
		x"43",	--3046
		x"43",	--3047
		x"93",	--3048
		x"20",	--3049
		x"93",	--3050
		x"20",	--3051
		x"43",	--3052
		x"43",	--3053
		x"f0",	--3054
		x"00",	--3055
		x"20",	--3056
		x"48",	--3057
		x"49",	--3058
		x"da",	--3059
		x"db",	--3060
		x"4d",	--3061
		x"00",	--3062
		x"4e",	--3063
		x"00",	--3064
		x"40",	--3065
		x"00",	--3066
		x"8f",	--3067
		x"4e",	--3068
		x"00",	--3069
		x"3f",	--3070
		x"c3",	--3071
		x"10",	--3072
		x"10",	--3073
		x"53",	--3074
		x"23",	--3075
		x"3f",	--3076
		x"12",	--3077
		x"12",	--3078
		x"12",	--3079
		x"93",	--3080
		x"2c",	--3081
		x"90",	--3082
		x"01",	--3083
		x"28",	--3084
		x"40",	--3085
		x"00",	--3086
		x"43",	--3087
		x"42",	--3088
		x"4e",	--3089
		x"4f",	--3090
		x"49",	--3091
		x"93",	--3092
		x"20",	--3093
		x"50",	--3094
		x"e9",	--3095
		x"4c",	--3096
		x"43",	--3097
		x"8e",	--3098
		x"7f",	--3099
		x"4a",	--3100
		x"41",	--3101
		x"41",	--3102
		x"41",	--3103
		x"41",	--3104
		x"90",	--3105
		x"01",	--3106
		x"28",	--3107
		x"42",	--3108
		x"43",	--3109
		x"40",	--3110
		x"00",	--3111
		x"4e",	--3112
		x"4f",	--3113
		x"49",	--3114
		x"93",	--3115
		x"27",	--3116
		x"c3",	--3117
		x"10",	--3118
		x"10",	--3119
		x"53",	--3120
		x"23",	--3121
		x"3f",	--3122
		x"40",	--3123
		x"00",	--3124
		x"43",	--3125
		x"40",	--3126
		x"00",	--3127
		x"3f",	--3128
		x"40",	--3129
		x"00",	--3130
		x"43",	--3131
		x"43",	--3132
		x"3f",	--3133
		x"12",	--3134
		x"12",	--3135
		x"12",	--3136
		x"12",	--3137
		x"12",	--3138
		x"4f",	--3139
		x"4f",	--3140
		x"00",	--3141
		x"4f",	--3142
		x"00",	--3143
		x"4d",	--3144
		x"00",	--3145
		x"4d",	--3146
		x"93",	--3147
		x"28",	--3148
		x"92",	--3149
		x"24",	--3150
		x"93",	--3151
		x"24",	--3152
		x"93",	--3153
		x"24",	--3154
		x"4d",	--3155
		x"00",	--3156
		x"90",	--3157
		x"ff",	--3158
		x"38",	--3159
		x"90",	--3160
		x"00",	--3161
		x"34",	--3162
		x"4e",	--3163
		x"4f",	--3164
		x"f0",	--3165
		x"00",	--3166
		x"f3",	--3167
		x"90",	--3168
		x"00",	--3169
		x"24",	--3170
		x"50",	--3171
		x"00",	--3172
		x"63",	--3173
		x"93",	--3174
		x"38",	--3175
		x"4b",	--3176
		x"50",	--3177
		x"00",	--3178
		x"c3",	--3179
		x"10",	--3180
		x"10",	--3181
		x"c3",	--3182
		x"10",	--3183
		x"10",	--3184
		x"c3",	--3185
		x"10",	--3186
		x"10",	--3187
		x"c3",	--3188
		x"10",	--3189
		x"10",	--3190
		x"c3",	--3191
		x"10",	--3192
		x"10",	--3193
		x"c3",	--3194
		x"10",	--3195
		x"10",	--3196
		x"c3",	--3197
		x"10",	--3198
		x"10",	--3199
		x"f3",	--3200
		x"f0",	--3201
		x"00",	--3202
		x"4d",	--3203
		x"3c",	--3204
		x"93",	--3205
		x"23",	--3206
		x"43",	--3207
		x"43",	--3208
		x"43",	--3209
		x"4d",	--3210
		x"5d",	--3211
		x"5d",	--3212
		x"5d",	--3213
		x"5d",	--3214
		x"5d",	--3215
		x"5d",	--3216
		x"5d",	--3217
		x"4f",	--3218
		x"f0",	--3219
		x"00",	--3220
		x"dd",	--3221
		x"4a",	--3222
		x"11",	--3223
		x"43",	--3224
		x"10",	--3225
		x"4c",	--3226
		x"df",	--3227
		x"4d",	--3228
		x"41",	--3229
		x"41",	--3230
		x"41",	--3231
		x"41",	--3232
		x"41",	--3233
		x"41",	--3234
		x"93",	--3235
		x"23",	--3236
		x"4e",	--3237
		x"4f",	--3238
		x"f0",	--3239
		x"00",	--3240
		x"f3",	--3241
		x"93",	--3242
		x"20",	--3243
		x"93",	--3244
		x"27",	--3245
		x"50",	--3246
		x"00",	--3247
		x"63",	--3248
		x"3f",	--3249
		x"c3",	--3250
		x"10",	--3251
		x"10",	--3252
		x"4b",	--3253
		x"50",	--3254
		x"00",	--3255
		x"3f",	--3256
		x"43",	--3257
		x"43",	--3258
		x"43",	--3259
		x"3f",	--3260
		x"d3",	--3261
		x"d0",	--3262
		x"00",	--3263
		x"f3",	--3264
		x"f0",	--3265
		x"00",	--3266
		x"43",	--3267
		x"3f",	--3268
		x"40",	--3269
		x"ff",	--3270
		x"8b",	--3271
		x"90",	--3272
		x"00",	--3273
		x"34",	--3274
		x"4e",	--3275
		x"4f",	--3276
		x"47",	--3277
		x"f0",	--3278
		x"00",	--3279
		x"24",	--3280
		x"c3",	--3281
		x"10",	--3282
		x"10",	--3283
		x"53",	--3284
		x"23",	--3285
		x"43",	--3286
		x"43",	--3287
		x"f0",	--3288
		x"00",	--3289
		x"24",	--3290
		x"58",	--3291
		x"69",	--3292
		x"53",	--3293
		x"23",	--3294
		x"53",	--3295
		x"63",	--3296
		x"fe",	--3297
		x"ff",	--3298
		x"43",	--3299
		x"43",	--3300
		x"93",	--3301
		x"20",	--3302
		x"93",	--3303
		x"20",	--3304
		x"43",	--3305
		x"43",	--3306
		x"4e",	--3307
		x"4f",	--3308
		x"dc",	--3309
		x"dd",	--3310
		x"48",	--3311
		x"49",	--3312
		x"f0",	--3313
		x"00",	--3314
		x"f3",	--3315
		x"90",	--3316
		x"00",	--3317
		x"24",	--3318
		x"50",	--3319
		x"00",	--3320
		x"63",	--3321
		x"48",	--3322
		x"49",	--3323
		x"c3",	--3324
		x"10",	--3325
		x"10",	--3326
		x"c3",	--3327
		x"10",	--3328
		x"10",	--3329
		x"c3",	--3330
		x"10",	--3331
		x"10",	--3332
		x"c3",	--3333
		x"10",	--3334
		x"10",	--3335
		x"c3",	--3336
		x"10",	--3337
		x"10",	--3338
		x"c3",	--3339
		x"10",	--3340
		x"10",	--3341
		x"c3",	--3342
		x"10",	--3343
		x"10",	--3344
		x"f3",	--3345
		x"f0",	--3346
		x"00",	--3347
		x"43",	--3348
		x"90",	--3349
		x"40",	--3350
		x"2f",	--3351
		x"43",	--3352
		x"3f",	--3353
		x"43",	--3354
		x"43",	--3355
		x"3f",	--3356
		x"93",	--3357
		x"23",	--3358
		x"48",	--3359
		x"49",	--3360
		x"f0",	--3361
		x"00",	--3362
		x"f3",	--3363
		x"93",	--3364
		x"24",	--3365
		x"50",	--3366
		x"00",	--3367
		x"63",	--3368
		x"3f",	--3369
		x"93",	--3370
		x"27",	--3371
		x"3f",	--3372
		x"12",	--3373
		x"12",	--3374
		x"4f",	--3375
		x"4f",	--3376
		x"00",	--3377
		x"f0",	--3378
		x"00",	--3379
		x"4f",	--3380
		x"00",	--3381
		x"c3",	--3382
		x"10",	--3383
		x"c3",	--3384
		x"10",	--3385
		x"c3",	--3386
		x"10",	--3387
		x"c3",	--3388
		x"10",	--3389
		x"c3",	--3390
		x"10",	--3391
		x"c3",	--3392
		x"10",	--3393
		x"c3",	--3394
		x"10",	--3395
		x"4d",	--3396
		x"4f",	--3397
		x"00",	--3398
		x"b0",	--3399
		x"00",	--3400
		x"43",	--3401
		x"6f",	--3402
		x"4f",	--3403
		x"00",	--3404
		x"93",	--3405
		x"20",	--3406
		x"93",	--3407
		x"24",	--3408
		x"40",	--3409
		x"ff",	--3410
		x"00",	--3411
		x"4a",	--3412
		x"4b",	--3413
		x"5c",	--3414
		x"6d",	--3415
		x"5c",	--3416
		x"6d",	--3417
		x"5c",	--3418
		x"6d",	--3419
		x"5c",	--3420
		x"6d",	--3421
		x"5c",	--3422
		x"6d",	--3423
		x"5c",	--3424
		x"6d",	--3425
		x"5c",	--3426
		x"6d",	--3427
		x"40",	--3428
		x"00",	--3429
		x"00",	--3430
		x"90",	--3431
		x"40",	--3432
		x"2c",	--3433
		x"40",	--3434
		x"ff",	--3435
		x"5c",	--3436
		x"6d",	--3437
		x"4f",	--3438
		x"53",	--3439
		x"90",	--3440
		x"40",	--3441
		x"2b",	--3442
		x"4a",	--3443
		x"00",	--3444
		x"4c",	--3445
		x"00",	--3446
		x"4d",	--3447
		x"00",	--3448
		x"41",	--3449
		x"41",	--3450
		x"41",	--3451
		x"90",	--3452
		x"00",	--3453
		x"24",	--3454
		x"50",	--3455
		x"ff",	--3456
		x"4d",	--3457
		x"00",	--3458
		x"40",	--3459
		x"00",	--3460
		x"00",	--3461
		x"4a",	--3462
		x"4b",	--3463
		x"5c",	--3464
		x"6d",	--3465
		x"5c",	--3466
		x"6d",	--3467
		x"5c",	--3468
		x"6d",	--3469
		x"5c",	--3470
		x"6d",	--3471
		x"5c",	--3472
		x"6d",	--3473
		x"5c",	--3474
		x"6d",	--3475
		x"5c",	--3476
		x"6d",	--3477
		x"4c",	--3478
		x"4d",	--3479
		x"d3",	--3480
		x"d0",	--3481
		x"40",	--3482
		x"4a",	--3483
		x"00",	--3484
		x"4b",	--3485
		x"00",	--3486
		x"41",	--3487
		x"41",	--3488
		x"41",	--3489
		x"93",	--3490
		x"23",	--3491
		x"43",	--3492
		x"00",	--3493
		x"41",	--3494
		x"41",	--3495
		x"41",	--3496
		x"93",	--3497
		x"24",	--3498
		x"4a",	--3499
		x"4b",	--3500
		x"f3",	--3501
		x"f0",	--3502
		x"00",	--3503
		x"93",	--3504
		x"20",	--3505
		x"93",	--3506
		x"24",	--3507
		x"43",	--3508
		x"00",	--3509
		x"3f",	--3510
		x"93",	--3511
		x"23",	--3512
		x"42",	--3513
		x"00",	--3514
		x"3f",	--3515
		x"43",	--3516
		x"00",	--3517
		x"3f",	--3518
		x"12",	--3519
		x"4f",	--3520
		x"93",	--3521
		x"28",	--3522
		x"4e",	--3523
		x"93",	--3524
		x"28",	--3525
		x"92",	--3526
		x"24",	--3527
		x"92",	--3528
		x"24",	--3529
		x"93",	--3530
		x"24",	--3531
		x"93",	--3532
		x"24",	--3533
		x"4f",	--3534
		x"00",	--3535
		x"9e",	--3536
		x"00",	--3537
		x"24",	--3538
		x"93",	--3539
		x"20",	--3540
		x"43",	--3541
		x"4e",	--3542
		x"41",	--3543
		x"41",	--3544
		x"93",	--3545
		x"24",	--3546
		x"93",	--3547
		x"00",	--3548
		x"23",	--3549
		x"43",	--3550
		x"4e",	--3551
		x"41",	--3552
		x"41",	--3553
		x"93",	--3554
		x"00",	--3555
		x"27",	--3556
		x"43",	--3557
		x"3f",	--3558
		x"4f",	--3559
		x"00",	--3560
		x"4e",	--3561
		x"00",	--3562
		x"9b",	--3563
		x"3b",	--3564
		x"9c",	--3565
		x"38",	--3566
		x"4f",	--3567
		x"00",	--3568
		x"4f",	--3569
		x"00",	--3570
		x"4e",	--3571
		x"00",	--3572
		x"4e",	--3573
		x"00",	--3574
		x"9f",	--3575
		x"2b",	--3576
		x"9e",	--3577
		x"28",	--3578
		x"9b",	--3579
		x"2b",	--3580
		x"9e",	--3581
		x"28",	--3582
		x"9f",	--3583
		x"28",	--3584
		x"9c",	--3585
		x"28",	--3586
		x"43",	--3587
		x"3f",	--3588
		x"93",	--3589
		x"23",	--3590
		x"43",	--3591
		x"3f",	--3592
		x"92",	--3593
		x"23",	--3594
		x"4e",	--3595
		x"00",	--3596
		x"4f",	--3597
		x"00",	--3598
		x"8f",	--3599
		x"3f",	--3600
		x"42",	--3601
		x"02",	--3602
		x"93",	--3603
		x"38",	--3604
		x"42",	--3605
		x"02",	--3606
		x"4f",	--3607
		x"00",	--3608
		x"53",	--3609
		x"4d",	--3610
		x"02",	--3611
		x"53",	--3612
		x"4e",	--3613
		x"02",	--3614
		x"41",	--3615
		x"43",	--3616
		x"41",	--3617
		x"12",	--3618
		x"12",	--3619
		x"83",	--3620
		x"4e",	--3621
		x"00",	--3622
		x"42",	--3623
		x"02",	--3624
		x"42",	--3625
		x"02",	--3626
		x"4e",	--3627
		x"4f",	--3628
		x"40",	--3629
		x"dc",	--3630
		x"12",	--3631
		x"de",	--3632
		x"9b",	--3633
		x"38",	--3634
		x"4a",	--3635
		x"5b",	--3636
		x"43",	--3637
		x"ff",	--3638
		x"3c",	--3639
		x"42",	--3640
		x"02",	--3641
		x"43",	--3642
		x"00",	--3643
		x"53",	--3644
		x"41",	--3645
		x"41",	--3646
		x"41",	--3647
		x"41",	--3648
		x"00",	--3649
		x"02",	--3650
		x"40",	--3651
		x"7f",	--3652
		x"02",	--3653
		x"41",	--3654
		x"50",	--3655
		x"00",	--3656
		x"41",	--3657
		x"00",	--3658
		x"12",	--3659
		x"dc",	--3660
		x"41",	--3661
		x"41",	--3662
		x"00",	--3663
		x"02",	--3664
		x"41",	--3665
		x"00",	--3666
		x"02",	--3667
		x"41",	--3668
		x"52",	--3669
		x"41",	--3670
		x"00",	--3671
		x"12",	--3672
		x"dc",	--3673
		x"41",	--3674
		x"4e",	--3675
		x"4f",	--3676
		x"02",	--3677
		x"40",	--3678
		x"7f",	--3679
		x"02",	--3680
		x"4d",	--3681
		x"4c",	--3682
		x"12",	--3683
		x"dc",	--3684
		x"41",	--3685
		x"4f",	--3686
		x"02",	--3687
		x"4e",	--3688
		x"02",	--3689
		x"4c",	--3690
		x"4d",	--3691
		x"12",	--3692
		x"dc",	--3693
		x"41",	--3694
		x"12",	--3695
		x"12",	--3696
		x"12",	--3697
		x"12",	--3698
		x"12",	--3699
		x"12",	--3700
		x"12",	--3701
		x"12",	--3702
		x"82",	--3703
		x"4f",	--3704
		x"4e",	--3705
		x"00",	--3706
		x"4d",	--3707
		x"41",	--3708
		x"00",	--3709
		x"41",	--3710
		x"00",	--3711
		x"4d",	--3712
		x"4d",	--3713
		x"10",	--3714
		x"44",	--3715
		x"4f",	--3716
		x"b0",	--3717
		x"00",	--3718
		x"24",	--3719
		x"40",	--3720
		x"00",	--3721
		x"00",	--3722
		x"4f",	--3723
		x"10",	--3724
		x"f3",	--3725
		x"24",	--3726
		x"40",	--3727
		x"00",	--3728
		x"3c",	--3729
		x"40",	--3730
		x"00",	--3731
		x"4e",	--3732
		x"00",	--3733
		x"41",	--3734
		x"53",	--3735
		x"3c",	--3736
		x"f0",	--3737
		x"00",	--3738
		x"24",	--3739
		x"40",	--3740
		x"00",	--3741
		x"00",	--3742
		x"3c",	--3743
		x"93",	--3744
		x"24",	--3745
		x"4d",	--3746
		x"00",	--3747
		x"41",	--3748
		x"53",	--3749
		x"3c",	--3750
		x"41",	--3751
		x"4c",	--3752
		x"10",	--3753
		x"11",	--3754
		x"10",	--3755
		x"11",	--3756
		x"4c",	--3757
		x"41",	--3758
		x"41",	--3759
		x"10",	--3760
		x"11",	--3761
		x"10",	--3762
		x"11",	--3763
		x"4c",	--3764
		x"86",	--3765
		x"77",	--3766
		x"4f",	--3767
		x"10",	--3768
		x"4e",	--3769
		x"00",	--3770
		x"f2",	--3771
		x"24",	--3772
		x"45",	--3773
		x"3c",	--3774
		x"43",	--3775
		x"4f",	--3776
		x"b0",	--3777
		x"00",	--3778
		x"20",	--3779
		x"41",	--3780
		x"00",	--3781
		x"53",	--3782
		x"53",	--3783
		x"93",	--3784
		x"00",	--3785
		x"23",	--3786
		x"81",	--3787
		x"00",	--3788
		x"9a",	--3789
		x"28",	--3790
		x"8a",	--3791
		x"3c",	--3792
		x"43",	--3793
		x"b3",	--3794
		x"00",	--3795
		x"24",	--3796
		x"95",	--3797
		x"28",	--3798
		x"85",	--3799
		x"3c",	--3800
		x"43",	--3801
		x"4d",	--3802
		x"9d",	--3803
		x"2c",	--3804
		x"47",	--3805
		x"93",	--3806
		x"38",	--3807
		x"40",	--3808
		x"00",	--3809
		x"00",	--3810
		x"43",	--3811
		x"43",	--3812
		x"3c",	--3813
		x"41",	--3814
		x"56",	--3815
		x"4f",	--3816
		x"11",	--3817
		x"53",	--3818
		x"12",	--3819
		x"3c",	--3820
		x"43",	--3821
		x"9a",	--3822
		x"3b",	--3823
		x"4a",	--3824
		x"40",	--3825
		x"00",	--3826
		x"00",	--3827
		x"8b",	--3828
		x"3c",	--3829
		x"41",	--3830
		x"00",	--3831
		x"11",	--3832
		x"12",	--3833
		x"53",	--3834
		x"45",	--3835
		x"5b",	--3836
		x"99",	--3837
		x"2b",	--3838
		x"3c",	--3839
		x"43",	--3840
		x"43",	--3841
		x"3c",	--3842
		x"53",	--3843
		x"41",	--3844
		x"56",	--3845
		x"4f",	--3846
		x"11",	--3847
		x"53",	--3848
		x"12",	--3849
		x"9a",	--3850
		x"3b",	--3851
		x"b3",	--3852
		x"00",	--3853
		x"24",	--3854
		x"44",	--3855
		x"3c",	--3856
		x"41",	--3857
		x"00",	--3858
		x"8b",	--3859
		x"3c",	--3860
		x"40",	--3861
		x"00",	--3862
		x"12",	--3863
		x"53",	--3864
		x"93",	--3865
		x"23",	--3866
		x"44",	--3867
		x"54",	--3868
		x"3f",	--3869
		x"53",	--3870
		x"11",	--3871
		x"12",	--3872
		x"53",	--3873
		x"4a",	--3874
		x"5b",	--3875
		x"4f",	--3876
		x"93",	--3877
		x"24",	--3878
		x"93",	--3879
		x"23",	--3880
		x"3c",	--3881
		x"40",	--3882
		x"00",	--3883
		x"12",	--3884
		x"53",	--3885
		x"99",	--3886
		x"2b",	--3887
		x"4b",	--3888
		x"52",	--3889
		x"41",	--3890
		x"41",	--3891
		x"41",	--3892
		x"41",	--3893
		x"41",	--3894
		x"41",	--3895
		x"41",	--3896
		x"41",	--3897
		x"41",	--3898
		x"12",	--3899
		x"12",	--3900
		x"12",	--3901
		x"12",	--3902
		x"12",	--3903
		x"12",	--3904
		x"12",	--3905
		x"12",	--3906
		x"50",	--3907
		x"ff",	--3908
		x"4f",	--3909
		x"00",	--3910
		x"4e",	--3911
		x"4d",	--3912
		x"4e",	--3913
		x"00",	--3914
		x"43",	--3915
		x"00",	--3916
		x"43",	--3917
		x"00",	--3918
		x"43",	--3919
		x"00",	--3920
		x"43",	--3921
		x"00",	--3922
		x"43",	--3923
		x"00",	--3924
		x"43",	--3925
		x"00",	--3926
		x"43",	--3927
		x"43",	--3928
		x"00",	--3929
		x"41",	--3930
		x"50",	--3931
		x"00",	--3932
		x"4e",	--3933
		x"00",	--3934
		x"40",	--3935
		x"e4",	--3936
		x"46",	--3937
		x"53",	--3938
		x"4f",	--3939
		x"00",	--3940
		x"93",	--3941
		x"20",	--3942
		x"90",	--3943
		x"00",	--3944
		x"20",	--3945
		x"43",	--3946
		x"00",	--3947
		x"43",	--3948
		x"00",	--3949
		x"46",	--3950
		x"00",	--3951
		x"43",	--3952
		x"00",	--3953
		x"43",	--3954
		x"00",	--3955
		x"43",	--3956
		x"00",	--3957
		x"43",	--3958
		x"00",	--3959
		x"43",	--3960
		x"00",	--3961
		x"40",	--3962
		x"e4",	--3963
		x"47",	--3964
		x"11",	--3965
		x"4e",	--3966
		x"12",	--3967
		x"00",	--3968
		x"53",	--3969
		x"00",	--3970
		x"40",	--3971
		x"e4",	--3972
		x"90",	--3973
		x"00",	--3974
		x"24",	--3975
		x"90",	--3976
		x"00",	--3977
		x"34",	--3978
		x"90",	--3979
		x"00",	--3980
		x"24",	--3981
		x"90",	--3982
		x"00",	--3983
		x"34",	--3984
		x"90",	--3985
		x"00",	--3986
		x"24",	--3987
		x"90",	--3988
		x"00",	--3989
		x"34",	--3990
		x"90",	--3991
		x"00",	--3992
		x"24",	--3993
		x"90",	--3994
		x"00",	--3995
		x"27",	--3996
		x"90",	--3997
		x"00",	--3998
		x"20",	--3999
		x"3c",	--4000
		x"90",	--4001
		x"00",	--4002
		x"24",	--4003
		x"90",	--4004
		x"00",	--4005
		x"24",	--4006
		x"90",	--4007
		x"00",	--4008
		x"20",	--4009
		x"3c",	--4010
		x"90",	--4011
		x"00",	--4012
		x"38",	--4013
		x"90",	--4014
		x"00",	--4015
		x"20",	--4016
		x"3c",	--4017
		x"90",	--4018
		x"00",	--4019
		x"24",	--4020
		x"90",	--4021
		x"00",	--4022
		x"34",	--4023
		x"90",	--4024
		x"00",	--4025
		x"24",	--4026
		x"90",	--4027
		x"00",	--4028
		x"24",	--4029
		x"90",	--4030
		x"00",	--4031
		x"20",	--4032
		x"3c",	--4033
		x"90",	--4034
		x"00",	--4035
		x"24",	--4036
		x"90",	--4037
		x"00",	--4038
		x"34",	--4039
		x"90",	--4040
		x"00",	--4041
		x"20",	--4042
		x"3c",	--4043
		x"90",	--4044
		x"00",	--4045
		x"24",	--4046
		x"90",	--4047
		x"00",	--4048
		x"24",	--4049
		x"41",	--4050
		x"00",	--4051
		x"41",	--4052
		x"00",	--4053
		x"89",	--4054
		x"40",	--4055
		x"e4",	--4056
		x"42",	--4057
		x"00",	--4058
		x"3c",	--4059
		x"d2",	--4060
		x"00",	--4061
		x"40",	--4062
		x"e4",	--4063
		x"41",	--4064
		x"f3",	--4065
		x"41",	--4066
		x"24",	--4067
		x"f0",	--4068
		x"ff",	--4069
		x"d3",	--4070
		x"3c",	--4071
		x"d3",	--4072
		x"4e",	--4073
		x"00",	--4074
		x"40",	--4075
		x"e4",	--4076
		x"d0",	--4077
		x"00",	--4078
		x"00",	--4079
		x"40",	--4080
		x"e4",	--4081
		x"40",	--4082
		x"00",	--4083
		x"00",	--4084
		x"40",	--4085
		x"e4",	--4086
		x"90",	--4087
		x"00",	--4088
		x"00",	--4089
		x"20",	--4090
		x"40",	--4091
		x"e4",	--4092
		x"40",	--4093
		x"00",	--4094
		x"00",	--4095
		x"40",	--4096
		x"e4",	--4097
		x"93",	--4098
		x"00",	--4099
		x"24",	--4100
		x"40",	--4101
		x"e4",	--4102
		x"43",	--4103
		x"00",	--4104
		x"40",	--4105
		x"e4",	--4106
		x"45",	--4107
		x"53",	--4108
		x"45",	--4109
		x"93",	--4110
		x"38",	--4111
		x"4a",	--4112
		x"00",	--4113
		x"3c",	--4114
		x"93",	--4115
		x"00",	--4116
		x"24",	--4117
		x"40",	--4118
		x"e4",	--4119
		x"d0",	--4120
		x"00",	--4121
		x"00",	--4122
		x"e3",	--4123
		x"4a",	--4124
		x"00",	--4125
		x"53",	--4126
		x"00",	--4127
		x"4e",	--4128
		x"3c",	--4129
		x"93",	--4130
		x"00",	--4131
		x"20",	--4132
		x"93",	--4133
		x"00",	--4134
		x"20",	--4135
		x"41",	--4136
		x"f0",	--4137
		x"00",	--4138
		x"43",	--4139
		x"24",	--4140
		x"43",	--4141
		x"4e",	--4142
		x"11",	--4143
		x"43",	--4144
		x"10",	--4145
		x"41",	--4146
		x"f0",	--4147
		x"00",	--4148
		x"de",	--4149
		x"4a",	--4150
		x"00",	--4151
		x"40",	--4152
		x"e4",	--4153
		x"41",	--4154
		x"00",	--4155
		x"5a",	--4156
		x"4a",	--4157
		x"5c",	--4158
		x"5c",	--4159
		x"5c",	--4160
		x"4a",	--4161
		x"00",	--4162
		x"50",	--4163
		x"ff",	--4164
		x"00",	--4165
		x"11",	--4166
		x"5e",	--4167
		x"00",	--4168
		x"43",	--4169
		x"00",	--4170
		x"40",	--4171
		x"e4",	--4172
		x"45",	--4173
		x"53",	--4174
		x"45",	--4175
		x"93",	--4176
		x"00",	--4177
		x"20",	--4178
		x"93",	--4179
		x"00",	--4180
		x"27",	--4181
		x"4e",	--4182
		x"00",	--4183
		x"43",	--4184
		x"00",	--4185
		x"41",	--4186
		x"52",	--4187
		x"3c",	--4188
		x"45",	--4189
		x"53",	--4190
		x"45",	--4191
		x"93",	--4192
		x"00",	--4193
		x"24",	--4194
		x"d2",	--4195
		x"00",	--4196
		x"41",	--4197
		x"00",	--4198
		x"4f",	--4199
		x"00",	--4200
		x"3c",	--4201
		x"93",	--4202
		x"00",	--4203
		x"24",	--4204
		x"41",	--4205
		x"00",	--4206
		x"00",	--4207
		x"93",	--4208
		x"20",	--4209
		x"40",	--4210
		x"ea",	--4211
		x"12",	--4212
		x"00",	--4213
		x"12",	--4214
		x"00",	--4215
		x"41",	--4216
		x"00",	--4217
		x"41",	--4218
		x"00",	--4219
		x"12",	--4220
		x"dc",	--4221
		x"52",	--4222
		x"5f",	--4223
		x"00",	--4224
		x"47",	--4225
		x"40",	--4226
		x"e4",	--4227
		x"45",	--4228
		x"53",	--4229
		x"45",	--4230
		x"49",	--4231
		x"00",	--4232
		x"43",	--4233
		x"93",	--4234
		x"20",	--4235
		x"43",	--4236
		x"5e",	--4237
		x"5e",	--4238
		x"5e",	--4239
		x"41",	--4240
		x"f0",	--4241
		x"ff",	--4242
		x"de",	--4243
		x"4a",	--4244
		x"00",	--4245
		x"47",	--4246
		x"40",	--4247
		x"00",	--4248
		x"00",	--4249
		x"3c",	--4250
		x"d3",	--4251
		x"00",	--4252
		x"3c",	--4253
		x"d2",	--4254
		x"00",	--4255
		x"40",	--4256
		x"00",	--4257
		x"00",	--4258
		x"3c",	--4259
		x"40",	--4260
		x"00",	--4261
		x"00",	--4262
		x"41",	--4263
		x"b3",	--4264
		x"24",	--4265
		x"45",	--4266
		x"52",	--4267
		x"45",	--4268
		x"45",	--4269
		x"00",	--4270
		x"45",	--4271
		x"00",	--4272
		x"45",	--4273
		x"00",	--4274
		x"48",	--4275
		x"00",	--4276
		x"47",	--4277
		x"00",	--4278
		x"46",	--4279
		x"00",	--4280
		x"4b",	--4281
		x"00",	--4282
		x"43",	--4283
		x"00",	--4284
		x"93",	--4285
		x"20",	--4286
		x"93",	--4287
		x"20",	--4288
		x"93",	--4289
		x"20",	--4290
		x"93",	--4291
		x"24",	--4292
		x"43",	--4293
		x"00",	--4294
		x"5b",	--4295
		x"43",	--4296
		x"6b",	--4297
		x"4b",	--4298
		x"00",	--4299
		x"4c",	--4300
		x"3c",	--4301
		x"f3",	--4302
		x"45",	--4303
		x"24",	--4304
		x"52",	--4305
		x"45",	--4306
		x"45",	--4307
		x"00",	--4308
		x"48",	--4309
		x"00",	--4310
		x"4b",	--4311
		x"00",	--4312
		x"43",	--4313
		x"00",	--4314
		x"93",	--4315
		x"20",	--4316
		x"3c",	--4317
		x"53",	--4318
		x"45",	--4319
		x"4b",	--4320
		x"00",	--4321
		x"43",	--4322
		x"00",	--4323
		x"93",	--4324
		x"24",	--4325
		x"43",	--4326
		x"00",	--4327
		x"5b",	--4328
		x"43",	--4329
		x"6b",	--4330
		x"4b",	--4331
		x"00",	--4332
		x"47",	--4333
		x"b2",	--4334
		x"00",	--4335
		x"24",	--4336
		x"93",	--4337
		x"00",	--4338
		x"20",	--4339
		x"41",	--4340
		x"90",	--4341
		x"00",	--4342
		x"00",	--4343
		x"20",	--4344
		x"d0",	--4345
		x"00",	--4346
		x"3c",	--4347
		x"92",	--4348
		x"00",	--4349
		x"20",	--4350
		x"d0",	--4351
		x"00",	--4352
		x"48",	--4353
		x"00",	--4354
		x"41",	--4355
		x"b2",	--4356
		x"24",	--4357
		x"93",	--4358
		x"00",	--4359
		x"24",	--4360
		x"40",	--4361
		x"00",	--4362
		x"00",	--4363
		x"b3",	--4364
		x"24",	--4365
		x"e3",	--4366
		x"00",	--4367
		x"e3",	--4368
		x"00",	--4369
		x"e3",	--4370
		x"00",	--4371
		x"e3",	--4372
		x"00",	--4373
		x"53",	--4374
		x"00",	--4375
		x"63",	--4376
		x"00",	--4377
		x"63",	--4378
		x"00",	--4379
		x"63",	--4380
		x"00",	--4381
		x"3c",	--4382
		x"b3",	--4383
		x"24",	--4384
		x"41",	--4385
		x"00",	--4386
		x"41",	--4387
		x"00",	--4388
		x"e3",	--4389
		x"e3",	--4390
		x"4a",	--4391
		x"4b",	--4392
		x"53",	--4393
		x"63",	--4394
		x"4e",	--4395
		x"00",	--4396
		x"4f",	--4397
		x"00",	--4398
		x"3c",	--4399
		x"41",	--4400
		x"00",	--4401
		x"e3",	--4402
		x"53",	--4403
		x"4a",	--4404
		x"00",	--4405
		x"43",	--4406
		x"00",	--4407
		x"b3",	--4408
		x"24",	--4409
		x"41",	--4410
		x"00",	--4411
		x"41",	--4412
		x"00",	--4413
		x"00",	--4414
		x"41",	--4415
		x"00",	--4416
		x"41",	--4417
		x"00",	--4418
		x"41",	--4419
		x"50",	--4420
		x"00",	--4421
		x"46",	--4422
		x"41",	--4423
		x"00",	--4424
		x"00",	--4425
		x"41",	--4426
		x"00",	--4427
		x"10",	--4428
		x"11",	--4429
		x"10",	--4430
		x"11",	--4431
		x"4b",	--4432
		x"00",	--4433
		x"4b",	--4434
		x"00",	--4435
		x"4b",	--4436
		x"00",	--4437
		x"12",	--4438
		x"00",	--4439
		x"12",	--4440
		x"00",	--4441
		x"12",	--4442
		x"00",	--4443
		x"12",	--4444
		x"00",	--4445
		x"49",	--4446
		x"41",	--4447
		x"00",	--4448
		x"48",	--4449
		x"44",	--4450
		x"12",	--4451
		x"e6",	--4452
		x"52",	--4453
		x"4c",	--4454
		x"90",	--4455
		x"00",	--4456
		x"34",	--4457
		x"50",	--4458
		x"00",	--4459
		x"4b",	--4460
		x"00",	--4461
		x"3c",	--4462
		x"4c",	--4463
		x"b3",	--4464
		x"00",	--4465
		x"24",	--4466
		x"40",	--4467
		x"00",	--4468
		x"3c",	--4469
		x"40",	--4470
		x"00",	--4471
		x"5b",	--4472
		x"4a",	--4473
		x"00",	--4474
		x"47",	--4475
		x"53",	--4476
		x"12",	--4477
		x"00",	--4478
		x"12",	--4479
		x"00",	--4480
		x"12",	--4481
		x"00",	--4482
		x"12",	--4483
		x"00",	--4484
		x"49",	--4485
		x"41",	--4486
		x"00",	--4487
		x"48",	--4488
		x"44",	--4489
		x"12",	--4490
		x"e6",	--4491
		x"52",	--4492
		x"4c",	--4493
		x"4d",	--4494
		x"00",	--4495
		x"4e",	--4496
		x"4f",	--4497
		x"53",	--4498
		x"93",	--4499
		x"23",	--4500
		x"93",	--4501
		x"23",	--4502
		x"93",	--4503
		x"23",	--4504
		x"93",	--4505
		x"23",	--4506
		x"43",	--4507
		x"00",	--4508
		x"43",	--4509
		x"00",	--4510
		x"43",	--4511
		x"00",	--4512
		x"43",	--4513
		x"00",	--4514
		x"3c",	--4515
		x"b3",	--4516
		x"24",	--4517
		x"41",	--4518
		x"00",	--4519
		x"41",	--4520
		x"00",	--4521
		x"41",	--4522
		x"50",	--4523
		x"00",	--4524
		x"41",	--4525
		x"00",	--4526
		x"10",	--4527
		x"11",	--4528
		x"10",	--4529
		x"11",	--4530
		x"41",	--4531
		x"00",	--4532
		x"49",	--4533
		x"44",	--4534
		x"47",	--4535
		x"12",	--4536
		x"e5",	--4537
		x"4e",	--4538
		x"90",	--4539
		x"00",	--4540
		x"34",	--4541
		x"50",	--4542
		x"00",	--4543
		x"4b",	--4544
		x"00",	--4545
		x"3c",	--4546
		x"4e",	--4547
		x"b3",	--4548
		x"00",	--4549
		x"24",	--4550
		x"40",	--4551
		x"00",	--4552
		x"3c",	--4553
		x"40",	--4554
		x"00",	--4555
		x"5b",	--4556
		x"4a",	--4557
		x"00",	--4558
		x"48",	--4559
		x"53",	--4560
		x"41",	--4561
		x"00",	--4562
		x"49",	--4563
		x"44",	--4564
		x"47",	--4565
		x"12",	--4566
		x"e5",	--4567
		x"4e",	--4568
		x"4f",	--4569
		x"53",	--4570
		x"93",	--4571
		x"23",	--4572
		x"93",	--4573
		x"23",	--4574
		x"43",	--4575
		x"00",	--4576
		x"43",	--4577
		x"00",	--4578
		x"3c",	--4579
		x"41",	--4580
		x"00",	--4581
		x"41",	--4582
		x"50",	--4583
		x"00",	--4584
		x"41",	--4585
		x"00",	--4586
		x"47",	--4587
		x"12",	--4588
		x"e5",	--4589
		x"4f",	--4590
		x"90",	--4591
		x"00",	--4592
		x"34",	--4593
		x"50",	--4594
		x"00",	--4595
		x"4d",	--4596
		x"00",	--4597
		x"3c",	--4598
		x"4f",	--4599
		x"b3",	--4600
		x"00",	--4601
		x"24",	--4602
		x"40",	--4603
		x"00",	--4604
		x"3c",	--4605
		x"40",	--4606
		x"00",	--4607
		x"5d",	--4608
		x"4c",	--4609
		x"00",	--4610
		x"48",	--4611
		x"53",	--4612
		x"41",	--4613
		x"00",	--4614
		x"47",	--4615
		x"12",	--4616
		x"e5",	--4617
		x"4f",	--4618
		x"53",	--4619
		x"93",	--4620
		x"23",	--4621
		x"43",	--4622
		x"00",	--4623
		x"90",	--4624
		x"00",	--4625
		x"00",	--4626
		x"24",	--4627
		x"43",	--4628
		x"00",	--4629
		x"93",	--4630
		x"00",	--4631
		x"24",	--4632
		x"41",	--4633
		x"50",	--4634
		x"00",	--4635
		x"4f",	--4636
		x"00",	--4637
		x"41",	--4638
		x"00",	--4639
		x"10",	--4640
		x"11",	--4641
		x"10",	--4642
		x"11",	--4643
		x"4a",	--4644
		x"00",	--4645
		x"46",	--4646
		x"00",	--4647
		x"46",	--4648
		x"10",	--4649
		x"11",	--4650
		x"10",	--4651
		x"11",	--4652
		x"4a",	--4653
		x"00",	--4654
		x"41",	--4655
		x"00",	--4656
		x"41",	--4657
		x"00",	--4658
		x"81",	--4659
		x"00",	--4660
		x"71",	--4661
		x"00",	--4662
		x"83",	--4663
		x"91",	--4664
		x"00",	--4665
		x"2c",	--4666
		x"d3",	--4667
		x"00",	--4668
		x"41",	--4669
		x"00",	--4670
		x"8c",	--4671
		x"4e",	--4672
		x"00",	--4673
		x"3c",	--4674
		x"93",	--4675
		x"00",	--4676
		x"24",	--4677
		x"41",	--4678
		x"00",	--4679
		x"00",	--4680
		x"12",	--4681
		x"00",	--4682
		x"12",	--4683
		x"00",	--4684
		x"41",	--4685
		x"00",	--4686
		x"46",	--4687
		x"53",	--4688
		x"41",	--4689
		x"00",	--4690
		x"12",	--4691
		x"dc",	--4692
		x"52",	--4693
		x"5f",	--4694
		x"00",	--4695
		x"3c",	--4696
		x"49",	--4697
		x"11",	--4698
		x"12",	--4699
		x"00",	--4700
		x"49",	--4701
		x"58",	--4702
		x"91",	--4703
		x"00",	--4704
		x"2b",	--4705
		x"49",	--4706
		x"00",	--4707
		x"4e",	--4708
		x"00",	--4709
		x"43",	--4710
		x"3c",	--4711
		x"41",	--4712
		x"00",	--4713
		x"00",	--4714
		x"43",	--4715
		x"00",	--4716
		x"43",	--4717
		x"00",	--4718
		x"3c",	--4719
		x"4e",	--4720
		x"43",	--4721
		x"00",	--4722
		x"43",	--4723
		x"00",	--4724
		x"43",	--4725
		x"41",	--4726
		x"00",	--4727
		x"46",	--4728
		x"93",	--4729
		x"24",	--4730
		x"40",	--4731
		x"de",	--4732
		x"41",	--4733
		x"00",	--4734
		x"50",	--4735
		x"00",	--4736
		x"41",	--4737
		x"41",	--4738
		x"41",	--4739
		x"41",	--4740
		x"41",	--4741
		x"41",	--4742
		x"41",	--4743
		x"41",	--4744
		x"41",	--4745
		x"43",	--4746
		x"93",	--4747
		x"34",	--4748
		x"40",	--4749
		x"00",	--4750
		x"e3",	--4751
		x"53",	--4752
		x"93",	--4753
		x"34",	--4754
		x"e3",	--4755
		x"e3",	--4756
		x"53",	--4757
		x"12",	--4758
		x"12",	--4759
		x"e5",	--4760
		x"41",	--4761
		x"b3",	--4762
		x"24",	--4763
		x"e3",	--4764
		x"53",	--4765
		x"b3",	--4766
		x"24",	--4767
		x"e3",	--4768
		x"53",	--4769
		x"41",	--4770
		x"12",	--4771
		x"e5",	--4772
		x"4e",	--4773
		x"41",	--4774
		x"12",	--4775
		x"12",	--4776
		x"12",	--4777
		x"40",	--4778
		x"00",	--4779
		x"4c",	--4780
		x"4d",	--4781
		x"43",	--4782
		x"43",	--4783
		x"5e",	--4784
		x"6f",	--4785
		x"6c",	--4786
		x"6d",	--4787
		x"9b",	--4788
		x"28",	--4789
		x"20",	--4790
		x"9a",	--4791
		x"28",	--4792
		x"8a",	--4793
		x"7b",	--4794
		x"d3",	--4795
		x"83",	--4796
		x"23",	--4797
		x"41",	--4798
		x"41",	--4799
		x"41",	--4800
		x"41",	--4801
		x"12",	--4802
		x"e5",	--4803
		x"4c",	--4804
		x"4d",	--4805
		x"41",	--4806
		x"12",	--4807
		x"43",	--4808
		x"93",	--4809
		x"34",	--4810
		x"40",	--4811
		x"00",	--4812
		x"e3",	--4813
		x"e3",	--4814
		x"53",	--4815
		x"63",	--4816
		x"93",	--4817
		x"34",	--4818
		x"e3",	--4819
		x"e3",	--4820
		x"e3",	--4821
		x"53",	--4822
		x"63",	--4823
		x"12",	--4824
		x"e5",	--4825
		x"b3",	--4826
		x"24",	--4827
		x"e3",	--4828
		x"e3",	--4829
		x"53",	--4830
		x"63",	--4831
		x"b3",	--4832
		x"24",	--4833
		x"e3",	--4834
		x"e3",	--4835
		x"53",	--4836
		x"63",	--4837
		x"41",	--4838
		x"41",	--4839
		x"12",	--4840
		x"e5",	--4841
		x"4c",	--4842
		x"4d",	--4843
		x"41",	--4844
		x"40",	--4845
		x"00",	--4846
		x"4e",	--4847
		x"43",	--4848
		x"5f",	--4849
		x"6e",	--4850
		x"9d",	--4851
		x"28",	--4852
		x"8d",	--4853
		x"d3",	--4854
		x"83",	--4855
		x"23",	--4856
		x"41",	--4857
		x"12",	--4858
		x"e5",	--4859
		x"4e",	--4860
		x"41",	--4861
		x"12",	--4862
		x"12",	--4863
		x"12",	--4864
		x"12",	--4865
		x"12",	--4866
		x"00",	--4867
		x"48",	--4868
		x"49",	--4869
		x"4a",	--4870
		x"4b",	--4871
		x"43",	--4872
		x"43",	--4873
		x"43",	--4874
		x"43",	--4875
		x"5c",	--4876
		x"6d",	--4877
		x"6e",	--4878
		x"6f",	--4879
		x"68",	--4880
		x"69",	--4881
		x"6a",	--4882
		x"6b",	--4883
		x"97",	--4884
		x"28",	--4885
		x"20",	--4886
		x"96",	--4887
		x"28",	--4888
		x"20",	--4889
		x"95",	--4890
		x"28",	--4891
		x"20",	--4892
		x"94",	--4893
		x"28",	--4894
		x"84",	--4895
		x"75",	--4896
		x"76",	--4897
		x"77",	--4898
		x"d3",	--4899
		x"83",	--4900
		x"00",	--4901
		x"23",	--4902
		x"53",	--4903
		x"41",	--4904
		x"41",	--4905
		x"41",	--4906
		x"41",	--4907
		x"41",	--4908
		x"12",	--4909
		x"12",	--4910
		x"12",	--4911
		x"12",	--4912
		x"41",	--4913
		x"00",	--4914
		x"41",	--4915
		x"00",	--4916
		x"41",	--4917
		x"00",	--4918
		x"41",	--4919
		x"00",	--4920
		x"12",	--4921
		x"e5",	--4922
		x"41",	--4923
		x"41",	--4924
		x"41",	--4925
		x"41",	--4926
		x"41",	--4927
		x"12",	--4928
		x"12",	--4929
		x"12",	--4930
		x"12",	--4931
		x"41",	--4932
		x"00",	--4933
		x"41",	--4934
		x"00",	--4935
		x"41",	--4936
		x"00",	--4937
		x"41",	--4938
		x"00",	--4939
		x"12",	--4940
		x"e5",	--4941
		x"48",	--4942
		x"49",	--4943
		x"4a",	--4944
		x"4b",	--4945
		x"41",	--4946
		x"41",	--4947
		x"41",	--4948
		x"41",	--4949
		x"41",	--4950
		x"12",	--4951
		x"12",	--4952
		x"12",	--4953
		x"12",	--4954
		x"12",	--4955
		x"41",	--4956
		x"00",	--4957
		x"41",	--4958
		x"00",	--4959
		x"41",	--4960
		x"00",	--4961
		x"41",	--4962
		x"00",	--4963
		x"12",	--4964
		x"e5",	--4965
		x"41",	--4966
		x"00",	--4967
		x"48",	--4968
		x"00",	--4969
		x"49",	--4970
		x"00",	--4971
		x"4a",	--4972
		x"00",	--4973
		x"4b",	--4974
		x"00",	--4975
		x"41",	--4976
		x"41",	--4977
		x"41",	--4978
		x"41",	--4979
		x"41",	--4980
		x"41",	--4981
		x"13",	--4982
		x"d0",	--4983
		x"00",	--4984
		x"3f",	--4985
		x"61",	--4986
		x"74",	--4987
		x"6e",	--4988
		x"20",	--4989
		x"6f",	--4990
		x"20",	--4991
		x"20",	--4992
		x"65",	--4993
		x"20",	--4994
		x"62",	--4995
		x"6e",	--4996
		x"66",	--4997
		x"6c",	--4998
		x"0d",	--4999
		x"00",	--5000
		x"65",	--5001
		x"73",	--5002
		x"6f",	--5003
		x"6c",	--5004
		x"20",	--5005
		x"6f",	--5006
		x"20",	--5007
		x"65",	--5008
		x"20",	--5009
		x"68",	--5010
		x"74",	--5011
		x"0a",	--5012
		x"53",	--5013
		x"6f",	--5014
		x"0d",	--5015
		x"00",	--5016
		x"72",	--5017
		x"6f",	--5018
		x"3a",	--5019
		x"6d",	--5020
		x"73",	--5021
		x"69",	--5022
		x"67",	--5023
		x"61",	--5024
		x"67",	--5025
		x"6d",	--5026
		x"6e",	--5027
		x"0d",	--5028
		x"00",	--5029
		x"6f",	--5030
		x"72",	--5031
		x"63",	--5032
		x"20",	--5033
		x"73",	--5034
		x"67",	--5035
		x"3a",	--5036
		x"0a",	--5037
		x"09",	--5038
		x"73",	--5039
		x"4c",	--5040
		x"46",	--5041
		x"20",	--5042
		x"49",	--5043
		x"48",	--5044
		x"20",	--5045
		x"54",	--5046
		x"4d",	--5047
		x"4f",	--5048
		x"54",	--5049
		x"0d",	--5050
		x"00",	--5051
		x"64",	--5052
		x"25",	--5053
		x"0d",	--5054
		x"00",	--5055
		x"6c",	--5056
		x"20",	--5057
		x"6c",	--5058
		x"00",	--5059
		x"73",	--5060
		x"0a",	--5061
		x"25",	--5062
		x"20",	--5063
		x"64",	--5064
		x"0a",	--5065
		x"00",	--5066
		x"c5",	--5067
		x"c5",	--5068
		x"c5",	--5069
		x"c5",	--5070
		x"c5",	--5071
		x"c6",	--5072
		x"c5",	--5073
		x"c5",	--5074
		x"0a",	--5075
		x"3d",	--5076
		x"3d",	--5077
		x"3d",	--5078
		x"4d",	--5079
		x"72",	--5080
		x"65",	--5081
		x"20",	--5082
		x"43",	--5083
		x"20",	--5084
		x"3d",	--5085
		x"3d",	--5086
		x"3d",	--5087
		x"0a",	--5088
		x"69",	--5089
		x"74",	--5090
		x"72",	--5091
		x"63",	--5092
		x"69",	--5093
		x"65",	--5094
		x"6d",	--5095
		x"64",	--5096
		x"00",	--5097
		x"72",	--5098
		x"74",	--5099
		x"00",	--5100
		x"65",	--5101
		x"64",	--5102
		x"62",	--5103
		x"7a",	--5104
		x"65",	--5105
		x"00",	--5106
		x"77",	--5107
		x"00",	--5108
		x"6e",	--5109
		x"6f",	--5110
		x"65",	--5111
		x"00",	--5112
		x"70",	--5113
		x"65",	--5114
		x"20",	--5115
		x"6f",	--5116
		x"74",	--5117
		x"6f",	--5118
		x"6c",	--5119
		x"72",	--5120
		x"73",	--5121
		x"65",	--5122
		x"64",	--5123
		x"63",	--5124
		x"6e",	--5125
		x"69",	--5126
		x"75",	--5127
		x"61",	--5128
		x"69",	--5129
		x"6e",	--5130
		x"62",	--5131
		x"6f",	--5132
		x"6c",	--5133
		x"61",	--5134
		x"65",	--5135
		x"00",	--5136
		x"0a",	--5137
		x"08",	--5138
		x"08",	--5139
		x"25",	--5140
		x"00",	--5141
		x"72",	--5142
		x"74",	--5143
		x"0a",	--5144
		x"00",	--5145
		x"72",	--5146
		x"6f",	--5147
		x"3a",	--5148
		x"6d",	--5149
		x"73",	--5150
		x"69",	--5151
		x"67",	--5152
		x"61",	--5153
		x"67",	--5154
		x"6d",	--5155
		x"6e",	--5156
		x"0d",	--5157
		x"00",	--5158
		x"6f",	--5159
		x"72",	--5160
		x"63",	--5161
		x"20",	--5162
		x"73",	--5163
		x"67",	--5164
		x"3a",	--5165
		x"0a",	--5166
		x"09",	--5167
		x"73",	--5168
		x"52",	--5169
		x"47",	--5170
		x"53",	--5171
		x"45",	--5172
		x"20",	--5173
		x"41",	--5174
		x"55",	--5175
		x"0d",	--5176
		x"00",	--5177
		x"3d",	--5178
		x"64",	--5179
		x"76",	--5180
		x"25",	--5181
		x"0d",	--5182
		x"00",	--5183
		x"25",	--5184
		x"20",	--5185
		x"45",	--5186
		x"49",	--5187
		x"54",	--5188
		x"52",	--5189
		x"0a",	--5190
		x"72",	--5191
		x"61",	--5192
		x"0a",	--5193
		x"00",	--5194
		x"63",	--5195
		x"69",	--5196
		x"20",	--5197
		x"6f",	--5198
		x"20",	--5199
		x"20",	--5200
		x"75",	--5201
		x"62",	--5202
		x"72",	--5203
		x"0a",	--5204
		x"25",	--5205
		x"20",	--5206
		x"73",	--5207
		x"0a",	--5208
		x"25",	--5209
		x"3a",	--5210
		x"6e",	--5211
		x"20",	--5212
		x"75",	--5213
		x"68",	--5214
		x"63",	--5215
		x"6d",	--5216
		x"61",	--5217
		x"64",	--5218
		x"0a",	--5219
		x"00",	--5220
		x"ce",	--5221
		x"cd",	--5222
		x"cd",	--5223
		x"cd",	--5224
		x"cd",	--5225
		x"cd",	--5226
		x"cd",	--5227
		x"cd",	--5228
		x"cd",	--5229
		x"cd",	--5230
		x"cd",	--5231
		x"cd",	--5232
		x"cd",	--5233
		x"cd",	--5234
		x"cd",	--5235
		x"cd",	--5236
		x"cd",	--5237
		x"cd",	--5238
		x"cd",	--5239
		x"cd",	--5240
		x"cd",	--5241
		x"cd",	--5242
		x"cd",	--5243
		x"cd",	--5244
		x"cd",	--5245
		x"cd",	--5246
		x"cd",	--5247
		x"cd",	--5248
		x"cd",	--5249
		x"ce",	--5250
		x"cd",	--5251
		x"cd",	--5252
		x"cd",	--5253
		x"cd",	--5254
		x"cd",	--5255
		x"cd",	--5256
		x"cd",	--5257
		x"cd",	--5258
		x"cd",	--5259
		x"cd",	--5260
		x"cd",	--5261
		x"cd",	--5262
		x"cd",	--5263
		x"cd",	--5264
		x"cd",	--5265
		x"cd",	--5266
		x"cd",	--5267
		x"cd",	--5268
		x"cd",	--5269
		x"cd",	--5270
		x"cd",	--5271
		x"cd",	--5272
		x"cd",	--5273
		x"cd",	--5274
		x"cd",	--5275
		x"cd",	--5276
		x"cd",	--5277
		x"cd",	--5278
		x"cd",	--5279
		x"cd",	--5280
		x"cd",	--5281
		x"ce",	--5282
		x"ce",	--5283
		x"ce",	--5284
		x"cd",	--5285
		x"cd",	--5286
		x"cd",	--5287
		x"cd",	--5288
		x"cd",	--5289
		x"cd",	--5290
		x"cd",	--5291
		x"ce",	--5292
		x"cd",	--5293
		x"ce",	--5294
		x"cd",	--5295
		x"cd",	--5296
		x"cd",	--5297
		x"cd",	--5298
		x"ce",	--5299
		x"cd",	--5300
		x"cd",	--5301
		x"cd",	--5302
		x"ce",	--5303
		x"ce",	--5304
		x"31",	--5305
		x"33",	--5306
		x"35",	--5307
		x"37",	--5308
		x"39",	--5309
		x"62",	--5310
		x"64",	--5311
		x"66",	--5312
		x"00",	--5313
		x"00",	--5314
		x"00",	--5315
		x"00",	--5316
		x"00",	--5317
		x"01",	--5318
		x"02",	--5319
		x"03",	--5320
		x"03",	--5321
		x"04",	--5322
		x"04",	--5323
		x"04",	--5324
		x"04",	--5325
		x"05",	--5326
		x"05",	--5327
		x"05",	--5328
		x"05",	--5329
		x"05",	--5330
		x"05",	--5331
		x"05",	--5332
		x"05",	--5333
		x"06",	--5334
		x"06",	--5335
		x"06",	--5336
		x"06",	--5337
		x"06",	--5338
		x"06",	--5339
		x"06",	--5340
		x"06",	--5341
		x"06",	--5342
		x"06",	--5343
		x"06",	--5344
		x"06",	--5345
		x"06",	--5346
		x"06",	--5347
		x"06",	--5348
		x"06",	--5349
		x"07",	--5350
		x"07",	--5351
		x"07",	--5352
		x"07",	--5353
		x"07",	--5354
		x"07",	--5355
		x"07",	--5356
		x"07",	--5357
		x"07",	--5358
		x"07",	--5359
		x"07",	--5360
		x"07",	--5361
		x"07",	--5362
		x"07",	--5363
		x"07",	--5364
		x"07",	--5365
		x"07",	--5366
		x"07",	--5367
		x"07",	--5368
		x"07",	--5369
		x"07",	--5370
		x"07",	--5371
		x"07",	--5372
		x"07",	--5373
		x"07",	--5374
		x"07",	--5375
		x"07",	--5376
		x"07",	--5377
		x"07",	--5378
		x"07",	--5379
		x"07",	--5380
		x"07",	--5381
		x"08",	--5382
		x"08",	--5383
		x"08",	--5384
		x"08",	--5385
		x"08",	--5386
		x"08",	--5387
		x"08",	--5388
		x"08",	--5389
		x"08",	--5390
		x"08",	--5391
		x"08",	--5392
		x"08",	--5393
		x"08",	--5394
		x"08",	--5395
		x"08",	--5396
		x"08",	--5397
		x"08",	--5398
		x"08",	--5399
		x"08",	--5400
		x"08",	--5401
		x"08",	--5402
		x"08",	--5403
		x"08",	--5404
		x"08",	--5405
		x"08",	--5406
		x"08",	--5407
		x"08",	--5408
		x"08",	--5409
		x"08",	--5410
		x"08",	--5411
		x"08",	--5412
		x"08",	--5413
		x"08",	--5414
		x"08",	--5415
		x"08",	--5416
		x"08",	--5417
		x"08",	--5418
		x"08",	--5419
		x"08",	--5420
		x"08",	--5421
		x"08",	--5422
		x"08",	--5423
		x"08",	--5424
		x"08",	--5425
		x"08",	--5426
		x"08",	--5427
		x"08",	--5428
		x"08",	--5429
		x"08",	--5430
		x"08",	--5431
		x"08",	--5432
		x"08",	--5433
		x"08",	--5434
		x"08",	--5435
		x"08",	--5436
		x"08",	--5437
		x"08",	--5438
		x"08",	--5439
		x"08",	--5440
		x"08",	--5441
		x"08",	--5442
		x"08",	--5443
		x"08",	--5444
		x"08",	--5445
		x"6e",	--5446
		x"6c",	--5447
		x"29",	--5448
		x"00",	--5449
		x"ff",	--5450
		x"ff",	--5451
		x"65",	--5452
		x"70",	--5453
		x"00",	--5454
		x"ff",	--5455
		x"ff",	--5456
		x"ff",	--5457
		x"ff",	--5458
		x"ff",	--5459
		x"ff",	--5460
		x"ff",	--5461
		x"ff",	--5462
		x"ff",	--5463
		x"ff",	--5464
		x"ff",	--5465
		x"ff",	--5466
		x"ff",	--5467
		x"ff",	--5468
		x"ff",	--5469
		x"ff",	--5470
		x"ff",	--5471
		x"ff",	--5472
		x"ff",	--5473
		x"ff",	--5474
		x"ff",	--5475
		x"ff",	--5476
		x"ff",	--5477
		x"ff",	--5478
		x"ff",	--5479
		x"ff",	--5480
		x"ff",	--5481
		x"ff",	--5482
		x"ff",	--5483
		x"ff",	--5484
		x"ff",	--5485
		x"ff",	--5486
		x"ff",	--5487
		x"ff",	--5488
		x"ff",	--5489
		x"ff",	--5490
		x"ff",	--5491
		x"ff",	--5492
		x"ff",	--5493
		x"ff",	--5494
		x"ff",	--5495
		x"ff",	--5496
		x"ff",	--5497
		x"ff",	--5498
		x"ff",	--5499
		x"ff",	--5500
		x"ff",	--5501
		x"ff",	--5502
		x"ff",	--5503
		x"ff",	--5504
		x"ff",	--5505
		x"ff",	--5506
		x"ff",	--5507
		x"ff",	--5508
		x"ff",	--5509
		x"ff",	--5510
		x"ff",	--5511
		x"ff",	--5512
		x"ff",	--5513
		x"ff",	--5514
		x"ff",	--5515
		x"ff",	--5516
		x"ff",	--5517
		x"ff",	--5518
		x"ff",	--5519
		x"ff",	--5520
		x"ff",	--5521
		x"ff",	--5522
		x"ff",	--5523
		x"ff",	--5524
		x"ff",	--5525
		x"ff",	--5526
		x"ff",	--5527
		x"ff",	--5528
		x"ff",	--5529
		x"ff",	--5530
		x"ff",	--5531
		x"ff",	--5532
		x"ff",	--5533
		x"ff",	--5534
		x"ff",	--5535
		x"ff",	--5536
		x"ff",	--5537
		x"ff",	--5538
		x"ff",	--5539
		x"ff",	--5540
		x"ff",	--5541
		x"ff",	--5542
		x"ff",	--5543
		x"ff",	--5544
		x"ff",	--5545
		x"ff",	--5546
		x"ff",	--5547
		x"ff",	--5548
		x"ff",	--5549
		x"ff",	--5550
		x"ff",	--5551
		x"ff",	--5552
		x"ff",	--5553
		x"ff",	--5554
		x"ff",	--5555
		x"ff",	--5556
		x"ff",	--5557
		x"ff",	--5558
		x"ff",	--5559
		x"ff",	--5560
		x"ff",	--5561
		x"ff",	--5562
		x"ff",	--5563
		x"ff",	--5564
		x"ff",	--5565
		x"ff",	--5566
		x"ff",	--5567
		x"ff",	--5568
		x"ff",	--5569
		x"ff",	--5570
		x"ff",	--5571
		x"ff",	--5572
		x"ff",	--5573
		x"ff",	--5574
		x"ff",	--5575
		x"ff",	--5576
		x"ff",	--5577
		x"ff",	--5578
		x"ff",	--5579
		x"ff",	--5580
		x"ff",	--5581
		x"ff",	--5582
		x"ff",	--5583
		x"ff",	--5584
		x"ff",	--5585
		x"ff",	--5586
		x"ff",	--5587
		x"ff",	--5588
		x"ff",	--5589
		x"ff",	--5590
		x"ff",	--5591
		x"ff",	--5592
		x"ff",	--5593
		x"ff",	--5594
		x"ff",	--5595
		x"ff",	--5596
		x"ff",	--5597
		x"ff",	--5598
		x"ff",	--5599
		x"ff",	--5600
		x"ff",	--5601
		x"ff",	--5602
		x"ff",	--5603
		x"ff",	--5604
		x"ff",	--5605
		x"ff",	--5606
		x"ff",	--5607
		x"ff",	--5608
		x"ff",	--5609
		x"ff",	--5610
		x"ff",	--5611
		x"ff",	--5612
		x"ff",	--5613
		x"ff",	--5614
		x"ff",	--5615
		x"ff",	--5616
		x"ff",	--5617
		x"ff",	--5618
		x"ff",	--5619
		x"ff",	--5620
		x"ff",	--5621
		x"ff",	--5622
		x"ff",	--5623
		x"ff",	--5624
		x"ff",	--5625
		x"ff",	--5626
		x"ff",	--5627
		x"ff",	--5628
		x"ff",	--5629
		x"ff",	--5630
		x"ff",	--5631
		x"ff",	--5632
		x"ff",	--5633
		x"ff",	--5634
		x"ff",	--5635
		x"ff",	--5636
		x"ff",	--5637
		x"ff",	--5638
		x"ff",	--5639
		x"ff",	--5640
		x"ff",	--5641
		x"ff",	--5642
		x"ff",	--5643
		x"ff",	--5644
		x"ff",	--5645
		x"ff",	--5646
		x"ff",	--5647
		x"ff",	--5648
		x"ff",	--5649
		x"ff",	--5650
		x"ff",	--5651
		x"ff",	--5652
		x"ff",	--5653
		x"ff",	--5654
		x"ff",	--5655
		x"ff",	--5656
		x"ff",	--5657
		x"ff",	--5658
		x"ff",	--5659
		x"ff",	--5660
		x"ff",	--5661
		x"ff",	--5662
		x"ff",	--5663
		x"ff",	--5664
		x"ff",	--5665
		x"ff",	--5666
		x"ff",	--5667
		x"ff",	--5668
		x"ff",	--5669
		x"ff",	--5670
		x"ff",	--5671
		x"ff",	--5672
		x"ff",	--5673
		x"ff",	--5674
		x"ff",	--5675
		x"ff",	--5676
		x"ff",	--5677
		x"ff",	--5678
		x"ff",	--5679
		x"ff",	--5680
		x"ff",	--5681
		x"ff",	--5682
		x"ff",	--5683
		x"ff",	--5684
		x"ff",	--5685
		x"ff",	--5686
		x"ff",	--5687
		x"ff",	--5688
		x"ff",	--5689
		x"ff",	--5690
		x"ff",	--5691
		x"ff",	--5692
		x"ff",	--5693
		x"ff",	--5694
		x"ff",	--5695
		x"ff",	--5696
		x"ff",	--5697
		x"ff",	--5698
		x"ff",	--5699
		x"ff",	--5700
		x"ff",	--5701
		x"ff",	--5702
		x"ff",	--5703
		x"ff",	--5704
		x"ff",	--5705
		x"ff",	--5706
		x"ff",	--5707
		x"ff",	--5708
		x"ff",	--5709
		x"ff",	--5710
		x"ff",	--5711
		x"ff",	--5712
		x"ff",	--5713
		x"ff",	--5714
		x"ff",	--5715
		x"ff",	--5716
		x"ff",	--5717
		x"ff",	--5718
		x"ff",	--5719
		x"ff",	--5720
		x"ff",	--5721
		x"ff",	--5722
		x"ff",	--5723
		x"ff",	--5724
		x"ff",	--5725
		x"ff",	--5726
		x"ff",	--5727
		x"ff",	--5728
		x"ff",	--5729
		x"ff",	--5730
		x"ff",	--5731
		x"ff",	--5732
		x"ff",	--5733
		x"ff",	--5734
		x"ff",	--5735
		x"ff",	--5736
		x"ff",	--5737
		x"ff",	--5738
		x"ff",	--5739
		x"ff",	--5740
		x"ff",	--5741
		x"ff",	--5742
		x"ff",	--5743
		x"ff",	--5744
		x"ff",	--5745
		x"ff",	--5746
		x"ff",	--5747
		x"ff",	--5748
		x"ff",	--5749
		x"ff",	--5750
		x"ff",	--5751
		x"ff",	--5752
		x"ff",	--5753
		x"ff",	--5754
		x"ff",	--5755
		x"ff",	--5756
		x"ff",	--5757
		x"ff",	--5758
		x"ff",	--5759
		x"ff",	--5760
		x"ff",	--5761
		x"ff",	--5762
		x"ff",	--5763
		x"ff",	--5764
		x"ff",	--5765
		x"ff",	--5766
		x"ff",	--5767
		x"ff",	--5768
		x"ff",	--5769
		x"ff",	--5770
		x"ff",	--5771
		x"ff",	--5772
		x"ff",	--5773
		x"ff",	--5774
		x"ff",	--5775
		x"ff",	--5776
		x"ff",	--5777
		x"ff",	--5778
		x"ff",	--5779
		x"ff",	--5780
		x"ff",	--5781
		x"ff",	--5782
		x"ff",	--5783
		x"ff",	--5784
		x"ff",	--5785
		x"ff",	--5786
		x"ff",	--5787
		x"ff",	--5788
		x"ff",	--5789
		x"ff",	--5790
		x"ff",	--5791
		x"ff",	--5792
		x"ff",	--5793
		x"ff",	--5794
		x"ff",	--5795
		x"ff",	--5796
		x"ff",	--5797
		x"ff",	--5798
		x"ff",	--5799
		x"ff",	--5800
		x"ff",	--5801
		x"ff",	--5802
		x"ff",	--5803
		x"ff",	--5804
		x"ff",	--5805
		x"ff",	--5806
		x"ff",	--5807
		x"ff",	--5808
		x"ff",	--5809
		x"ff",	--5810
		x"ff",	--5811
		x"ff",	--5812
		x"ff",	--5813
		x"ff",	--5814
		x"ff",	--5815
		x"ff",	--5816
		x"ff",	--5817
		x"ff",	--5818
		x"ff",	--5819
		x"ff",	--5820
		x"ff",	--5821
		x"ff",	--5822
		x"ff",	--5823
		x"ff",	--5824
		x"ff",	--5825
		x"ff",	--5826
		x"ff",	--5827
		x"ff",	--5828
		x"ff",	--5829
		x"ff",	--5830
		x"ff",	--5831
		x"ff",	--5832
		x"ff",	--5833
		x"ff",	--5834
		x"ff",	--5835
		x"ff",	--5836
		x"ff",	--5837
		x"ff",	--5838
		x"ff",	--5839
		x"ff",	--5840
		x"ff",	--5841
		x"ff",	--5842
		x"ff",	--5843
		x"ff",	--5844
		x"ff",	--5845
		x"ff",	--5846
		x"ff",	--5847
		x"ff",	--5848
		x"ff",	--5849
		x"ff",	--5850
		x"ff",	--5851
		x"ff",	--5852
		x"ff",	--5853
		x"ff",	--5854
		x"ff",	--5855
		x"ff",	--5856
		x"ff",	--5857
		x"ff",	--5858
		x"ff",	--5859
		x"ff",	--5860
		x"ff",	--5861
		x"ff",	--5862
		x"ff",	--5863
		x"ff",	--5864
		x"ff",	--5865
		x"ff",	--5866
		x"ff",	--5867
		x"ff",	--5868
		x"ff",	--5869
		x"ff",	--5870
		x"ff",	--5871
		x"ff",	--5872
		x"ff",	--5873
		x"ff",	--5874
		x"ff",	--5875
		x"ff",	--5876
		x"ff",	--5877
		x"ff",	--5878
		x"ff",	--5879
		x"ff",	--5880
		x"ff",	--5881
		x"ff",	--5882
		x"ff",	--5883
		x"ff",	--5884
		x"ff",	--5885
		x"ff",	--5886
		x"ff",	--5887
		x"ff",	--5888
		x"ff",	--5889
		x"ff",	--5890
		x"ff",	--5891
		x"ff",	--5892
		x"ff",	--5893
		x"ff",	--5894
		x"ff",	--5895
		x"ff",	--5896
		x"ff",	--5897
		x"ff",	--5898
		x"ff",	--5899
		x"ff",	--5900
		x"ff",	--5901
		x"ff",	--5902
		x"ff",	--5903
		x"ff",	--5904
		x"ff",	--5905
		x"ff",	--5906
		x"ff",	--5907
		x"ff",	--5908
		x"ff",	--5909
		x"ff",	--5910
		x"ff",	--5911
		x"ff",	--5912
		x"ff",	--5913
		x"ff",	--5914
		x"ff",	--5915
		x"ff",	--5916
		x"ff",	--5917
		x"ff",	--5918
		x"ff",	--5919
		x"ff",	--5920
		x"ff",	--5921
		x"ff",	--5922
		x"ff",	--5923
		x"ff",	--5924
		x"ff",	--5925
		x"ff",	--5926
		x"ff",	--5927
		x"ff",	--5928
		x"ff",	--5929
		x"ff",	--5930
		x"ff",	--5931
		x"ff",	--5932
		x"ff",	--5933
		x"ff",	--5934
		x"ff",	--5935
		x"ff",	--5936
		x"ff",	--5937
		x"ff",	--5938
		x"ff",	--5939
		x"ff",	--5940
		x"ff",	--5941
		x"ff",	--5942
		x"ff",	--5943
		x"ff",	--5944
		x"ff",	--5945
		x"ff",	--5946
		x"ff",	--5947
		x"ff",	--5948
		x"ff",	--5949
		x"ff",	--5950
		x"ff",	--5951
		x"ff",	--5952
		x"ff",	--5953
		x"ff",	--5954
		x"ff",	--5955
		x"ff",	--5956
		x"ff",	--5957
		x"ff",	--5958
		x"ff",	--5959
		x"ff",	--5960
		x"ff",	--5961
		x"ff",	--5962
		x"ff",	--5963
		x"ff",	--5964
		x"ff",	--5965
		x"ff",	--5966
		x"ff",	--5967
		x"ff",	--5968
		x"ff",	--5969
		x"ff",	--5970
		x"ff",	--5971
		x"ff",	--5972
		x"ff",	--5973
		x"ff",	--5974
		x"ff",	--5975
		x"ff",	--5976
		x"ff",	--5977
		x"ff",	--5978
		x"ff",	--5979
		x"ff",	--5980
		x"ff",	--5981
		x"ff",	--5982
		x"ff",	--5983
		x"ff",	--5984
		x"ff",	--5985
		x"ff",	--5986
		x"ff",	--5987
		x"ff",	--5988
		x"ff",	--5989
		x"ff",	--5990
		x"ff",	--5991
		x"ff",	--5992
		x"ff",	--5993
		x"ff",	--5994
		x"ff",	--5995
		x"ff",	--5996
		x"ff",	--5997
		x"ff",	--5998
		x"ff",	--5999
		x"ff",	--6000
		x"ff",	--6001
		x"ff",	--6002
		x"ff",	--6003
		x"ff",	--6004
		x"ff",	--6005
		x"ff",	--6006
		x"ff",	--6007
		x"ff",	--6008
		x"ff",	--6009
		x"ff",	--6010
		x"ff",	--6011
		x"ff",	--6012
		x"ff",	--6013
		x"ff",	--6014
		x"ff",	--6015
		x"ff",	--6016
		x"ff",	--6017
		x"ff",	--6018
		x"ff",	--6019
		x"ff",	--6020
		x"ff",	--6021
		x"ff",	--6022
		x"ff",	--6023
		x"ff",	--6024
		x"ff",	--6025
		x"ff",	--6026
		x"ff",	--6027
		x"ff",	--6028
		x"ff",	--6029
		x"ff",	--6030
		x"ff",	--6031
		x"ff",	--6032
		x"ff",	--6033
		x"ff",	--6034
		x"ff",	--6035
		x"ff",	--6036
		x"ff",	--6037
		x"ff",	--6038
		x"ff",	--6039
		x"ff",	--6040
		x"ff",	--6041
		x"ff",	--6042
		x"ff",	--6043
		x"ff",	--6044
		x"ff",	--6045
		x"ff",	--6046
		x"ff",	--6047
		x"ff",	--6048
		x"ff",	--6049
		x"ff",	--6050
		x"ff",	--6051
		x"ff",	--6052
		x"ff",	--6053
		x"ff",	--6054
		x"ff",	--6055
		x"ff",	--6056
		x"ff",	--6057
		x"ff",	--6058
		x"ff",	--6059
		x"ff",	--6060
		x"ff",	--6061
		x"ff",	--6062
		x"ff",	--6063
		x"ff",	--6064
		x"ff",	--6065
		x"ff",	--6066
		x"ff",	--6067
		x"ff",	--6068
		x"ff",	--6069
		x"ff",	--6070
		x"ff",	--6071
		x"ff",	--6072
		x"ff",	--6073
		x"ff",	--6074
		x"ff",	--6075
		x"ff",	--6076
		x"ff",	--6077
		x"ff",	--6078
		x"ff",	--6079
		x"ff",	--6080
		x"ff",	--6081
		x"ff",	--6082
		x"ff",	--6083
		x"ff",	--6084
		x"ff",	--6085
		x"ff",	--6086
		x"ff",	--6087
		x"ff",	--6088
		x"ff",	--6089
		x"ff",	--6090
		x"ff",	--6091
		x"ff",	--6092
		x"ff",	--6093
		x"ff",	--6094
		x"ff",	--6095
		x"ff",	--6096
		x"ff",	--6097
		x"ff",	--6098
		x"ff",	--6099
		x"ff",	--6100
		x"ff",	--6101
		x"ff",	--6102
		x"ff",	--6103
		x"ff",	--6104
		x"ff",	--6105
		x"ff",	--6106
		x"ff",	--6107
		x"ff",	--6108
		x"ff",	--6109
		x"ff",	--6110
		x"ff",	--6111
		x"ff",	--6112
		x"ff",	--6113
		x"ff",	--6114
		x"ff",	--6115
		x"ff",	--6116
		x"ff",	--6117
		x"ff",	--6118
		x"ff",	--6119
		x"ff",	--6120
		x"ff",	--6121
		x"ff",	--6122
		x"ff",	--6123
		x"ff",	--6124
		x"ff",	--6125
		x"ff",	--6126
		x"ff",	--6127
		x"ff",	--6128
		x"ff",	--6129
		x"ff",	--6130
		x"ff",	--6131
		x"ff",	--6132
		x"ff",	--6133
		x"ff",	--6134
		x"ff",	--6135
		x"ff",	--6136
		x"ff",	--6137
		x"ff",	--6138
		x"ff",	--6139
		x"ff",	--6140
		x"ff",	--6141
		x"ff",	--6142
		x"ff",	--6143
		x"ff",	--6144
		x"ff",	--6145
		x"ff",	--6146
		x"ff",	--6147
		x"ff",	--6148
		x"ff",	--6149
		x"ff",	--6150
		x"ff",	--6151
		x"ff",	--6152
		x"ff",	--6153
		x"ff",	--6154
		x"ff",	--6155
		x"ff",	--6156
		x"ff",	--6157
		x"ff",	--6158
		x"ff",	--6159
		x"ff",	--6160
		x"ff",	--6161
		x"ff",	--6162
		x"ff",	--6163
		x"ff",	--6164
		x"ff",	--6165
		x"ff",	--6166
		x"ff",	--6167
		x"ff",	--6168
		x"ff",	--6169
		x"ff",	--6170
		x"ff",	--6171
		x"ff",	--6172
		x"ff",	--6173
		x"ff",	--6174
		x"ff",	--6175
		x"ff",	--6176
		x"ff",	--6177
		x"ff",	--6178
		x"ff",	--6179
		x"ff",	--6180
		x"ff",	--6181
		x"ff",	--6182
		x"ff",	--6183
		x"ff",	--6184
		x"ff",	--6185
		x"ff",	--6186
		x"ff",	--6187
		x"ff",	--6188
		x"ff",	--6189
		x"ff",	--6190
		x"ff",	--6191
		x"ff",	--6192
		x"ff",	--6193
		x"ff",	--6194
		x"ff",	--6195
		x"ff",	--6196
		x"ff",	--6197
		x"ff",	--6198
		x"ff",	--6199
		x"ff",	--6200
		x"ff",	--6201
		x"ff",	--6202
		x"ff",	--6203
		x"ff",	--6204
		x"ff",	--6205
		x"ff",	--6206
		x"ff",	--6207
		x"ff",	--6208
		x"ff",	--6209
		x"ff",	--6210
		x"ff",	--6211
		x"ff",	--6212
		x"ff",	--6213
		x"ff",	--6214
		x"ff",	--6215
		x"ff",	--6216
		x"ff",	--6217
		x"ff",	--6218
		x"ff",	--6219
		x"ff",	--6220
		x"ff",	--6221
		x"ff",	--6222
		x"ff",	--6223
		x"ff",	--6224
		x"ff",	--6225
		x"ff",	--6226
		x"ff",	--6227
		x"ff",	--6228
		x"ff",	--6229
		x"ff",	--6230
		x"ff",	--6231
		x"ff",	--6232
		x"ff",	--6233
		x"ff",	--6234
		x"ff",	--6235
		x"ff",	--6236
		x"ff",	--6237
		x"ff",	--6238
		x"ff",	--6239
		x"ff",	--6240
		x"ff",	--6241
		x"ff",	--6242
		x"ff",	--6243
		x"ff",	--6244
		x"ff",	--6245
		x"ff",	--6246
		x"ff",	--6247
		x"ff",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"ff",	--6252
		x"ff",	--6253
		x"ff",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"c2",	--8176
		x"c2",	--8177
		x"c2",	--8178
		x"c2",	--8179
		x"c2",	--8180
		x"c2",	--8181
		x"c2",	--8182
		x"ce",	--8183
		x"ca",	--8184
		x"c2",	--8185
		x"c2",	--8186
		x"c2",	--8187
		x"c2",	--8188
		x"c2",	--8189
		x"c2",	--8190
		x"c0");	--8191

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
