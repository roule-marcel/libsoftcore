library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"e0",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"0a",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"e0",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"98",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"d6",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"e0",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"0a",	--29
		x"f9",	--30
		x"31",	--31
		x"be",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"12",	--44
		x"b0",	--45
		x"c8",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"de",	--50
		x"b0",	--51
		x"d6",	--52
		x"21",	--53
		x"3d",	--54
		x"fb",	--55
		x"3e",	--56
		x"7a",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"f8",	--61
		x"3d",	--62
		x"0c",	--63
		x"3e",	--64
		x"00",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"f8",	--69
		x"3d",	--70
		x"12",	--71
		x"3e",	--72
		x"74",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"f8",	--77
		x"3d",	--78
		x"17",	--79
		x"3e",	--80
		x"e2",	--81
		x"7f",	--82
		x"70",	--83
		x"b0",	--84
		x"f8",	--85
		x"3d",	--86
		x"1b",	--87
		x"3e",	--88
		x"e4",	--89
		x"7f",	--90
		x"65",	--91
		x"b0",	--92
		x"f8",	--93
		x"3d",	--94
		x"23",	--95
		x"3e",	--96
		x"78",	--97
		x"7f",	--98
		x"62",	--99
		x"b0",	--100
		x"f8",	--101
		x"0e",	--102
		x"0f",	--103
		x"b0",	--104
		x"8e",	--105
		x"2c",	--106
		x"3d",	--107
		x"20",	--108
		x"3e",	--109
		x"80",	--110
		x"0f",	--111
		x"3f",	--112
		x"0e",	--113
		x"b0",	--114
		x"9e",	--115
		x"0f",	--116
		x"3f",	--117
		x"0e",	--118
		x"b0",	--119
		x"e6",	--120
		x"2c",	--121
		x"3d",	--122
		x"20",	--123
		x"3e",	--124
		x"88",	--125
		x"0f",	--126
		x"2f",	--127
		x"b0",	--128
		x"9e",	--129
		x"0f",	--130
		x"2f",	--131
		x"b0",	--132
		x"e6",	--133
		x"0e",	--134
		x"2e",	--135
		x"0f",	--136
		x"3f",	--137
		x"0e",	--138
		x"b0",	--139
		x"d8",	--140
		x"3e",	--141
		x"98",	--142
		x"0f",	--143
		x"2f",	--144
		x"b0",	--145
		x"ec",	--146
		x"3e",	--147
		x"9c",	--148
		x"0f",	--149
		x"b0",	--150
		x"ec",	--151
		x"0e",	--152
		x"0f",	--153
		x"2f",	--154
		x"b0",	--155
		x"da",	--156
		x"b0",	--157
		x"c4",	--158
		x"0e",	--159
		x"3f",	--160
		x"8c",	--161
		x"b0",	--162
		x"d4",	--163
		x"0d",	--164
		x"1e",	--165
		x"b0",	--166
		x"18",	--167
		x"f2",	--168
		x"80",	--169
		x"19",	--170
		x"32",	--171
		x"0b",	--172
		x"b0",	--173
		x"30",	--174
		x"0f",	--175
		x"fc",	--176
		x"b0",	--177
		x"58",	--178
		x"7f",	--179
		x"15",	--180
		x"7f",	--181
		x"0d",	--182
		x"1b",	--183
		x"30",	--184
		x"2e",	--185
		x"b0",	--186
		x"d6",	--187
		x"21",	--188
		x"3f",	--189
		x"18",	--190
		x"0f",	--191
		x"0b",	--192
		x"cb",	--193
		x"00",	--194
		x"0e",	--195
		x"5f",	--196
		x"18",	--197
		x"b0",	--198
		x"2c",	--199
		x"0b",	--200
		x"e3",	--201
		x"0b",	--202
		x"e1",	--203
		x"3b",	--204
		x"30",	--205
		x"31",	--206
		x"b0",	--207
		x"d6",	--208
		x"21",	--209
		x"da",	--210
		x"3b",	--211
		x"28",	--212
		x"d7",	--213
		x"82",	--214
		x"0c",	--215
		x"0c",	--216
		x"4e",	--217
		x"8e",	--218
		x"0e",	--219
		x"30",	--220
		x"35",	--221
		x"81",	--222
		x"44",	--223
		x"b0",	--224
		x"d6",	--225
		x"21",	--226
		x"1f",	--227
		x"40",	--228
		x"3e",	--229
		x"18",	--230
		x"0e",	--231
		x"0e",	--232
		x"ce",	--233
		x"00",	--234
		x"1b",	--235
		x"c0",	--236
		x"30",	--237
		x"2c",	--238
		x"8f",	--239
		x"00",	--240
		x"8f",	--241
		x"02",	--242
		x"8f",	--243
		x"04",	--244
		x"8f",	--245
		x"06",	--246
		x"8f",	--247
		x"08",	--248
		x"8f",	--249
		x"0a",	--250
		x"30",	--251
		x"8f",	--252
		x"06",	--253
		x"8f",	--254
		x"08",	--255
		x"8f",	--256
		x"0a",	--257
		x"30",	--258
		x"8f",	--259
		x"00",	--260
		x"30",	--261
		x"8f",	--262
		x"02",	--263
		x"30",	--264
		x"8f",	--265
		x"04",	--266
		x"30",	--267
		x"8f",	--268
		x"06",	--269
		x"30",	--270
		x"1d",	--271
		x"06",	--272
		x"0d",	--273
		x"0e",	--274
		x"1d",	--275
		x"08",	--276
		x"8f",	--277
		x"08",	--278
		x"02",	--279
		x"32",	--280
		x"03",	--281
		x"82",	--282
		x"32",	--283
		x"a2",	--284
		x"38",	--285
		x"1c",	--286
		x"3a",	--287
		x"32",	--288
		x"02",	--289
		x"32",	--290
		x"03",	--291
		x"82",	--292
		x"32",	--293
		x"92",	--294
		x"02",	--295
		x"38",	--296
		x"1d",	--297
		x"3a",	--298
		x"32",	--299
		x"0d",	--300
		x"1e",	--301
		x"0a",	--302
		x"02",	--303
		x"32",	--304
		x"03",	--305
		x"82",	--306
		x"32",	--307
		x"92",	--308
		x"04",	--309
		x"38",	--310
		x"1f",	--311
		x"3a",	--312
		x"32",	--313
		x"0f",	--314
		x"30",	--315
		x"b2",	--316
		x"00",	--317
		x"92",	--318
		x"b2",	--319
		x"30",	--320
		x"94",	--321
		x"b2",	--322
		x"41",	--323
		x"96",	--324
		x"30",	--325
		x"34",	--326
		x"b0",	--327
		x"d6",	--328
		x"92",	--329
		x"90",	--330
		x"b1",	--331
		x"52",	--332
		x"00",	--333
		x"b0",	--334
		x"d6",	--335
		x"21",	--336
		x"0f",	--337
		x"30",	--338
		x"0b",	--339
		x"0a",	--340
		x"0a",	--341
		x"3b",	--342
		x"00",	--343
		x"0d",	--344
		x"0e",	--345
		x"1f",	--346
		x"1a",	--347
		x"b0",	--348
		x"3a",	--349
		x"0d",	--350
		x"0e",	--351
		x"1f",	--352
		x"18",	--353
		x"b0",	--354
		x"3a",	--355
		x"30",	--356
		x"6b",	--357
		x"b0",	--358
		x"d6",	--359
		x"21",	--360
		x"3a",	--361
		x"3b",	--362
		x"30",	--363
		x"82",	--364
		x"1a",	--365
		x"82",	--366
		x"18",	--367
		x"30",	--368
		x"0b",	--369
		x"0a",	--370
		x"21",	--371
		x"0a",	--372
		x"0b",	--373
		x"b2",	--374
		x"00",	--375
		x"47",	--376
		x"3a",	--377
		x"03",	--378
		x"4c",	--379
		x"37",	--380
		x"0e",	--381
		x"1f",	--382
		x"02",	--383
		x"b0",	--384
		x"d0",	--385
		x"0a",	--386
		x"0e",	--387
		x"1f",	--388
		x"04",	--389
		x"b0",	--390
		x"d0",	--391
		x"0b",	--392
		x"0f",	--393
		x"0a",	--394
		x"30",	--395
		x"b8",	--396
		x"b0",	--397
		x"d6",	--398
		x"31",	--399
		x"06",	--400
		x"0e",	--401
		x"0f",	--402
		x"b0",	--403
		x"4a",	--404
		x"0c",	--405
		x"3d",	--406
		x"c8",	--407
		x"b0",	--408
		x"1a",	--409
		x"0d",	--410
		x"0e",	--411
		x"1f",	--412
		x"1a",	--413
		x"b0",	--414
		x"3a",	--415
		x"0e",	--416
		x"0f",	--417
		x"b0",	--418
		x"4a",	--419
		x"0c",	--420
		x"3d",	--421
		x"c8",	--422
		x"b0",	--423
		x"1a",	--424
		x"0d",	--425
		x"0e",	--426
		x"1f",	--427
		x"18",	--428
		x"b0",	--429
		x"3a",	--430
		x"0f",	--431
		x"21",	--432
		x"3a",	--433
		x"3b",	--434
		x"30",	--435
		x"0e",	--436
		x"1f",	--437
		x"06",	--438
		x"b0",	--439
		x"d0",	--440
		x"1d",	--441
		x"0e",	--442
		x"1f",	--443
		x"00",	--444
		x"b0",	--445
		x"18",	--446
		x"bd",	--447
		x"0e",	--448
		x"3f",	--449
		x"a6",	--450
		x"b0",	--451
		x"d4",	--452
		x"82",	--453
		x"00",	--454
		x"b1",	--455
		x"30",	--456
		x"72",	--457
		x"b0",	--458
		x"d6",	--459
		x"b1",	--460
		x"8c",	--461
		x"00",	--462
		x"b0",	--463
		x"d6",	--464
		x"a1",	--465
		x"00",	--466
		x"30",	--467
		x"9d",	--468
		x"b0",	--469
		x"d6",	--470
		x"21",	--471
		x"3f",	--472
		x"d6",	--473
		x"1f",	--474
		x"1e",	--475
		x"2e",	--476
		x"1f",	--477
		x"1c",	--478
		x"2f",	--479
		x"2e",	--480
		x"1e",	--481
		x"02",	--482
		x"2f",	--483
		x"1f",	--484
		x"02",	--485
		x"30",	--486
		x"c0",	--487
		x"b0",	--488
		x"d6",	--489
		x"31",	--490
		x"0a",	--491
		x"30",	--492
		x"82",	--493
		x"1c",	--494
		x"82",	--495
		x"1e",	--496
		x"30",	--497
		x"0b",	--498
		x"0a",	--499
		x"09",	--500
		x"21",	--501
		x"0a",	--502
		x"0b",	--503
		x"81",	--504
		x"00",	--505
		x"1f",	--506
		x"1a",	--507
		x"b2",	--508
		x"02",	--509
		x"36",	--510
		x"92",	--511
		x"0a",	--512
		x"0e",	--513
		x"1f",	--514
		x"02",	--515
		x"b0",	--516
		x"d0",	--517
		x"09",	--518
		x"3a",	--519
		x"03",	--520
		x"1b",	--521
		x"0d",	--522
		x"0e",	--523
		x"1f",	--524
		x"02",	--525
		x"b0",	--526
		x"18",	--527
		x"0f",	--528
		x"21",	--529
		x"39",	--530
		x"3a",	--531
		x"3b",	--532
		x"30",	--533
		x"82",	--534
		x"0a",	--535
		x"13",	--536
		x"82",	--537
		x"0a",	--538
		x"1f",	--539
		x"02",	--540
		x"b0",	--541
		x"40",	--542
		x"0f",	--543
		x"21",	--544
		x"39",	--545
		x"3a",	--546
		x"3b",	--547
		x"30",	--548
		x"0e",	--549
		x"1f",	--550
		x"04",	--551
		x"b0",	--552
		x"d0",	--553
		x"0d",	--554
		x"df",	--555
		x"0f",	--556
		x"b0",	--557
		x"b4",	--558
		x"0f",	--559
		x"21",	--560
		x"39",	--561
		x"3a",	--562
		x"3b",	--563
		x"30",	--564
		x"0e",	--565
		x"3f",	--566
		x"b4",	--567
		x"b0",	--568
		x"d4",	--569
		x"82",	--570
		x"02",	--571
		x"c2",	--572
		x"1f",	--573
		x"82",	--574
		x"0c",	--575
		x"01",	--576
		x"0f",	--577
		x"82",	--578
		x"0c",	--579
		x"0f",	--580
		x"30",	--581
		x"1e",	--582
		x"0e",	--583
		x"3e",	--584
		x"06",	--585
		x"0f",	--586
		x"0f",	--587
		x"10",	--588
		x"ce",	--589
		x"c2",	--590
		x"19",	--591
		x"3e",	--592
		x"07",	--593
		x"03",	--594
		x"82",	--595
		x"0e",	--596
		x"30",	--597
		x"1e",	--598
		x"82",	--599
		x"0e",	--600
		x"30",	--601
		x"f2",	--602
		x"0e",	--603
		x"19",	--604
		x"f2",	--605
		x"f2",	--606
		x"0a",	--607
		x"19",	--608
		x"ee",	--609
		x"e2",	--610
		x"19",	--611
		x"eb",	--612
		x"f2",	--613
		x"0d",	--614
		x"19",	--615
		x"e7",	--616
		x"f2",	--617
		x"09",	--618
		x"19",	--619
		x"e3",	--620
		x"f2",	--621
		x"03",	--622
		x"19",	--623
		x"df",	--624
		x"f2",	--625
		x"07",	--626
		x"19",	--627
		x"db",	--628
		x"5e",	--629
		x"19",	--630
		x"4e",	--631
		x"0f",	--632
		x"03",	--633
		x"c2",	--634
		x"19",	--635
		x"30",	--636
		x"c2",	--637
		x"19",	--638
		x"30",	--639
		x"0b",	--640
		x"0a",	--641
		x"21",	--642
		x"0a",	--643
		x"0b",	--644
		x"30",	--645
		x"38",	--646
		x"b0",	--647
		x"d6",	--648
		x"21",	--649
		x"3a",	--650
		x"03",	--651
		x"1b",	--652
		x"0e",	--653
		x"1f",	--654
		x"02",	--655
		x"b0",	--656
		x"d0",	--657
		x"0a",	--658
		x"0e",	--659
		x"1f",	--660
		x"04",	--661
		x"b0",	--662
		x"d0",	--663
		x"0b",	--664
		x"0f",	--665
		x"0a",	--666
		x"30",	--667
		x"80",	--668
		x"b0",	--669
		x"d6",	--670
		x"31",	--671
		x"06",	--672
		x"8a",	--673
		x"00",	--674
		x"0f",	--675
		x"21",	--676
		x"3a",	--677
		x"3b",	--678
		x"30",	--679
		x"30",	--680
		x"40",	--681
		x"b0",	--682
		x"d6",	--683
		x"b1",	--684
		x"5a",	--685
		x"00",	--686
		x"b0",	--687
		x"d6",	--688
		x"a1",	--689
		x"00",	--690
		x"30",	--691
		x"6b",	--692
		x"b0",	--693
		x"d6",	--694
		x"21",	--695
		x"3f",	--696
		x"ea",	--697
		x"0b",	--698
		x"21",	--699
		x"0b",	--700
		x"1f",	--701
		x"17",	--702
		x"16",	--703
		x"30",	--704
		x"9b",	--705
		x"b0",	--706
		x"d6",	--707
		x"21",	--708
		x"0e",	--709
		x"1f",	--710
		x"02",	--711
		x"b0",	--712
		x"d0",	--713
		x"2f",	--714
		x"0f",	--715
		x"30",	--716
		x"80",	--717
		x"b0",	--718
		x"d6",	--719
		x"31",	--720
		x"06",	--721
		x"0f",	--722
		x"21",	--723
		x"3b",	--724
		x"30",	--725
		x"30",	--726
		x"40",	--727
		x"b0",	--728
		x"d6",	--729
		x"b1",	--730
		x"5a",	--731
		x"00",	--732
		x"b0",	--733
		x"d6",	--734
		x"a1",	--735
		x"00",	--736
		x"30",	--737
		x"8c",	--738
		x"b0",	--739
		x"d6",	--740
		x"21",	--741
		x"3f",	--742
		x"eb",	--743
		x"0b",	--744
		x"0a",	--745
		x"8e",	--746
		x"00",	--747
		x"6d",	--748
		x"4d",	--749
		x"5e",	--750
		x"1f",	--751
		x"0a",	--752
		x"0c",	--753
		x"0f",	--754
		x"7b",	--755
		x"0a",	--756
		x"2b",	--757
		x"0c",	--758
		x"0c",	--759
		x"0c",	--760
		x"0c",	--761
		x"8d",	--762
		x"0c",	--763
		x"3c",	--764
		x"d0",	--765
		x"1a",	--766
		x"7d",	--767
		x"4d",	--768
		x"17",	--769
		x"7d",	--770
		x"78",	--771
		x"1a",	--772
		x"4b",	--773
		x"7b",	--774
		x"d0",	--775
		x"0a",	--776
		x"e9",	--777
		x"7b",	--778
		x"0a",	--779
		x"34",	--780
		x"0c",	--781
		x"0b",	--782
		x"0b",	--783
		x"0b",	--784
		x"0c",	--785
		x"8d",	--786
		x"0c",	--787
		x"3c",	--788
		x"d0",	--789
		x"7d",	--790
		x"4d",	--791
		x"e9",	--792
		x"9e",	--793
		x"00",	--794
		x"0f",	--795
		x"3a",	--796
		x"3b",	--797
		x"30",	--798
		x"1a",	--799
		x"de",	--800
		x"4b",	--801
		x"7b",	--802
		x"9f",	--803
		x"7b",	--804
		x"06",	--805
		x"0a",	--806
		x"0c",	--807
		x"0c",	--808
		x"0c",	--809
		x"0c",	--810
		x"8d",	--811
		x"0c",	--812
		x"3c",	--813
		x"a9",	--814
		x"1a",	--815
		x"ce",	--816
		x"4b",	--817
		x"7b",	--818
		x"bf",	--819
		x"7b",	--820
		x"06",	--821
		x"0a",	--822
		x"0c",	--823
		x"0c",	--824
		x"0c",	--825
		x"0c",	--826
		x"8d",	--827
		x"0c",	--828
		x"3c",	--829
		x"c9",	--830
		x"1a",	--831
		x"be",	--832
		x"8d",	--833
		x"0d",	--834
		x"30",	--835
		x"a2",	--836
		x"b0",	--837
		x"d6",	--838
		x"21",	--839
		x"0c",	--840
		x"0f",	--841
		x"3a",	--842
		x"3b",	--843
		x"30",	--844
		x"0c",	--845
		x"ca",	--846
		x"0b",	--847
		x"0a",	--848
		x"0b",	--849
		x"0a",	--850
		x"8f",	--851
		x"00",	--852
		x"8f",	--853
		x"02",	--854
		x"8f",	--855
		x"04",	--856
		x"0c",	--857
		x"0d",	--858
		x"3e",	--859
		x"00",	--860
		x"3f",	--861
		x"6e",	--862
		x"b0",	--863
		x"be",	--864
		x"8b",	--865
		x"02",	--866
		x"02",	--867
		x"32",	--868
		x"03",	--869
		x"82",	--870
		x"32",	--871
		x"b2",	--872
		x"18",	--873
		x"38",	--874
		x"9b",	--875
		x"3a",	--876
		x"06",	--877
		x"32",	--878
		x"0f",	--879
		x"3a",	--880
		x"3b",	--881
		x"30",	--882
		x"0b",	--883
		x"09",	--884
		x"08",	--885
		x"8f",	--886
		x"06",	--887
		x"bf",	--888
		x"00",	--889
		x"08",	--890
		x"2b",	--891
		x"1e",	--892
		x"02",	--893
		x"0f",	--894
		x"b0",	--895
		x"4a",	--896
		x"0c",	--897
		x"3d",	--898
		x"00",	--899
		x"b0",	--900
		x"f6",	--901
		x"08",	--902
		x"09",	--903
		x"1e",	--904
		x"06",	--905
		x"0f",	--906
		x"b0",	--907
		x"4a",	--908
		x"0c",	--909
		x"0d",	--910
		x"0e",	--911
		x"0f",	--912
		x"b0",	--913
		x"a6",	--914
		x"b0",	--915
		x"86",	--916
		x"8b",	--917
		x"04",	--918
		x"9b",	--919
		x"00",	--920
		x"38",	--921
		x"39",	--922
		x"3b",	--923
		x"30",	--924
		x"0b",	--925
		x"0a",	--926
		x"09",	--927
		x"0a",	--928
		x"0b",	--929
		x"8f",	--930
		x"06",	--931
		x"8f",	--932
		x"08",	--933
		x"29",	--934
		x"1e",	--935
		x"02",	--936
		x"0f",	--937
		x"b0",	--938
		x"4a",	--939
		x"0c",	--940
		x"0d",	--941
		x"0e",	--942
		x"0f",	--943
		x"b0",	--944
		x"f6",	--945
		x"0a",	--946
		x"0b",	--947
		x"1e",	--948
		x"06",	--949
		x"0f",	--950
		x"b0",	--951
		x"4a",	--952
		x"0c",	--953
		x"0d",	--954
		x"0e",	--955
		x"0f",	--956
		x"b0",	--957
		x"a6",	--958
		x"b0",	--959
		x"86",	--960
		x"89",	--961
		x"04",	--962
		x"39",	--963
		x"3a",	--964
		x"3b",	--965
		x"30",	--966
		x"0b",	--967
		x"0a",	--968
		x"92",	--969
		x"10",	--970
		x"14",	--971
		x"3b",	--972
		x"24",	--973
		x"0a",	--974
		x"2b",	--975
		x"5f",	--976
		x"fc",	--977
		x"8f",	--978
		x"0f",	--979
		x"30",	--980
		x"b7",	--981
		x"b0",	--982
		x"d6",	--983
		x"31",	--984
		x"06",	--985
		x"1a",	--986
		x"3b",	--987
		x"06",	--988
		x"1a",	--989
		x"10",	--990
		x"ef",	--991
		x"0f",	--992
		x"3a",	--993
		x"3b",	--994
		x"30",	--995
		x"1e",	--996
		x"10",	--997
		x"3e",	--998
		x"20",	--999
		x"12",	--1000
		x"0f",	--1001
		x"0f",	--1002
		x"0f",	--1003
		x"0f",	--1004
		x"3f",	--1005
		x"20",	--1006
		x"ff",	--1007
		x"68",	--1008
		x"00",	--1009
		x"bf",	--1010
		x"8e",	--1011
		x"02",	--1012
		x"bf",	--1013
		x"04",	--1014
		x"04",	--1015
		x"1e",	--1016
		x"82",	--1017
		x"10",	--1018
		x"30",	--1019
		x"0b",	--1020
		x"1b",	--1021
		x"10",	--1022
		x"3b",	--1023
		x"20",	--1024
		x"12",	--1025
		x"0c",	--1026
		x"0c",	--1027
		x"0c",	--1028
		x"0c",	--1029
		x"3c",	--1030
		x"20",	--1031
		x"cc",	--1032
		x"00",	--1033
		x"8c",	--1034
		x"02",	--1035
		x"8c",	--1036
		x"04",	--1037
		x"1b",	--1038
		x"82",	--1039
		x"10",	--1040
		x"0f",	--1041
		x"3b",	--1042
		x"30",	--1043
		x"3f",	--1044
		x"fc",	--1045
		x"0b",	--1046
		x"31",	--1047
		x"f0",	--1048
		x"1b",	--1049
		x"10",	--1050
		x"1b",	--1051
		x"0f",	--1052
		x"5f",	--1053
		x"20",	--1054
		x"16",	--1055
		x"3d",	--1056
		x"26",	--1057
		x"0c",	--1058
		x"05",	--1059
		x"3d",	--1060
		x"06",	--1061
		x"cd",	--1062
		x"fa",	--1063
		x"0e",	--1064
		x"1c",	--1065
		x"0c",	--1066
		x"f8",	--1067
		x"30",	--1068
		x"bf",	--1069
		x"b0",	--1070
		x"d6",	--1071
		x"21",	--1072
		x"3f",	--1073
		x"31",	--1074
		x"10",	--1075
		x"3b",	--1076
		x"30",	--1077
		x"0c",	--1078
		x"81",	--1079
		x"00",	--1080
		x"6d",	--1081
		x"4d",	--1082
		x"24",	--1083
		x"1e",	--1084
		x"1f",	--1085
		x"06",	--1086
		x"6d",	--1087
		x"4d",	--1088
		x"11",	--1089
		x"1e",	--1090
		x"3f",	--1091
		x"0e",	--1092
		x"7d",	--1093
		x"20",	--1094
		x"f7",	--1095
		x"ce",	--1096
		x"ff",	--1097
		x"0d",	--1098
		x"0d",	--1099
		x"0d",	--1100
		x"8d",	--1101
		x"00",	--1102
		x"1f",	--1103
		x"6d",	--1104
		x"4d",	--1105
		x"ef",	--1106
		x"0e",	--1107
		x"0e",	--1108
		x"0c",	--1109
		x"0c",	--1110
		x"3c",	--1111
		x"20",	--1112
		x"0e",	--1113
		x"9c",	--1114
		x"02",	--1115
		x"31",	--1116
		x"10",	--1117
		x"3b",	--1118
		x"30",	--1119
		x"1f",	--1120
		x"f1",	--1121
		x"b2",	--1122
		x"d2",	--1123
		x"60",	--1124
		x"b2",	--1125
		x"b8",	--1126
		x"72",	--1127
		x"0f",	--1128
		x"30",	--1129
		x"0b",	--1130
		x"0b",	--1131
		x"1f",	--1132
		x"12",	--1133
		x"3f",	--1134
		x"20",	--1135
		x"19",	--1136
		x"0c",	--1137
		x"0c",	--1138
		x"0d",	--1139
		x"0d",	--1140
		x"0d",	--1141
		x"0d",	--1142
		x"0d",	--1143
		x"3d",	--1144
		x"e0",	--1145
		x"8d",	--1146
		x"00",	--1147
		x"8d",	--1148
		x"02",	--1149
		x"8d",	--1150
		x"08",	--1151
		x"8d",	--1152
		x"0a",	--1153
		x"8d",	--1154
		x"0c",	--1155
		x"0e",	--1156
		x"1e",	--1157
		x"82",	--1158
		x"12",	--1159
		x"3b",	--1160
		x"30",	--1161
		x"3f",	--1162
		x"fc",	--1163
		x"0f",	--1164
		x"0c",	--1165
		x"0c",	--1166
		x"0c",	--1167
		x"0c",	--1168
		x"0c",	--1169
		x"3c",	--1170
		x"e0",	--1171
		x"8c",	--1172
		x"02",	--1173
		x"8c",	--1174
		x"04",	--1175
		x"8c",	--1176
		x"06",	--1177
		x"8c",	--1178
		x"08",	--1179
		x"9c",	--1180
		x"00",	--1181
		x"0f",	--1182
		x"30",	--1183
		x"0f",	--1184
		x"0e",	--1185
		x"0e",	--1186
		x"0e",	--1187
		x"0e",	--1188
		x"0e",	--1189
		x"8e",	--1190
		x"e0",	--1191
		x"0f",	--1192
		x"30",	--1193
		x"0f",	--1194
		x"0e",	--1195
		x"0d",	--1196
		x"0c",	--1197
		x"0b",	--1198
		x"0a",	--1199
		x"09",	--1200
		x"08",	--1201
		x"07",	--1202
		x"92",	--1203
		x"12",	--1204
		x"33",	--1205
		x"3a",	--1206
		x"e0",	--1207
		x"0b",	--1208
		x"2b",	--1209
		x"08",	--1210
		x"38",	--1211
		x"07",	--1212
		x"37",	--1213
		x"06",	--1214
		x"09",	--1215
		x"0f",	--1216
		x"1f",	--1217
		x"8b",	--1218
		x"00",	--1219
		x"19",	--1220
		x"3a",	--1221
		x"0e",	--1222
		x"3b",	--1223
		x"0e",	--1224
		x"38",	--1225
		x"0e",	--1226
		x"37",	--1227
		x"0e",	--1228
		x"19",	--1229
		x"12",	--1230
		x"19",	--1231
		x"8a",	--1232
		x"00",	--1233
		x"f1",	--1234
		x"2f",	--1235
		x"1f",	--1236
		x"02",	--1237
		x"ea",	--1238
		x"8b",	--1239
		x"00",	--1240
		x"1f",	--1241
		x"0a",	--1242
		x"9b",	--1243
		x"08",	--1244
		x"88",	--1245
		x"00",	--1246
		x"e4",	--1247
		x"2f",	--1248
		x"1f",	--1249
		x"87",	--1250
		x"00",	--1251
		x"2f",	--1252
		x"de",	--1253
		x"8a",	--1254
		x"00",	--1255
		x"db",	--1256
		x"b2",	--1257
		x"fe",	--1258
		x"60",	--1259
		x"37",	--1260
		x"38",	--1261
		x"39",	--1262
		x"3a",	--1263
		x"3b",	--1264
		x"3c",	--1265
		x"3d",	--1266
		x"3e",	--1267
		x"3f",	--1268
		x"00",	--1269
		x"8f",	--1270
		x"00",	--1271
		x"0f",	--1272
		x"30",	--1273
		x"2f",	--1274
		x"2f",	--1275
		x"30",	--1276
		x"5e",	--1277
		x"81",	--1278
		x"3e",	--1279
		x"fc",	--1280
		x"c2",	--1281
		x"84",	--1282
		x"0f",	--1283
		x"30",	--1284
		x"3f",	--1285
		x"0f",	--1286
		x"5f",	--1287
		x"7e",	--1288
		x"8f",	--1289
		x"b0",	--1290
		x"fa",	--1291
		x"30",	--1292
		x"0b",	--1293
		x"0b",	--1294
		x"0e",	--1295
		x"0e",	--1296
		x"0e",	--1297
		x"0e",	--1298
		x"0e",	--1299
		x"0f",	--1300
		x"b0",	--1301
		x"0a",	--1302
		x"0f",	--1303
		x"b0",	--1304
		x"0a",	--1305
		x"3b",	--1306
		x"30",	--1307
		x"0b",	--1308
		x"0a",	--1309
		x"0a",	--1310
		x"3b",	--1311
		x"07",	--1312
		x"0e",	--1313
		x"4d",	--1314
		x"7d",	--1315
		x"0f",	--1316
		x"03",	--1317
		x"0e",	--1318
		x"7d",	--1319
		x"fd",	--1320
		x"1e",	--1321
		x"0a",	--1322
		x"3f",	--1323
		x"31",	--1324
		x"b0",	--1325
		x"fa",	--1326
		x"3b",	--1327
		x"3b",	--1328
		x"ef",	--1329
		x"3a",	--1330
		x"3b",	--1331
		x"30",	--1332
		x"3f",	--1333
		x"30",	--1334
		x"f5",	--1335
		x"0b",	--1336
		x"0b",	--1337
		x"0e",	--1338
		x"8e",	--1339
		x"8e",	--1340
		x"0f",	--1341
		x"b0",	--1342
		x"1a",	--1343
		x"0f",	--1344
		x"b0",	--1345
		x"1a",	--1346
		x"3b",	--1347
		x"30",	--1348
		x"0b",	--1349
		x"0a",	--1350
		x"0a",	--1351
		x"0b",	--1352
		x"0d",	--1353
		x"8d",	--1354
		x"8d",	--1355
		x"0f",	--1356
		x"b0",	--1357
		x"1a",	--1358
		x"0f",	--1359
		x"b0",	--1360
		x"1a",	--1361
		x"0c",	--1362
		x"0d",	--1363
		x"8d",	--1364
		x"8c",	--1365
		x"4d",	--1366
		x"0d",	--1367
		x"0f",	--1368
		x"b0",	--1369
		x"1a",	--1370
		x"0f",	--1371
		x"b0",	--1372
		x"1a",	--1373
		x"3a",	--1374
		x"3b",	--1375
		x"30",	--1376
		x"0b",	--1377
		x"0a",	--1378
		x"09",	--1379
		x"0a",	--1380
		x"0e",	--1381
		x"19",	--1382
		x"09",	--1383
		x"39",	--1384
		x"0b",	--1385
		x"0d",	--1386
		x"0d",	--1387
		x"6f",	--1388
		x"8f",	--1389
		x"b0",	--1390
		x"1a",	--1391
		x"0b",	--1392
		x"0e",	--1393
		x"1b",	--1394
		x"3b",	--1395
		x"07",	--1396
		x"05",	--1397
		x"3f",	--1398
		x"20",	--1399
		x"b0",	--1400
		x"fa",	--1401
		x"ef",	--1402
		x"3f",	--1403
		x"3a",	--1404
		x"b0",	--1405
		x"fa",	--1406
		x"ea",	--1407
		x"39",	--1408
		x"3a",	--1409
		x"3b",	--1410
		x"30",	--1411
		x"0b",	--1412
		x"0a",	--1413
		x"09",	--1414
		x"0a",	--1415
		x"0e",	--1416
		x"17",	--1417
		x"09",	--1418
		x"39",	--1419
		x"0b",	--1420
		x"6f",	--1421
		x"8f",	--1422
		x"b0",	--1423
		x"0a",	--1424
		x"0b",	--1425
		x"0e",	--1426
		x"1b",	--1427
		x"3b",	--1428
		x"07",	--1429
		x"f6",	--1430
		x"3f",	--1431
		x"20",	--1432
		x"b0",	--1433
		x"fa",	--1434
		x"6f",	--1435
		x"8f",	--1436
		x"b0",	--1437
		x"0a",	--1438
		x"0b",	--1439
		x"f2",	--1440
		x"39",	--1441
		x"3a",	--1442
		x"3b",	--1443
		x"30",	--1444
		x"0b",	--1445
		x"0a",	--1446
		x"09",	--1447
		x"31",	--1448
		x"ec",	--1449
		x"0b",	--1450
		x"0f",	--1451
		x"34",	--1452
		x"3b",	--1453
		x"0a",	--1454
		x"38",	--1455
		x"09",	--1456
		x"0a",	--1457
		x"0a",	--1458
		x"3e",	--1459
		x"0a",	--1460
		x"0f",	--1461
		x"b0",	--1462
		x"76",	--1463
		x"7f",	--1464
		x"30",	--1465
		x"ca",	--1466
		x"00",	--1467
		x"19",	--1468
		x"3e",	--1469
		x"0a",	--1470
		x"0f",	--1471
		x"b0",	--1472
		x"44",	--1473
		x"0b",	--1474
		x"3f",	--1475
		x"0a",	--1476
		x"eb",	--1477
		x"0a",	--1478
		x"1a",	--1479
		x"09",	--1480
		x"3e",	--1481
		x"0a",	--1482
		x"0f",	--1483
		x"b0",	--1484
		x"76",	--1485
		x"7f",	--1486
		x"30",	--1487
		x"c9",	--1488
		x"00",	--1489
		x"3a",	--1490
		x"0f",	--1491
		x"0f",	--1492
		x"6f",	--1493
		x"8f",	--1494
		x"b0",	--1495
		x"fa",	--1496
		x"0a",	--1497
		x"f7",	--1498
		x"31",	--1499
		x"14",	--1500
		x"39",	--1501
		x"3a",	--1502
		x"3b",	--1503
		x"30",	--1504
		x"3f",	--1505
		x"2d",	--1506
		x"b0",	--1507
		x"fa",	--1508
		x"3b",	--1509
		x"1b",	--1510
		x"c5",	--1511
		x"1a",	--1512
		x"09",	--1513
		x"dd",	--1514
		x"0b",	--1515
		x"0a",	--1516
		x"09",	--1517
		x"0b",	--1518
		x"3b",	--1519
		x"39",	--1520
		x"6f",	--1521
		x"4f",	--1522
		x"0b",	--1523
		x"1a",	--1524
		x"8f",	--1525
		x"b0",	--1526
		x"fa",	--1527
		x"0a",	--1528
		x"09",	--1529
		x"19",	--1530
		x"5f",	--1531
		x"01",	--1532
		x"4f",	--1533
		x"10",	--1534
		x"7f",	--1535
		x"25",	--1536
		x"f3",	--1537
		x"0a",	--1538
		x"1a",	--1539
		x"5f",	--1540
		x"01",	--1541
		x"7f",	--1542
		x"db",	--1543
		x"7f",	--1544
		x"54",	--1545
		x"ee",	--1546
		x"4f",	--1547
		x"0f",	--1548
		x"10",	--1549
		x"d6",	--1550
		x"39",	--1551
		x"3a",	--1552
		x"3b",	--1553
		x"30",	--1554
		x"09",	--1555
		x"29",	--1556
		x"1e",	--1557
		x"02",	--1558
		x"2f",	--1559
		x"b0",	--1560
		x"c2",	--1561
		x"0b",	--1562
		x"dd",	--1563
		x"09",	--1564
		x"29",	--1565
		x"2f",	--1566
		x"b0",	--1567
		x"70",	--1568
		x"0b",	--1569
		x"d6",	--1570
		x"0f",	--1571
		x"2b",	--1572
		x"29",	--1573
		x"6f",	--1574
		x"4f",	--1575
		x"d0",	--1576
		x"19",	--1577
		x"8f",	--1578
		x"b0",	--1579
		x"fa",	--1580
		x"7f",	--1581
		x"4f",	--1582
		x"fa",	--1583
		x"c8",	--1584
		x"09",	--1585
		x"29",	--1586
		x"1e",	--1587
		x"02",	--1588
		x"2f",	--1589
		x"b0",	--1590
		x"08",	--1591
		x"0b",	--1592
		x"bf",	--1593
		x"09",	--1594
		x"29",	--1595
		x"2e",	--1596
		x"0f",	--1597
		x"8f",	--1598
		x"8f",	--1599
		x"8f",	--1600
		x"8f",	--1601
		x"b0",	--1602
		x"8a",	--1603
		x"0b",	--1604
		x"b3",	--1605
		x"09",	--1606
		x"29",	--1607
		x"2f",	--1608
		x"b0",	--1609
		x"4a",	--1610
		x"0b",	--1611
		x"ac",	--1612
		x"09",	--1613
		x"29",	--1614
		x"2f",	--1615
		x"b0",	--1616
		x"fa",	--1617
		x"0b",	--1618
		x"a5",	--1619
		x"09",	--1620
		x"29",	--1621
		x"2f",	--1622
		x"b0",	--1623
		x"1a",	--1624
		x"0b",	--1625
		x"9e",	--1626
		x"09",	--1627
		x"29",	--1628
		x"2f",	--1629
		x"b0",	--1630
		x"38",	--1631
		x"0b",	--1632
		x"97",	--1633
		x"3f",	--1634
		x"25",	--1635
		x"b0",	--1636
		x"fa",	--1637
		x"92",	--1638
		x"0f",	--1639
		x"0e",	--1640
		x"1f",	--1641
		x"14",	--1642
		x"df",	--1643
		x"85",	--1644
		x"a0",	--1645
		x"1f",	--1646
		x"14",	--1647
		x"3f",	--1648
		x"3f",	--1649
		x"13",	--1650
		x"92",	--1651
		x"14",	--1652
		x"1e",	--1653
		x"14",	--1654
		x"1f",	--1655
		x"16",	--1656
		x"0e",	--1657
		x"02",	--1658
		x"92",	--1659
		x"16",	--1660
		x"f2",	--1661
		x"10",	--1662
		x"81",	--1663
		x"3e",	--1664
		x"3f",	--1665
		x"b1",	--1666
		x"f0",	--1667
		x"00",	--1668
		x"00",	--1669
		x"82",	--1670
		x"14",	--1671
		x"ec",	--1672
		x"0c",	--1673
		x"0d",	--1674
		x"3e",	--1675
		x"00",	--1676
		x"3f",	--1677
		x"6e",	--1678
		x"b0",	--1679
		x"7e",	--1680
		x"3e",	--1681
		x"82",	--1682
		x"82",	--1683
		x"f2",	--1684
		x"11",	--1685
		x"80",	--1686
		x"30",	--1687
		x"1e",	--1688
		x"14",	--1689
		x"1f",	--1690
		x"16",	--1691
		x"0e",	--1692
		x"05",	--1693
		x"1f",	--1694
		x"14",	--1695
		x"1f",	--1696
		x"16",	--1697
		x"30",	--1698
		x"1d",	--1699
		x"14",	--1700
		x"1e",	--1701
		x"16",	--1702
		x"3f",	--1703
		x"40",	--1704
		x"0f",	--1705
		x"0f",	--1706
		x"30",	--1707
		x"1f",	--1708
		x"16",	--1709
		x"5f",	--1710
		x"a0",	--1711
		x"1d",	--1712
		x"16",	--1713
		x"1e",	--1714
		x"14",	--1715
		x"0d",	--1716
		x"0b",	--1717
		x"1e",	--1718
		x"16",	--1719
		x"3e",	--1720
		x"3f",	--1721
		x"03",	--1722
		x"82",	--1723
		x"16",	--1724
		x"30",	--1725
		x"92",	--1726
		x"16",	--1727
		x"30",	--1728
		x"4f",	--1729
		x"30",	--1730
		x"0b",	--1731
		x"0a",	--1732
		x"0a",	--1733
		x"0b",	--1734
		x"0c",	--1735
		x"3d",	--1736
		x"00",	--1737
		x"b0",	--1738
		x"6a",	--1739
		x"0f",	--1740
		x"07",	--1741
		x"0e",	--1742
		x"0f",	--1743
		x"b0",	--1744
		x"ba",	--1745
		x"3a",	--1746
		x"3b",	--1747
		x"30",	--1748
		x"0c",	--1749
		x"3d",	--1750
		x"00",	--1751
		x"0e",	--1752
		x"0f",	--1753
		x"b0",	--1754
		x"a6",	--1755
		x"b0",	--1756
		x"ba",	--1757
		x"0e",	--1758
		x"3f",	--1759
		x"00",	--1760
		x"3a",	--1761
		x"3b",	--1762
		x"30",	--1763
		x"0b",	--1764
		x"0a",	--1765
		x"09",	--1766
		x"08",	--1767
		x"07",	--1768
		x"06",	--1769
		x"05",	--1770
		x"04",	--1771
		x"31",	--1772
		x"fa",	--1773
		x"08",	--1774
		x"6b",	--1775
		x"6b",	--1776
		x"67",	--1777
		x"6c",	--1778
		x"6c",	--1779
		x"e9",	--1780
		x"6b",	--1781
		x"02",	--1782
		x"30",	--1783
		x"48",	--1784
		x"6c",	--1785
		x"e3",	--1786
		x"6c",	--1787
		x"bb",	--1788
		x"6b",	--1789
		x"df",	--1790
		x"91",	--1791
		x"02",	--1792
		x"00",	--1793
		x"1b",	--1794
		x"02",	--1795
		x"14",	--1796
		x"04",	--1797
		x"15",	--1798
		x"06",	--1799
		x"16",	--1800
		x"04",	--1801
		x"17",	--1802
		x"06",	--1803
		x"2c",	--1804
		x"0c",	--1805
		x"09",	--1806
		x"0c",	--1807
		x"bf",	--1808
		x"39",	--1809
		x"20",	--1810
		x"50",	--1811
		x"1c",	--1812
		x"d7",	--1813
		x"81",	--1814
		x"02",	--1815
		x"81",	--1816
		x"04",	--1817
		x"4c",	--1818
		x"7c",	--1819
		x"1f",	--1820
		x"0b",	--1821
		x"0a",	--1822
		x"0b",	--1823
		x"12",	--1824
		x"0b",	--1825
		x"0a",	--1826
		x"7c",	--1827
		x"fb",	--1828
		x"81",	--1829
		x"02",	--1830
		x"81",	--1831
		x"04",	--1832
		x"1c",	--1833
		x"0d",	--1834
		x"79",	--1835
		x"1f",	--1836
		x"04",	--1837
		x"0c",	--1838
		x"0d",	--1839
		x"79",	--1840
		x"fc",	--1841
		x"3c",	--1842
		x"3d",	--1843
		x"0c",	--1844
		x"0d",	--1845
		x"1a",	--1846
		x"0b",	--1847
		x"0c",	--1848
		x"02",	--1849
		x"0d",	--1850
		x"e5",	--1851
		x"16",	--1852
		x"02",	--1853
		x"17",	--1854
		x"04",	--1855
		x"06",	--1856
		x"07",	--1857
		x"5f",	--1858
		x"01",	--1859
		x"5f",	--1860
		x"01",	--1861
		x"28",	--1862
		x"c8",	--1863
		x"01",	--1864
		x"a8",	--1865
		x"02",	--1866
		x"0e",	--1867
		x"0f",	--1868
		x"0e",	--1869
		x"0f",	--1870
		x"88",	--1871
		x"04",	--1872
		x"88",	--1873
		x"06",	--1874
		x"f8",	--1875
		x"03",	--1876
		x"00",	--1877
		x"0f",	--1878
		x"4d",	--1879
		x"0f",	--1880
		x"31",	--1881
		x"06",	--1882
		x"34",	--1883
		x"35",	--1884
		x"36",	--1885
		x"37",	--1886
		x"38",	--1887
		x"39",	--1888
		x"3a",	--1889
		x"3b",	--1890
		x"30",	--1891
		x"2b",	--1892
		x"67",	--1893
		x"81",	--1894
		x"00",	--1895
		x"04",	--1896
		x"05",	--1897
		x"5f",	--1898
		x"01",	--1899
		x"5f",	--1900
		x"01",	--1901
		x"d8",	--1902
		x"4f",	--1903
		x"68",	--1904
		x"0e",	--1905
		x"0f",	--1906
		x"0e",	--1907
		x"0f",	--1908
		x"0f",	--1909
		x"69",	--1910
		x"c8",	--1911
		x"01",	--1912
		x"a8",	--1913
		x"02",	--1914
		x"88",	--1915
		x"04",	--1916
		x"88",	--1917
		x"06",	--1918
		x"0c",	--1919
		x"0d",	--1920
		x"3c",	--1921
		x"3d",	--1922
		x"3d",	--1923
		x"ff",	--1924
		x"05",	--1925
		x"3d",	--1926
		x"00",	--1927
		x"17",	--1928
		x"3c",	--1929
		x"15",	--1930
		x"1b",	--1931
		x"02",	--1932
		x"3b",	--1933
		x"0e",	--1934
		x"0f",	--1935
		x"0a",	--1936
		x"3b",	--1937
		x"0c",	--1938
		x"0d",	--1939
		x"3c",	--1940
		x"3d",	--1941
		x"3d",	--1942
		x"ff",	--1943
		x"f5",	--1944
		x"3c",	--1945
		x"88",	--1946
		x"04",	--1947
		x"88",	--1948
		x"06",	--1949
		x"88",	--1950
		x"02",	--1951
		x"f8",	--1952
		x"03",	--1953
		x"00",	--1954
		x"0f",	--1955
		x"b3",	--1956
		x"0c",	--1957
		x"0d",	--1958
		x"1c",	--1959
		x"0d",	--1960
		x"12",	--1961
		x"0f",	--1962
		x"0e",	--1963
		x"0a",	--1964
		x"0b",	--1965
		x"0a",	--1966
		x"0b",	--1967
		x"88",	--1968
		x"04",	--1969
		x"88",	--1970
		x"06",	--1971
		x"98",	--1972
		x"02",	--1973
		x"0f",	--1974
		x"a1",	--1975
		x"6b",	--1976
		x"9f",	--1977
		x"ad",	--1978
		x"00",	--1979
		x"9d",	--1980
		x"02",	--1981
		x"02",	--1982
		x"9d",	--1983
		x"04",	--1984
		x"04",	--1985
		x"9d",	--1986
		x"06",	--1987
		x"06",	--1988
		x"5e",	--1989
		x"01",	--1990
		x"5e",	--1991
		x"01",	--1992
		x"cd",	--1993
		x"01",	--1994
		x"0f",	--1995
		x"8c",	--1996
		x"06",	--1997
		x"07",	--1998
		x"9a",	--1999
		x"39",	--2000
		x"19",	--2001
		x"39",	--2002
		x"20",	--2003
		x"8f",	--2004
		x"3e",	--2005
		x"3c",	--2006
		x"b6",	--2007
		x"c1",	--2008
		x"0e",	--2009
		x"0f",	--2010
		x"0e",	--2011
		x"0f",	--2012
		x"97",	--2013
		x"0f",	--2014
		x"79",	--2015
		x"d8",	--2016
		x"01",	--2017
		x"a8",	--2018
		x"02",	--2019
		x"3e",	--2020
		x"3f",	--2021
		x"1e",	--2022
		x"0f",	--2023
		x"88",	--2024
		x"04",	--2025
		x"88",	--2026
		x"06",	--2027
		x"92",	--2028
		x"0c",	--2029
		x"7b",	--2030
		x"81",	--2031
		x"00",	--2032
		x"81",	--2033
		x"02",	--2034
		x"81",	--2035
		x"04",	--2036
		x"4d",	--2037
		x"7d",	--2038
		x"1f",	--2039
		x"0c",	--2040
		x"4b",	--2041
		x"0c",	--2042
		x"0d",	--2043
		x"12",	--2044
		x"0d",	--2045
		x"0c",	--2046
		x"7b",	--2047
		x"fb",	--2048
		x"81",	--2049
		x"02",	--2050
		x"81",	--2051
		x"04",	--2052
		x"1c",	--2053
		x"0d",	--2054
		x"79",	--2055
		x"1f",	--2056
		x"04",	--2057
		x"0c",	--2058
		x"0d",	--2059
		x"79",	--2060
		x"fc",	--2061
		x"3c",	--2062
		x"3d",	--2063
		x"0c",	--2064
		x"0d",	--2065
		x"1a",	--2066
		x"0b",	--2067
		x"0c",	--2068
		x"04",	--2069
		x"0d",	--2070
		x"02",	--2071
		x"0a",	--2072
		x"0b",	--2073
		x"14",	--2074
		x"02",	--2075
		x"15",	--2076
		x"04",	--2077
		x"04",	--2078
		x"05",	--2079
		x"49",	--2080
		x"0a",	--2081
		x"0b",	--2082
		x"18",	--2083
		x"6c",	--2084
		x"33",	--2085
		x"df",	--2086
		x"01",	--2087
		x"01",	--2088
		x"2f",	--2089
		x"3f",	--2090
		x"90",	--2091
		x"2c",	--2092
		x"31",	--2093
		x"e0",	--2094
		x"81",	--2095
		x"04",	--2096
		x"81",	--2097
		x"06",	--2098
		x"81",	--2099
		x"00",	--2100
		x"81",	--2101
		x"02",	--2102
		x"0e",	--2103
		x"3e",	--2104
		x"18",	--2105
		x"0f",	--2106
		x"2f",	--2107
		x"b0",	--2108
		x"7c",	--2109
		x"0e",	--2110
		x"3e",	--2111
		x"10",	--2112
		x"0f",	--2113
		x"b0",	--2114
		x"7c",	--2115
		x"0d",	--2116
		x"3d",	--2117
		x"0e",	--2118
		x"3e",	--2119
		x"10",	--2120
		x"0f",	--2121
		x"3f",	--2122
		x"18",	--2123
		x"b0",	--2124
		x"c8",	--2125
		x"b0",	--2126
		x"9e",	--2127
		x"31",	--2128
		x"20",	--2129
		x"30",	--2130
		x"31",	--2131
		x"e0",	--2132
		x"81",	--2133
		x"04",	--2134
		x"81",	--2135
		x"06",	--2136
		x"81",	--2137
		x"00",	--2138
		x"81",	--2139
		x"02",	--2140
		x"0e",	--2141
		x"3e",	--2142
		x"18",	--2143
		x"0f",	--2144
		x"2f",	--2145
		x"b0",	--2146
		x"7c",	--2147
		x"0e",	--2148
		x"3e",	--2149
		x"10",	--2150
		x"0f",	--2151
		x"b0",	--2152
		x"7c",	--2153
		x"d1",	--2154
		x"11",	--2155
		x"0d",	--2156
		x"3d",	--2157
		x"0e",	--2158
		x"3e",	--2159
		x"10",	--2160
		x"0f",	--2161
		x"3f",	--2162
		x"18",	--2163
		x"b0",	--2164
		x"c8",	--2165
		x"b0",	--2166
		x"9e",	--2167
		x"31",	--2168
		x"20",	--2169
		x"30",	--2170
		x"0b",	--2171
		x"0a",	--2172
		x"09",	--2173
		x"08",	--2174
		x"07",	--2175
		x"06",	--2176
		x"05",	--2177
		x"04",	--2178
		x"31",	--2179
		x"dc",	--2180
		x"81",	--2181
		x"04",	--2182
		x"81",	--2183
		x"06",	--2184
		x"81",	--2185
		x"00",	--2186
		x"81",	--2187
		x"02",	--2188
		x"0e",	--2189
		x"3e",	--2190
		x"18",	--2191
		x"0f",	--2192
		x"2f",	--2193
		x"b0",	--2194
		x"7c",	--2195
		x"0e",	--2196
		x"3e",	--2197
		x"10",	--2198
		x"0f",	--2199
		x"b0",	--2200
		x"7c",	--2201
		x"5f",	--2202
		x"18",	--2203
		x"6f",	--2204
		x"b6",	--2205
		x"5e",	--2206
		x"10",	--2207
		x"6e",	--2208
		x"d9",	--2209
		x"6f",	--2210
		x"ae",	--2211
		x"6e",	--2212
		x"e2",	--2213
		x"6f",	--2214
		x"ac",	--2215
		x"6e",	--2216
		x"d1",	--2217
		x"14",	--2218
		x"1c",	--2219
		x"15",	--2220
		x"1e",	--2221
		x"18",	--2222
		x"14",	--2223
		x"19",	--2224
		x"16",	--2225
		x"3c",	--2226
		x"20",	--2227
		x"0e",	--2228
		x"0f",	--2229
		x"06",	--2230
		x"07",	--2231
		x"81",	--2232
		x"20",	--2233
		x"81",	--2234
		x"22",	--2235
		x"0a",	--2236
		x"0b",	--2237
		x"81",	--2238
		x"20",	--2239
		x"08",	--2240
		x"08",	--2241
		x"09",	--2242
		x"12",	--2243
		x"05",	--2244
		x"04",	--2245
		x"b1",	--2246
		x"20",	--2247
		x"19",	--2248
		x"14",	--2249
		x"0d",	--2250
		x"0a",	--2251
		x"0b",	--2252
		x"0e",	--2253
		x"0f",	--2254
		x"1c",	--2255
		x"0d",	--2256
		x"0b",	--2257
		x"03",	--2258
		x"0b",	--2259
		x"0c",	--2260
		x"0d",	--2261
		x"0e",	--2262
		x"0f",	--2263
		x"06",	--2264
		x"07",	--2265
		x"09",	--2266
		x"e5",	--2267
		x"16",	--2268
		x"07",	--2269
		x"e2",	--2270
		x"0a",	--2271
		x"f5",	--2272
		x"f2",	--2273
		x"81",	--2274
		x"20",	--2275
		x"81",	--2276
		x"22",	--2277
		x"0c",	--2278
		x"1a",	--2279
		x"1a",	--2280
		x"1a",	--2281
		x"12",	--2282
		x"06",	--2283
		x"26",	--2284
		x"81",	--2285
		x"0a",	--2286
		x"5d",	--2287
		x"d1",	--2288
		x"11",	--2289
		x"19",	--2290
		x"83",	--2291
		x"c1",	--2292
		x"09",	--2293
		x"0c",	--2294
		x"3c",	--2295
		x"3f",	--2296
		x"00",	--2297
		x"18",	--2298
		x"1d",	--2299
		x"0a",	--2300
		x"3d",	--2301
		x"1a",	--2302
		x"20",	--2303
		x"1b",	--2304
		x"22",	--2305
		x"0c",	--2306
		x"0e",	--2307
		x"0f",	--2308
		x"0b",	--2309
		x"2a",	--2310
		x"0a",	--2311
		x"0b",	--2312
		x"3d",	--2313
		x"3f",	--2314
		x"00",	--2315
		x"f5",	--2316
		x"81",	--2317
		x"20",	--2318
		x"81",	--2319
		x"22",	--2320
		x"81",	--2321
		x"0a",	--2322
		x"0c",	--2323
		x"0d",	--2324
		x"3c",	--2325
		x"7f",	--2326
		x"0d",	--2327
		x"3c",	--2328
		x"40",	--2329
		x"44",	--2330
		x"81",	--2331
		x"0c",	--2332
		x"81",	--2333
		x"0e",	--2334
		x"f1",	--2335
		x"03",	--2336
		x"08",	--2337
		x"0f",	--2338
		x"3f",	--2339
		x"b0",	--2340
		x"9e",	--2341
		x"31",	--2342
		x"24",	--2343
		x"34",	--2344
		x"35",	--2345
		x"36",	--2346
		x"37",	--2347
		x"38",	--2348
		x"39",	--2349
		x"3a",	--2350
		x"3b",	--2351
		x"30",	--2352
		x"1e",	--2353
		x"0f",	--2354
		x"d3",	--2355
		x"3a",	--2356
		x"03",	--2357
		x"08",	--2358
		x"1e",	--2359
		x"10",	--2360
		x"1c",	--2361
		x"20",	--2362
		x"1d",	--2363
		x"22",	--2364
		x"12",	--2365
		x"0d",	--2366
		x"0c",	--2367
		x"06",	--2368
		x"07",	--2369
		x"06",	--2370
		x"37",	--2371
		x"00",	--2372
		x"81",	--2373
		x"20",	--2374
		x"81",	--2375
		x"22",	--2376
		x"12",	--2377
		x"0f",	--2378
		x"0e",	--2379
		x"1a",	--2380
		x"0f",	--2381
		x"e7",	--2382
		x"81",	--2383
		x"0a",	--2384
		x"a6",	--2385
		x"6e",	--2386
		x"36",	--2387
		x"5f",	--2388
		x"d1",	--2389
		x"11",	--2390
		x"19",	--2391
		x"20",	--2392
		x"c1",	--2393
		x"19",	--2394
		x"0f",	--2395
		x"3f",	--2396
		x"18",	--2397
		x"c5",	--2398
		x"0d",	--2399
		x"ba",	--2400
		x"0c",	--2401
		x"0d",	--2402
		x"3c",	--2403
		x"80",	--2404
		x"0d",	--2405
		x"0c",	--2406
		x"b3",	--2407
		x"0d",	--2408
		x"b1",	--2409
		x"81",	--2410
		x"20",	--2411
		x"03",	--2412
		x"81",	--2413
		x"22",	--2414
		x"ab",	--2415
		x"3e",	--2416
		x"40",	--2417
		x"0f",	--2418
		x"3e",	--2419
		x"80",	--2420
		x"3f",	--2421
		x"a4",	--2422
		x"4d",	--2423
		x"7b",	--2424
		x"4f",	--2425
		x"de",	--2426
		x"5f",	--2427
		x"d1",	--2428
		x"11",	--2429
		x"19",	--2430
		x"06",	--2431
		x"c1",	--2432
		x"11",	--2433
		x"0f",	--2434
		x"3f",	--2435
		x"10",	--2436
		x"9e",	--2437
		x"4f",	--2438
		x"f8",	--2439
		x"6f",	--2440
		x"f1",	--2441
		x"3f",	--2442
		x"90",	--2443
		x"97",	--2444
		x"0b",	--2445
		x"0a",	--2446
		x"09",	--2447
		x"08",	--2448
		x"07",	--2449
		x"31",	--2450
		x"e8",	--2451
		x"81",	--2452
		x"04",	--2453
		x"81",	--2454
		x"06",	--2455
		x"81",	--2456
		x"00",	--2457
		x"81",	--2458
		x"02",	--2459
		x"0e",	--2460
		x"3e",	--2461
		x"10",	--2462
		x"0f",	--2463
		x"2f",	--2464
		x"b0",	--2465
		x"7c",	--2466
		x"0e",	--2467
		x"3e",	--2468
		x"0f",	--2469
		x"b0",	--2470
		x"7c",	--2471
		x"5f",	--2472
		x"10",	--2473
		x"6f",	--2474
		x"5d",	--2475
		x"5e",	--2476
		x"08",	--2477
		x"6e",	--2478
		x"82",	--2479
		x"d1",	--2480
		x"09",	--2481
		x"11",	--2482
		x"6f",	--2483
		x"58",	--2484
		x"6f",	--2485
		x"56",	--2486
		x"6e",	--2487
		x"6f",	--2488
		x"6e",	--2489
		x"4c",	--2490
		x"1d",	--2491
		x"12",	--2492
		x"1d",	--2493
		x"0a",	--2494
		x"81",	--2495
		x"12",	--2496
		x"1e",	--2497
		x"14",	--2498
		x"1f",	--2499
		x"16",	--2500
		x"18",	--2501
		x"0c",	--2502
		x"19",	--2503
		x"0e",	--2504
		x"0f",	--2505
		x"1e",	--2506
		x"0e",	--2507
		x"0f",	--2508
		x"3d",	--2509
		x"81",	--2510
		x"12",	--2511
		x"37",	--2512
		x"1f",	--2513
		x"0c",	--2514
		x"3d",	--2515
		x"00",	--2516
		x"0a",	--2517
		x"0b",	--2518
		x"0b",	--2519
		x"0a",	--2520
		x"0b",	--2521
		x"0e",	--2522
		x"0f",	--2523
		x"12",	--2524
		x"0d",	--2525
		x"0c",	--2526
		x"0e",	--2527
		x"0f",	--2528
		x"37",	--2529
		x"0b",	--2530
		x"0f",	--2531
		x"f7",	--2532
		x"f2",	--2533
		x"0e",	--2534
		x"f4",	--2535
		x"ef",	--2536
		x"09",	--2537
		x"e5",	--2538
		x"0e",	--2539
		x"e3",	--2540
		x"dd",	--2541
		x"0c",	--2542
		x"0d",	--2543
		x"3c",	--2544
		x"7f",	--2545
		x"0d",	--2546
		x"3c",	--2547
		x"40",	--2548
		x"1c",	--2549
		x"81",	--2550
		x"14",	--2551
		x"81",	--2552
		x"16",	--2553
		x"0f",	--2554
		x"3f",	--2555
		x"10",	--2556
		x"b0",	--2557
		x"9e",	--2558
		x"31",	--2559
		x"18",	--2560
		x"37",	--2561
		x"38",	--2562
		x"39",	--2563
		x"3a",	--2564
		x"3b",	--2565
		x"30",	--2566
		x"e1",	--2567
		x"10",	--2568
		x"0f",	--2569
		x"3f",	--2570
		x"10",	--2571
		x"f0",	--2572
		x"4f",	--2573
		x"fa",	--2574
		x"3f",	--2575
		x"90",	--2576
		x"eb",	--2577
		x"0d",	--2578
		x"e2",	--2579
		x"0c",	--2580
		x"0d",	--2581
		x"3c",	--2582
		x"80",	--2583
		x"0d",	--2584
		x"0c",	--2585
		x"db",	--2586
		x"0d",	--2587
		x"d9",	--2588
		x"0e",	--2589
		x"02",	--2590
		x"0f",	--2591
		x"d5",	--2592
		x"3a",	--2593
		x"40",	--2594
		x"0b",	--2595
		x"3a",	--2596
		x"80",	--2597
		x"3b",	--2598
		x"ce",	--2599
		x"81",	--2600
		x"14",	--2601
		x"81",	--2602
		x"16",	--2603
		x"81",	--2604
		x"12",	--2605
		x"0f",	--2606
		x"3f",	--2607
		x"10",	--2608
		x"cb",	--2609
		x"0f",	--2610
		x"3f",	--2611
		x"c8",	--2612
		x"31",	--2613
		x"e8",	--2614
		x"81",	--2615
		x"04",	--2616
		x"81",	--2617
		x"06",	--2618
		x"81",	--2619
		x"00",	--2620
		x"81",	--2621
		x"02",	--2622
		x"0e",	--2623
		x"3e",	--2624
		x"10",	--2625
		x"0f",	--2626
		x"2f",	--2627
		x"b0",	--2628
		x"7c",	--2629
		x"0e",	--2630
		x"3e",	--2631
		x"0f",	--2632
		x"b0",	--2633
		x"7c",	--2634
		x"e1",	--2635
		x"10",	--2636
		x"0d",	--2637
		x"e1",	--2638
		x"08",	--2639
		x"0a",	--2640
		x"0e",	--2641
		x"3e",	--2642
		x"0f",	--2643
		x"3f",	--2644
		x"10",	--2645
		x"b0",	--2646
		x"a0",	--2647
		x"31",	--2648
		x"18",	--2649
		x"30",	--2650
		x"3f",	--2651
		x"fb",	--2652
		x"31",	--2653
		x"f4",	--2654
		x"81",	--2655
		x"00",	--2656
		x"81",	--2657
		x"02",	--2658
		x"0e",	--2659
		x"2e",	--2660
		x"0f",	--2661
		x"b0",	--2662
		x"7c",	--2663
		x"5f",	--2664
		x"04",	--2665
		x"6f",	--2666
		x"28",	--2667
		x"27",	--2668
		x"6f",	--2669
		x"07",	--2670
		x"1d",	--2671
		x"06",	--2672
		x"0d",	--2673
		x"21",	--2674
		x"3d",	--2675
		x"1f",	--2676
		x"09",	--2677
		x"c1",	--2678
		x"05",	--2679
		x"26",	--2680
		x"3e",	--2681
		x"3f",	--2682
		x"ff",	--2683
		x"31",	--2684
		x"0c",	--2685
		x"30",	--2686
		x"1e",	--2687
		x"08",	--2688
		x"1f",	--2689
		x"0a",	--2690
		x"3c",	--2691
		x"1e",	--2692
		x"4c",	--2693
		x"4d",	--2694
		x"7d",	--2695
		x"1f",	--2696
		x"0f",	--2697
		x"c1",	--2698
		x"05",	--2699
		x"ef",	--2700
		x"3e",	--2701
		x"3f",	--2702
		x"1e",	--2703
		x"0f",	--2704
		x"31",	--2705
		x"0c",	--2706
		x"30",	--2707
		x"0e",	--2708
		x"0f",	--2709
		x"31",	--2710
		x"0c",	--2711
		x"30",	--2712
		x"12",	--2713
		x"0f",	--2714
		x"0e",	--2715
		x"7d",	--2716
		x"fb",	--2717
		x"eb",	--2718
		x"0e",	--2719
		x"3f",	--2720
		x"00",	--2721
		x"31",	--2722
		x"0c",	--2723
		x"30",	--2724
		x"0b",	--2725
		x"0a",	--2726
		x"09",	--2727
		x"08",	--2728
		x"31",	--2729
		x"0a",	--2730
		x"0b",	--2731
		x"c1",	--2732
		x"01",	--2733
		x"0e",	--2734
		x"0d",	--2735
		x"0b",	--2736
		x"0b",	--2737
		x"e1",	--2738
		x"00",	--2739
		x"0f",	--2740
		x"b0",	--2741
		x"9e",	--2742
		x"31",	--2743
		x"38",	--2744
		x"39",	--2745
		x"3a",	--2746
		x"3b",	--2747
		x"30",	--2748
		x"f1",	--2749
		x"03",	--2750
		x"00",	--2751
		x"b1",	--2752
		x"1e",	--2753
		x"02",	--2754
		x"81",	--2755
		x"04",	--2756
		x"81",	--2757
		x"06",	--2758
		x"0e",	--2759
		x"0f",	--2760
		x"b0",	--2761
		x"2c",	--2762
		x"3f",	--2763
		x"0f",	--2764
		x"18",	--2765
		x"e5",	--2766
		x"81",	--2767
		x"04",	--2768
		x"81",	--2769
		x"06",	--2770
		x"4e",	--2771
		x"7e",	--2772
		x"1f",	--2773
		x"06",	--2774
		x"3e",	--2775
		x"1e",	--2776
		x"0e",	--2777
		x"81",	--2778
		x"02",	--2779
		x"d7",	--2780
		x"91",	--2781
		x"04",	--2782
		x"04",	--2783
		x"91",	--2784
		x"06",	--2785
		x"06",	--2786
		x"7e",	--2787
		x"f8",	--2788
		x"f1",	--2789
		x"0e",	--2790
		x"3e",	--2791
		x"1e",	--2792
		x"1c",	--2793
		x"0d",	--2794
		x"48",	--2795
		x"78",	--2796
		x"1f",	--2797
		x"04",	--2798
		x"0c",	--2799
		x"0d",	--2800
		x"78",	--2801
		x"fc",	--2802
		x"3c",	--2803
		x"3d",	--2804
		x"0c",	--2805
		x"0d",	--2806
		x"18",	--2807
		x"09",	--2808
		x"0c",	--2809
		x"04",	--2810
		x"0d",	--2811
		x"02",	--2812
		x"08",	--2813
		x"09",	--2814
		x"7e",	--2815
		x"1f",	--2816
		x"0e",	--2817
		x"0d",	--2818
		x"0e",	--2819
		x"0d",	--2820
		x"0e",	--2821
		x"81",	--2822
		x"04",	--2823
		x"81",	--2824
		x"06",	--2825
		x"3e",	--2826
		x"1e",	--2827
		x"0e",	--2828
		x"81",	--2829
		x"02",	--2830
		x"a4",	--2831
		x"12",	--2832
		x"0b",	--2833
		x"0a",	--2834
		x"7e",	--2835
		x"fb",	--2836
		x"ec",	--2837
		x"0b",	--2838
		x"0a",	--2839
		x"09",	--2840
		x"1f",	--2841
		x"17",	--2842
		x"3e",	--2843
		x"00",	--2844
		x"2c",	--2845
		x"3a",	--2846
		x"18",	--2847
		x"0b",	--2848
		x"39",	--2849
		x"0c",	--2850
		x"0d",	--2851
		x"4f",	--2852
		x"4f",	--2853
		x"17",	--2854
		x"3c",	--2855
		x"98",	--2856
		x"6e",	--2857
		x"0f",	--2858
		x"0a",	--2859
		x"0b",	--2860
		x"0f",	--2861
		x"39",	--2862
		x"3a",	--2863
		x"3b",	--2864
		x"30",	--2865
		x"3f",	--2866
		x"00",	--2867
		x"0f",	--2868
		x"3a",	--2869
		x"0b",	--2870
		x"39",	--2871
		x"18",	--2872
		x"0c",	--2873
		x"0d",	--2874
		x"4f",	--2875
		x"4f",	--2876
		x"e9",	--2877
		x"12",	--2878
		x"0d",	--2879
		x"0c",	--2880
		x"7f",	--2881
		x"fb",	--2882
		x"e3",	--2883
		x"3a",	--2884
		x"10",	--2885
		x"0b",	--2886
		x"39",	--2887
		x"10",	--2888
		x"ef",	--2889
		x"3a",	--2890
		x"20",	--2891
		x"0b",	--2892
		x"09",	--2893
		x"ea",	--2894
		x"0b",	--2895
		x"0a",	--2896
		x"09",	--2897
		x"08",	--2898
		x"07",	--2899
		x"0d",	--2900
		x"1e",	--2901
		x"04",	--2902
		x"1f",	--2903
		x"06",	--2904
		x"5a",	--2905
		x"01",	--2906
		x"6c",	--2907
		x"6c",	--2908
		x"70",	--2909
		x"6c",	--2910
		x"6a",	--2911
		x"6c",	--2912
		x"36",	--2913
		x"0e",	--2914
		x"32",	--2915
		x"1b",	--2916
		x"02",	--2917
		x"3b",	--2918
		x"82",	--2919
		x"6d",	--2920
		x"3b",	--2921
		x"80",	--2922
		x"5e",	--2923
		x"0c",	--2924
		x"0d",	--2925
		x"3c",	--2926
		x"7f",	--2927
		x"0d",	--2928
		x"3c",	--2929
		x"40",	--2930
		x"40",	--2931
		x"3e",	--2932
		x"3f",	--2933
		x"0f",	--2934
		x"0f",	--2935
		x"4a",	--2936
		x"0d",	--2937
		x"3d",	--2938
		x"7f",	--2939
		x"12",	--2940
		x"0f",	--2941
		x"0e",	--2942
		x"12",	--2943
		x"0f",	--2944
		x"0e",	--2945
		x"12",	--2946
		x"0f",	--2947
		x"0e",	--2948
		x"12",	--2949
		x"0f",	--2950
		x"0e",	--2951
		x"12",	--2952
		x"0f",	--2953
		x"0e",	--2954
		x"12",	--2955
		x"0f",	--2956
		x"0e",	--2957
		x"12",	--2958
		x"0f",	--2959
		x"0e",	--2960
		x"3e",	--2961
		x"3f",	--2962
		x"7f",	--2963
		x"4d",	--2964
		x"05",	--2965
		x"0f",	--2966
		x"cc",	--2967
		x"4d",	--2968
		x"0e",	--2969
		x"0f",	--2970
		x"4d",	--2971
		x"0d",	--2972
		x"0d",	--2973
		x"0d",	--2974
		x"0d",	--2975
		x"0d",	--2976
		x"0d",	--2977
		x"0d",	--2978
		x"0c",	--2979
		x"3c",	--2980
		x"7f",	--2981
		x"0c",	--2982
		x"4f",	--2983
		x"0f",	--2984
		x"0f",	--2985
		x"0f",	--2986
		x"0d",	--2987
		x"0d",	--2988
		x"0f",	--2989
		x"37",	--2990
		x"38",	--2991
		x"39",	--2992
		x"3a",	--2993
		x"3b",	--2994
		x"30",	--2995
		x"0d",	--2996
		x"be",	--2997
		x"0c",	--2998
		x"0d",	--2999
		x"3c",	--3000
		x"80",	--3001
		x"0d",	--3002
		x"0c",	--3003
		x"02",	--3004
		x"0d",	--3005
		x"b8",	--3006
		x"3e",	--3007
		x"40",	--3008
		x"0f",	--3009
		x"b4",	--3010
		x"12",	--3011
		x"0f",	--3012
		x"0e",	--3013
		x"0d",	--3014
		x"3d",	--3015
		x"80",	--3016
		x"b2",	--3017
		x"7d",	--3018
		x"0e",	--3019
		x"0f",	--3020
		x"cd",	--3021
		x"0e",	--3022
		x"3f",	--3023
		x"10",	--3024
		x"3e",	--3025
		x"3f",	--3026
		x"7f",	--3027
		x"7d",	--3028
		x"c5",	--3029
		x"37",	--3030
		x"82",	--3031
		x"07",	--3032
		x"37",	--3033
		x"1a",	--3034
		x"4f",	--3035
		x"0c",	--3036
		x"0d",	--3037
		x"4b",	--3038
		x"7b",	--3039
		x"1f",	--3040
		x"05",	--3041
		x"12",	--3042
		x"0d",	--3043
		x"0c",	--3044
		x"7b",	--3045
		x"fb",	--3046
		x"18",	--3047
		x"09",	--3048
		x"77",	--3049
		x"1f",	--3050
		x"04",	--3051
		x"08",	--3052
		x"09",	--3053
		x"77",	--3054
		x"fc",	--3055
		x"38",	--3056
		x"39",	--3057
		x"08",	--3058
		x"09",	--3059
		x"1e",	--3060
		x"0f",	--3061
		x"08",	--3062
		x"04",	--3063
		x"09",	--3064
		x"02",	--3065
		x"0e",	--3066
		x"0f",	--3067
		x"08",	--3068
		x"09",	--3069
		x"08",	--3070
		x"09",	--3071
		x"0e",	--3072
		x"0f",	--3073
		x"3e",	--3074
		x"7f",	--3075
		x"0f",	--3076
		x"3e",	--3077
		x"40",	--3078
		x"26",	--3079
		x"38",	--3080
		x"3f",	--3081
		x"09",	--3082
		x"0e",	--3083
		x"0f",	--3084
		x"12",	--3085
		x"0f",	--3086
		x"0e",	--3087
		x"12",	--3088
		x"0f",	--3089
		x"0e",	--3090
		x"12",	--3091
		x"0f",	--3092
		x"0e",	--3093
		x"12",	--3094
		x"0f",	--3095
		x"0e",	--3096
		x"12",	--3097
		x"0f",	--3098
		x"0e",	--3099
		x"12",	--3100
		x"0f",	--3101
		x"0e",	--3102
		x"12",	--3103
		x"0f",	--3104
		x"0e",	--3105
		x"3e",	--3106
		x"3f",	--3107
		x"7f",	--3108
		x"5d",	--3109
		x"39",	--3110
		x"00",	--3111
		x"72",	--3112
		x"4d",	--3113
		x"70",	--3114
		x"08",	--3115
		x"09",	--3116
		x"da",	--3117
		x"0f",	--3118
		x"d8",	--3119
		x"0e",	--3120
		x"0f",	--3121
		x"3e",	--3122
		x"80",	--3123
		x"0f",	--3124
		x"0e",	--3125
		x"04",	--3126
		x"38",	--3127
		x"40",	--3128
		x"09",	--3129
		x"d0",	--3130
		x"0f",	--3131
		x"ce",	--3132
		x"f9",	--3133
		x"0b",	--3134
		x"0a",	--3135
		x"2a",	--3136
		x"5b",	--3137
		x"02",	--3138
		x"3b",	--3139
		x"7f",	--3140
		x"1d",	--3141
		x"02",	--3142
		x"12",	--3143
		x"0d",	--3144
		x"12",	--3145
		x"0d",	--3146
		x"12",	--3147
		x"0d",	--3148
		x"12",	--3149
		x"0d",	--3150
		x"12",	--3151
		x"0d",	--3152
		x"12",	--3153
		x"0d",	--3154
		x"12",	--3155
		x"0d",	--3156
		x"4d",	--3157
		x"5f",	--3158
		x"03",	--3159
		x"3f",	--3160
		x"80",	--3161
		x"0f",	--3162
		x"0f",	--3163
		x"ce",	--3164
		x"01",	--3165
		x"0d",	--3166
		x"2d",	--3167
		x"0a",	--3168
		x"51",	--3169
		x"be",	--3170
		x"82",	--3171
		x"02",	--3172
		x"0c",	--3173
		x"0d",	--3174
		x"0c",	--3175
		x"0d",	--3176
		x"0c",	--3177
		x"0d",	--3178
		x"0c",	--3179
		x"0d",	--3180
		x"0c",	--3181
		x"0d",	--3182
		x"0c",	--3183
		x"0d",	--3184
		x"0c",	--3185
		x"0d",	--3186
		x"0c",	--3187
		x"0d",	--3188
		x"fe",	--3189
		x"03",	--3190
		x"00",	--3191
		x"3d",	--3192
		x"00",	--3193
		x"0b",	--3194
		x"3f",	--3195
		x"81",	--3196
		x"0c",	--3197
		x"0d",	--3198
		x"0a",	--3199
		x"3f",	--3200
		x"3d",	--3201
		x"00",	--3202
		x"f9",	--3203
		x"8e",	--3204
		x"02",	--3205
		x"8e",	--3206
		x"04",	--3207
		x"8e",	--3208
		x"06",	--3209
		x"3a",	--3210
		x"3b",	--3211
		x"30",	--3212
		x"3d",	--3213
		x"ff",	--3214
		x"2a",	--3215
		x"3d",	--3216
		x"81",	--3217
		x"8e",	--3218
		x"02",	--3219
		x"fe",	--3220
		x"03",	--3221
		x"00",	--3222
		x"0c",	--3223
		x"0d",	--3224
		x"0c",	--3225
		x"0d",	--3226
		x"0c",	--3227
		x"0d",	--3228
		x"0c",	--3229
		x"0d",	--3230
		x"0c",	--3231
		x"0d",	--3232
		x"0c",	--3233
		x"0d",	--3234
		x"0c",	--3235
		x"0d",	--3236
		x"0c",	--3237
		x"0d",	--3238
		x"0a",	--3239
		x"0b",	--3240
		x"0a",	--3241
		x"3b",	--3242
		x"00",	--3243
		x"8e",	--3244
		x"04",	--3245
		x"8e",	--3246
		x"06",	--3247
		x"3a",	--3248
		x"3b",	--3249
		x"30",	--3250
		x"0b",	--3251
		x"ad",	--3252
		x"ee",	--3253
		x"00",	--3254
		x"3a",	--3255
		x"3b",	--3256
		x"30",	--3257
		x"0a",	--3258
		x"0c",	--3259
		x"0c",	--3260
		x"0d",	--3261
		x"0c",	--3262
		x"3d",	--3263
		x"10",	--3264
		x"0c",	--3265
		x"02",	--3266
		x"0d",	--3267
		x"08",	--3268
		x"de",	--3269
		x"00",	--3270
		x"e4",	--3271
		x"0b",	--3272
		x"f2",	--3273
		x"ee",	--3274
		x"00",	--3275
		x"e3",	--3276
		x"ce",	--3277
		x"00",	--3278
		x"dc",	--3279
		x"0b",	--3280
		x"6d",	--3281
		x"6d",	--3282
		x"12",	--3283
		x"6c",	--3284
		x"6c",	--3285
		x"0f",	--3286
		x"6d",	--3287
		x"41",	--3288
		x"6c",	--3289
		x"11",	--3290
		x"6d",	--3291
		x"0d",	--3292
		x"6c",	--3293
		x"14",	--3294
		x"5d",	--3295
		x"01",	--3296
		x"5d",	--3297
		x"01",	--3298
		x"14",	--3299
		x"4d",	--3300
		x"09",	--3301
		x"1e",	--3302
		x"0f",	--3303
		x"3b",	--3304
		x"30",	--3305
		x"6c",	--3306
		x"28",	--3307
		x"ce",	--3308
		x"01",	--3309
		x"f7",	--3310
		x"3e",	--3311
		x"0f",	--3312
		x"3b",	--3313
		x"30",	--3314
		x"cf",	--3315
		x"01",	--3316
		x"f0",	--3317
		x"3e",	--3318
		x"f8",	--3319
		x"1b",	--3320
		x"02",	--3321
		x"1c",	--3322
		x"02",	--3323
		x"0c",	--3324
		x"e6",	--3325
		x"0b",	--3326
		x"16",	--3327
		x"1b",	--3328
		x"04",	--3329
		x"1f",	--3330
		x"06",	--3331
		x"1c",	--3332
		x"04",	--3333
		x"1e",	--3334
		x"06",	--3335
		x"0e",	--3336
		x"da",	--3337
		x"0f",	--3338
		x"02",	--3339
		x"0c",	--3340
		x"d6",	--3341
		x"0f",	--3342
		x"06",	--3343
		x"0e",	--3344
		x"02",	--3345
		x"0b",	--3346
		x"02",	--3347
		x"0e",	--3348
		x"d1",	--3349
		x"4d",	--3350
		x"ce",	--3351
		x"3e",	--3352
		x"d6",	--3353
		x"6c",	--3354
		x"d7",	--3355
		x"5e",	--3356
		x"01",	--3357
		x"5f",	--3358
		x"01",	--3359
		x"0e",	--3360
		x"c5",	--3361
		x"0d",	--3362
		x"0f",	--3363
		x"04",	--3364
		x"3d",	--3365
		x"03",	--3366
		x"3f",	--3367
		x"1f",	--3368
		x"0e",	--3369
		x"03",	--3370
		x"5d",	--3371
		x"3e",	--3372
		x"1e",	--3373
		x"0d",	--3374
		x"b0",	--3375
		x"0a",	--3376
		x"3d",	--3377
		x"6d",	--3378
		x"02",	--3379
		x"3e",	--3380
		x"1e",	--3381
		x"5d",	--3382
		x"02",	--3383
		x"3f",	--3384
		x"1f",	--3385
		x"30",	--3386
		x"b0",	--3387
		x"44",	--3388
		x"0f",	--3389
		x"30",	--3390
		x"0b",	--3391
		x"0a",	--3392
		x"09",	--3393
		x"79",	--3394
		x"20",	--3395
		x"0a",	--3396
		x"0b",	--3397
		x"0c",	--3398
		x"0d",	--3399
		x"0e",	--3400
		x"0f",	--3401
		x"0c",	--3402
		x"0d",	--3403
		x"0d",	--3404
		x"06",	--3405
		x"02",	--3406
		x"0c",	--3407
		x"03",	--3408
		x"0c",	--3409
		x"0d",	--3410
		x"1e",	--3411
		x"19",	--3412
		x"f2",	--3413
		x"39",	--3414
		x"3a",	--3415
		x"3b",	--3416
		x"30",	--3417
		x"b0",	--3418
		x"7e",	--3419
		x"0e",	--3420
		x"0f",	--3421
		x"30",	--3422
		x"0b",	--3423
		x"0b",	--3424
		x"0f",	--3425
		x"06",	--3426
		x"3b",	--3427
		x"03",	--3428
		x"3e",	--3429
		x"3f",	--3430
		x"1e",	--3431
		x"0f",	--3432
		x"0d",	--3433
		x"05",	--3434
		x"5b",	--3435
		x"3c",	--3436
		x"3d",	--3437
		x"1c",	--3438
		x"0d",	--3439
		x"b0",	--3440
		x"7e",	--3441
		x"6b",	--3442
		x"04",	--3443
		x"3c",	--3444
		x"3d",	--3445
		x"1c",	--3446
		x"0d",	--3447
		x"5b",	--3448
		x"04",	--3449
		x"3e",	--3450
		x"3f",	--3451
		x"1e",	--3452
		x"0f",	--3453
		x"3b",	--3454
		x"30",	--3455
		x"b0",	--3456
		x"be",	--3457
		x"0e",	--3458
		x"0f",	--3459
		x"30",	--3460
		x"7c",	--3461
		x"10",	--3462
		x"0d",	--3463
		x"0e",	--3464
		x"0f",	--3465
		x"0e",	--3466
		x"0e",	--3467
		x"02",	--3468
		x"0e",	--3469
		x"1f",	--3470
		x"1c",	--3471
		x"f8",	--3472
		x"30",	--3473
		x"b0",	--3474
		x"0a",	--3475
		x"0f",	--3476
		x"30",	--3477
		x"00",	--3478
		x"32",	--3479
		x"f0",	--3480
		x"fd",	--3481
		x"57",	--3482
		x"69",	--3483
		x"69",	--3484
		x"67",	--3485
		x"66",	--3486
		x"72",	--3487
		x"61",	--3488
		x"6e",	--3489
		x"77",	--3490
		x"2e",	--3491
		x"69",	--3492
		x"20",	--3493
		x"69",	--3494
		x"65",	--3495
		x"0a",	--3496
		x"57",	--3497
		x"20",	--3498
		x"68",	--3499
		x"75",	--3500
		x"64",	--3501
		x"6e",	--3502
		x"74",	--3503
		x"73",	--3504
		x"65",	--3505
		x"74",	--3506
		x"61",	--3507
		x"0d",	--3508
		x"00",	--3509
		x"74",	--3510
		x"70",	--3511
		x"0a",	--3512
		x"65",	--3513
		x"72",	--3514
		x"72",	--3515
		x"20",	--3516
		x"69",	--3517
		x"73",	--3518
		x"6e",	--3519
		x"20",	--3520
		x"72",	--3521
		x"75",	--3522
		x"65",	--3523
		x"74",	--3524
		x"0a",	--3525
		x"63",	--3526
		x"72",	--3527
		x"65",	--3528
		x"74",	--3529
		x"75",	--3530
		x"61",	--3531
		x"65",	--3532
		x"0d",	--3533
		x"00",	--3534
		x"25",	--3535
		x"20",	--3536
		x"45",	--3537
		x"54",	--3538
		x"52",	--3539
		x"47",	--3540
		x"54",	--3541
		x"3c",	--3542
		x"49",	--3543
		x"45",	--3544
		x"55",	--3545
		x"3e",	--3546
		x"0a",	--3547
		x"25",	--3548
		x"20",	--3549
		x"64",	--3550
		x"0a",	--3551
		x"25",	--3552
		x"20",	--3553
		x"77",	--3554
		x"25",	--3555
		x"20",	--3556
		x"77",	--3557
		x"0a",	--3558
		x"9c",	--3559
		x"c4",	--3560
		x"ca",	--3561
		x"d2",	--3562
		x"da",	--3563
		x"e2",	--3564
		x"b4",	--3565
		x"bc",	--3566
		x"0d",	--3567
		x"3d",	--3568
		x"3d",	--3569
		x"3d",	--3570
		x"20",	--3571
		x"61",	--3572
		x"63",	--3573
		x"6c",	--3574
		x"4d",	--3575
		x"55",	--3576
		x"3d",	--3577
		x"3d",	--3578
		x"3d",	--3579
		x"0d",	--3580
		x"00",	--3581
		x"6e",	--3582
		x"65",	--3583
		x"61",	--3584
		x"74",	--3585
		x"76",	--3586
		x"20",	--3587
		x"6f",	--3588
		x"65",	--3589
		x"77",	--3590
		x"69",	--3591
		x"65",	--3592
		x"72",	--3593
		x"61",	--3594
		x"00",	--3595
		x"77",	--3596
		x"00",	--3597
		x"6e",	--3598
		x"6f",	--3599
		x"65",	--3600
		x"00",	--3601
		x"6f",	--3602
		x"74",	--3603
		x"6f",	--3604
		x"64",	--3605
		x"72",	--3606
		x"0d",	--3607
		x"00",	--3608
		x"20",	--3609
		x"00",	--3610
		x"63",	--3611
		x"77",	--3612
		x"69",	--3613
		x"65",	--3614
		x"0d",	--3615
		x"65",	--3616
		x"72",	--3617
		x"72",	--3618
		x"20",	--3619
		x"69",	--3620
		x"73",	--3621
		x"6e",	--3622
		x"20",	--3623
		x"72",	--3624
		x"75",	--3625
		x"65",	--3626
		x"74",	--3627
		x"0a",	--3628
		x"63",	--3629
		x"72",	--3630
		x"65",	--3631
		x"74",	--3632
		x"75",	--3633
		x"61",	--3634
		x"65",	--3635
		x"0d",	--3636
		x"00",	--3637
		x"25",	--3638
		x"20",	--3639
		x"45",	--3640
		x"49",	--3641
		x"54",	--3642
		x"52",	--3643
		x"56",	--3644
		x"4c",	--3645
		x"45",	--3646
		x"0a",	--3647
		x"72",	--3648
		x"25",	--3649
		x"20",	--3650
		x"3d",	--3651
		x"64",	--3652
		x"0a",	--3653
		x"09",	--3654
		x"73",	--3655
		x"52",	--3656
		x"47",	--3657
		x"53",	--3658
		x"45",	--3659
		x"0d",	--3660
		x"00",	--3661
		x"65",	--3662
		x"64",	--3663
		x"0d",	--3664
		x"25",	--3665
		x"20",	--3666
		x"73",	--3667
		x"6e",	--3668
		x"74",	--3669
		x"61",	--3670
		x"6e",	--3671
		x"6d",	--3672
		x"65",	--3673
		x"0d",	--3674
		x"00",	--3675
		x"63",	--3676
		x"25",	--3677
		x"0d",	--3678
		x"00",	--3679
		x"63",	--3680
		x"20",	--3681
		x"6f",	--3682
		x"73",	--3683
		x"63",	--3684
		x"20",	--3685
		x"6f",	--3686
		x"6d",	--3687
		x"6e",	--3688
		x"0d",	--3689
		x"00",	--3690
		x"c4",	--3691
		x"f2",	--3692
		x"f2",	--3693
		x"f2",	--3694
		x"f2",	--3695
		x"f2",	--3696
		x"f2",	--3697
		x"f2",	--3698
		x"f2",	--3699
		x"f2",	--3700
		x"f2",	--3701
		x"f2",	--3702
		x"f2",	--3703
		x"f2",	--3704
		x"f2",	--3705
		x"f2",	--3706
		x"f2",	--3707
		x"f2",	--3708
		x"f2",	--3709
		x"f2",	--3710
		x"f2",	--3711
		x"f2",	--3712
		x"f2",	--3713
		x"f2",	--3714
		x"f2",	--3715
		x"f2",	--3716
		x"f2",	--3717
		x"f2",	--3718
		x"f2",	--3719
		x"b6",	--3720
		x"f2",	--3721
		x"f2",	--3722
		x"f2",	--3723
		x"f2",	--3724
		x"f2",	--3725
		x"f2",	--3726
		x"f2",	--3727
		x"f2",	--3728
		x"f2",	--3729
		x"f2",	--3730
		x"f2",	--3731
		x"f2",	--3732
		x"f2",	--3733
		x"f2",	--3734
		x"f2",	--3735
		x"f2",	--3736
		x"f2",	--3737
		x"f2",	--3738
		x"f2",	--3739
		x"f2",	--3740
		x"f2",	--3741
		x"f2",	--3742
		x"f2",	--3743
		x"f2",	--3744
		x"f2",	--3745
		x"f2",	--3746
		x"f2",	--3747
		x"f2",	--3748
		x"f2",	--3749
		x"f2",	--3750
		x"f2",	--3751
		x"a8",	--3752
		x"9a",	--3753
		x"8c",	--3754
		x"f2",	--3755
		x"f2",	--3756
		x"f2",	--3757
		x"f2",	--3758
		x"f2",	--3759
		x"f2",	--3760
		x"f2",	--3761
		x"74",	--3762
		x"f2",	--3763
		x"62",	--3764
		x"f2",	--3765
		x"f2",	--3766
		x"f2",	--3767
		x"f2",	--3768
		x"46",	--3769
		x"f2",	--3770
		x"f2",	--3771
		x"f2",	--3772
		x"38",	--3773
		x"26",	--3774
		x"30",	--3775
		x"32",	--3776
		x"34",	--3777
		x"36",	--3778
		x"38",	--3779
		x"61",	--3780
		x"63",	--3781
		x"65",	--3782
		x"00",	--3783
		x"00",	--3784
		x"00",	--3785
		x"00",	--3786
		x"00",	--3787
		x"00",	--3788
		x"02",	--3789
		x"03",	--3790
		x"03",	--3791
		x"04",	--3792
		x"04",	--3793
		x"04",	--3794
		x"04",	--3795
		x"05",	--3796
		x"05",	--3797
		x"05",	--3798
		x"05",	--3799
		x"05",	--3800
		x"05",	--3801
		x"05",	--3802
		x"05",	--3803
		x"06",	--3804
		x"06",	--3805
		x"06",	--3806
		x"06",	--3807
		x"06",	--3808
		x"06",	--3809
		x"06",	--3810
		x"06",	--3811
		x"06",	--3812
		x"06",	--3813
		x"06",	--3814
		x"06",	--3815
		x"06",	--3816
		x"06",	--3817
		x"06",	--3818
		x"06",	--3819
		x"07",	--3820
		x"07",	--3821
		x"07",	--3822
		x"07",	--3823
		x"07",	--3824
		x"07",	--3825
		x"07",	--3826
		x"07",	--3827
		x"07",	--3828
		x"07",	--3829
		x"07",	--3830
		x"07",	--3831
		x"07",	--3832
		x"07",	--3833
		x"07",	--3834
		x"07",	--3835
		x"07",	--3836
		x"07",	--3837
		x"07",	--3838
		x"07",	--3839
		x"07",	--3840
		x"07",	--3841
		x"07",	--3842
		x"07",	--3843
		x"07",	--3844
		x"07",	--3845
		x"07",	--3846
		x"07",	--3847
		x"07",	--3848
		x"07",	--3849
		x"07",	--3850
		x"07",	--3851
		x"08",	--3852
		x"08",	--3853
		x"08",	--3854
		x"08",	--3855
		x"08",	--3856
		x"08",	--3857
		x"08",	--3858
		x"08",	--3859
		x"08",	--3860
		x"08",	--3861
		x"08",	--3862
		x"08",	--3863
		x"08",	--3864
		x"08",	--3865
		x"08",	--3866
		x"08",	--3867
		x"08",	--3868
		x"08",	--3869
		x"08",	--3870
		x"08",	--3871
		x"08",	--3872
		x"08",	--3873
		x"08",	--3874
		x"08",	--3875
		x"08",	--3876
		x"08",	--3877
		x"08",	--3878
		x"08",	--3879
		x"08",	--3880
		x"08",	--3881
		x"08",	--3882
		x"08",	--3883
		x"08",	--3884
		x"08",	--3885
		x"08",	--3886
		x"08",	--3887
		x"08",	--3888
		x"08",	--3889
		x"08",	--3890
		x"08",	--3891
		x"08",	--3892
		x"08",	--3893
		x"08",	--3894
		x"08",	--3895
		x"08",	--3896
		x"08",	--3897
		x"08",	--3898
		x"08",	--3899
		x"08",	--3900
		x"08",	--3901
		x"08",	--3902
		x"08",	--3903
		x"08",	--3904
		x"08",	--3905
		x"08",	--3906
		x"08",	--3907
		x"08",	--3908
		x"08",	--3909
		x"08",	--3910
		x"08",	--3911
		x"08",	--3912
		x"08",	--3913
		x"08",	--3914
		x"08",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"68",	--3918
		x"6c",	--3919
		x"00",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"da",	--4080
		x"da",	--4081
		x"da",	--4082
		x"da",	--4083
		x"da",	--4084
		x"da",	--4085
		x"da",	--4086
		x"ce",	--4087
		x"54",	--4088
		x"da",	--4089
		x"da",	--4090
		x"da",	--4091
		x"da",	--4092
		x"da",	--4093
		x"da",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"04",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"04",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fe",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"02",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"04",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"ed",	--44
		x"12",	--45
		x"e7",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"fb",	--50
		x"12",	--51
		x"eb",	--52
		x"53",	--53
		x"40",	--54
		x"fb",	--55
		x"40",	--56
		x"e4",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"e7",	--61
		x"40",	--62
		x"fc",	--63
		x"40",	--64
		x"e5",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"e7",	--69
		x"40",	--70
		x"fc",	--71
		x"40",	--72
		x"e5",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"e7",	--77
		x"40",	--78
		x"fc",	--79
		x"40",	--80
		x"e2",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"e7",	--85
		x"40",	--86
		x"fc",	--87
		x"40",	--88
		x"e3",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"e7",	--93
		x"40",	--94
		x"fc",	--95
		x"40",	--96
		x"e2",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"e7",	--101
		x"43",	--102
		x"43",	--103
		x"12",	--104
		x"e7",	--105
		x"43",	--106
		x"40",	--107
		x"4e",	--108
		x"40",	--109
		x"01",	--110
		x"41",	--111
		x"50",	--112
		x"00",	--113
		x"12",	--114
		x"e6",	--115
		x"41",	--116
		x"50",	--117
		x"00",	--118
		x"12",	--119
		x"e6",	--120
		x"43",	--121
		x"40",	--122
		x"4e",	--123
		x"40",	--124
		x"01",	--125
		x"41",	--126
		x"52",	--127
		x"12",	--128
		x"e6",	--129
		x"41",	--130
		x"52",	--131
		x"12",	--132
		x"e6",	--133
		x"41",	--134
		x"52",	--135
		x"41",	--136
		x"50",	--137
		x"00",	--138
		x"12",	--139
		x"e2",	--140
		x"40",	--141
		x"01",	--142
		x"41",	--143
		x"53",	--144
		x"12",	--145
		x"e9",	--146
		x"40",	--147
		x"01",	--148
		x"41",	--149
		x"12",	--150
		x"e9",	--151
		x"41",	--152
		x"41",	--153
		x"53",	--154
		x"12",	--155
		x"e3",	--156
		x"12",	--157
		x"e8",	--158
		x"43",	--159
		x"40",	--160
		x"e4",	--161
		x"12",	--162
		x"e8",	--163
		x"43",	--164
		x"43",	--165
		x"12",	--166
		x"e9",	--167
		x"40",	--168
		x"ff",	--169
		x"00",	--170
		x"d2",	--171
		x"43",	--172
		x"12",	--173
		x"ed",	--174
		x"93",	--175
		x"27",	--176
		x"12",	--177
		x"ed",	--178
		x"92",	--179
		x"24",	--180
		x"90",	--181
		x"00",	--182
		x"20",	--183
		x"12",	--184
		x"fc",	--185
		x"12",	--186
		x"eb",	--187
		x"53",	--188
		x"40",	--189
		x"00",	--190
		x"51",	--191
		x"5f",	--192
		x"43",	--193
		x"00",	--194
		x"4f",	--195
		x"41",	--196
		x"00",	--197
		x"12",	--198
		x"e8",	--199
		x"43",	--200
		x"3f",	--201
		x"93",	--202
		x"27",	--203
		x"53",	--204
		x"12",	--205
		x"fc",	--206
		x"12",	--207
		x"eb",	--208
		x"53",	--209
		x"3f",	--210
		x"90",	--211
		x"00",	--212
		x"2f",	--213
		x"93",	--214
		x"02",	--215
		x"24",	--216
		x"4f",	--217
		x"11",	--218
		x"12",	--219
		x"12",	--220
		x"fc",	--221
		x"4f",	--222
		x"00",	--223
		x"12",	--224
		x"eb",	--225
		x"52",	--226
		x"41",	--227
		x"00",	--228
		x"40",	--229
		x"00",	--230
		x"51",	--231
		x"5b",	--232
		x"4f",	--233
		x"00",	--234
		x"53",	--235
		x"3f",	--236
		x"40",	--237
		x"fb",	--238
		x"4e",	--239
		x"00",	--240
		x"4d",	--241
		x"00",	--242
		x"4c",	--243
		x"00",	--244
		x"43",	--245
		x"00",	--246
		x"43",	--247
		x"00",	--248
		x"43",	--249
		x"00",	--250
		x"41",	--251
		x"43",	--252
		x"00",	--253
		x"43",	--254
		x"00",	--255
		x"43",	--256
		x"00",	--257
		x"41",	--258
		x"4e",	--259
		x"00",	--260
		x"41",	--261
		x"4e",	--262
		x"00",	--263
		x"41",	--264
		x"4e",	--265
		x"00",	--266
		x"41",	--267
		x"4e",	--268
		x"00",	--269
		x"41",	--270
		x"4f",	--271
		x"00",	--272
		x"8e",	--273
		x"4d",	--274
		x"5f",	--275
		x"00",	--276
		x"4d",	--277
		x"00",	--278
		x"12",	--279
		x"c2",	--280
		x"43",	--281
		x"4e",	--282
		x"01",	--283
		x"4f",	--284
		x"01",	--285
		x"42",	--286
		x"01",	--287
		x"41",	--288
		x"12",	--289
		x"c2",	--290
		x"43",	--291
		x"4d",	--292
		x"01",	--293
		x"4f",	--294
		x"00",	--295
		x"01",	--296
		x"42",	--297
		x"01",	--298
		x"41",	--299
		x"5c",	--300
		x"8f",	--301
		x"00",	--302
		x"12",	--303
		x"c2",	--304
		x"43",	--305
		x"4e",	--306
		x"01",	--307
		x"4f",	--308
		x"00",	--309
		x"01",	--310
		x"42",	--311
		x"01",	--312
		x"41",	--313
		x"5d",	--314
		x"41",	--315
		x"40",	--316
		x"e0",	--317
		x"01",	--318
		x"40",	--319
		x"00",	--320
		x"01",	--321
		x"40",	--322
		x"02",	--323
		x"01",	--324
		x"12",	--325
		x"fb",	--326
		x"12",	--327
		x"eb",	--328
		x"43",	--329
		x"01",	--330
		x"40",	--331
		x"fb",	--332
		x"00",	--333
		x"12",	--334
		x"eb",	--335
		x"53",	--336
		x"43",	--337
		x"41",	--338
		x"12",	--339
		x"12",	--340
		x"43",	--341
		x"40",	--342
		x"3f",	--343
		x"4a",	--344
		x"4b",	--345
		x"42",	--346
		x"02",	--347
		x"12",	--348
		x"e7",	--349
		x"4a",	--350
		x"4b",	--351
		x"42",	--352
		x"02",	--353
		x"12",	--354
		x"e7",	--355
		x"12",	--356
		x"fb",	--357
		x"12",	--358
		x"eb",	--359
		x"53",	--360
		x"41",	--361
		x"41",	--362
		x"41",	--363
		x"4f",	--364
		x"02",	--365
		x"4e",	--366
		x"02",	--367
		x"41",	--368
		x"12",	--369
		x"12",	--370
		x"83",	--371
		x"4f",	--372
		x"4e",	--373
		x"93",	--374
		x"02",	--375
		x"24",	--376
		x"90",	--377
		x"00",	--378
		x"38",	--379
		x"20",	--380
		x"41",	--381
		x"4b",	--382
		x"00",	--383
		x"12",	--384
		x"e5",	--385
		x"4f",	--386
		x"41",	--387
		x"4b",	--388
		x"00",	--389
		x"12",	--390
		x"e5",	--391
		x"4f",	--392
		x"12",	--393
		x"12",	--394
		x"12",	--395
		x"fb",	--396
		x"12",	--397
		x"eb",	--398
		x"50",	--399
		x"00",	--400
		x"4a",	--401
		x"43",	--402
		x"12",	--403
		x"f5",	--404
		x"43",	--405
		x"40",	--406
		x"42",	--407
		x"12",	--408
		x"f3",	--409
		x"4e",	--410
		x"4f",	--411
		x"42",	--412
		x"02",	--413
		x"12",	--414
		x"e7",	--415
		x"4b",	--416
		x"43",	--417
		x"12",	--418
		x"f5",	--419
		x"43",	--420
		x"40",	--421
		x"42",	--422
		x"12",	--423
		x"f3",	--424
		x"4e",	--425
		x"4f",	--426
		x"42",	--427
		x"02",	--428
		x"12",	--429
		x"e7",	--430
		x"43",	--431
		x"53",	--432
		x"41",	--433
		x"41",	--434
		x"41",	--435
		x"41",	--436
		x"4b",	--437
		x"00",	--438
		x"12",	--439
		x"e5",	--440
		x"43",	--441
		x"4f",	--442
		x"42",	--443
		x"02",	--444
		x"12",	--445
		x"e9",	--446
		x"3f",	--447
		x"43",	--448
		x"40",	--449
		x"e2",	--450
		x"12",	--451
		x"e8",	--452
		x"4f",	--453
		x"02",	--454
		x"3f",	--455
		x"12",	--456
		x"fb",	--457
		x"12",	--458
		x"eb",	--459
		x"40",	--460
		x"fb",	--461
		x"00",	--462
		x"12",	--463
		x"eb",	--464
		x"4b",	--465
		x"00",	--466
		x"12",	--467
		x"fb",	--468
		x"12",	--469
		x"eb",	--470
		x"52",	--471
		x"43",	--472
		x"3f",	--473
		x"42",	--474
		x"02",	--475
		x"4f",	--476
		x"42",	--477
		x"02",	--478
		x"4f",	--479
		x"12",	--480
		x"12",	--481
		x"00",	--482
		x"12",	--483
		x"12",	--484
		x"00",	--485
		x"12",	--486
		x"fb",	--487
		x"12",	--488
		x"eb",	--489
		x"50",	--490
		x"00",	--491
		x"41",	--492
		x"4f",	--493
		x"02",	--494
		x"4e",	--495
		x"02",	--496
		x"41",	--497
		x"12",	--498
		x"12",	--499
		x"12",	--500
		x"83",	--501
		x"4f",	--502
		x"4e",	--503
		x"43",	--504
		x"00",	--505
		x"93",	--506
		x"24",	--507
		x"93",	--508
		x"02",	--509
		x"24",	--510
		x"43",	--511
		x"02",	--512
		x"41",	--513
		x"4b",	--514
		x"00",	--515
		x"12",	--516
		x"e5",	--517
		x"4f",	--518
		x"90",	--519
		x"00",	--520
		x"34",	--521
		x"43",	--522
		x"49",	--523
		x"42",	--524
		x"02",	--525
		x"12",	--526
		x"e9",	--527
		x"43",	--528
		x"53",	--529
		x"41",	--530
		x"41",	--531
		x"41",	--532
		x"41",	--533
		x"93",	--534
		x"02",	--535
		x"24",	--536
		x"43",	--537
		x"02",	--538
		x"42",	--539
		x"02",	--540
		x"12",	--541
		x"e9",	--542
		x"43",	--543
		x"53",	--544
		x"41",	--545
		x"41",	--546
		x"41",	--547
		x"41",	--548
		x"41",	--549
		x"4b",	--550
		x"00",	--551
		x"12",	--552
		x"e5",	--553
		x"4f",	--554
		x"3f",	--555
		x"43",	--556
		x"12",	--557
		x"e3",	--558
		x"43",	--559
		x"53",	--560
		x"41",	--561
		x"41",	--562
		x"41",	--563
		x"41",	--564
		x"43",	--565
		x"40",	--566
		x"e3",	--567
		x"12",	--568
		x"e8",	--569
		x"4f",	--570
		x"02",	--571
		x"3f",	--572
		x"43",	--573
		x"93",	--574
		x"02",	--575
		x"24",	--576
		x"43",	--577
		x"4f",	--578
		x"02",	--579
		x"43",	--580
		x"41",	--581
		x"42",	--582
		x"02",	--583
		x"92",	--584
		x"2c",	--585
		x"4e",	--586
		x"5f",	--587
		x"4f",	--588
		x"fb",	--589
		x"43",	--590
		x"00",	--591
		x"90",	--592
		x"00",	--593
		x"38",	--594
		x"43",	--595
		x"02",	--596
		x"41",	--597
		x"53",	--598
		x"4e",	--599
		x"02",	--600
		x"41",	--601
		x"40",	--602
		x"00",	--603
		x"00",	--604
		x"3f",	--605
		x"40",	--606
		x"00",	--607
		x"00",	--608
		x"3f",	--609
		x"42",	--610
		x"00",	--611
		x"3f",	--612
		x"40",	--613
		x"00",	--614
		x"00",	--615
		x"3f",	--616
		x"40",	--617
		x"00",	--618
		x"00",	--619
		x"3f",	--620
		x"40",	--621
		x"00",	--622
		x"00",	--623
		x"3f",	--624
		x"40",	--625
		x"00",	--626
		x"00",	--627
		x"3f",	--628
		x"42",	--629
		x"00",	--630
		x"4e",	--631
		x"be",	--632
		x"20",	--633
		x"df",	--634
		x"00",	--635
		x"41",	--636
		x"cf",	--637
		x"00",	--638
		x"41",	--639
		x"12",	--640
		x"12",	--641
		x"83",	--642
		x"4f",	--643
		x"4e",	--644
		x"12",	--645
		x"fc",	--646
		x"12",	--647
		x"eb",	--648
		x"53",	--649
		x"90",	--650
		x"00",	--651
		x"38",	--652
		x"41",	--653
		x"4b",	--654
		x"00",	--655
		x"12",	--656
		x"e5",	--657
		x"4f",	--658
		x"41",	--659
		x"4b",	--660
		x"00",	--661
		x"12",	--662
		x"e5",	--663
		x"4f",	--664
		x"12",	--665
		x"12",	--666
		x"12",	--667
		x"fc",	--668
		x"12",	--669
		x"eb",	--670
		x"50",	--671
		x"00",	--672
		x"4b",	--673
		x"00",	--674
		x"43",	--675
		x"53",	--676
		x"41",	--677
		x"41",	--678
		x"41",	--679
		x"12",	--680
		x"fc",	--681
		x"12",	--682
		x"eb",	--683
		x"40",	--684
		x"fc",	--685
		x"00",	--686
		x"12",	--687
		x"eb",	--688
		x"4b",	--689
		x"00",	--690
		x"12",	--691
		x"fc",	--692
		x"12",	--693
		x"eb",	--694
		x"52",	--695
		x"43",	--696
		x"3f",	--697
		x"12",	--698
		x"83",	--699
		x"4e",	--700
		x"93",	--701
		x"24",	--702
		x"38",	--703
		x"12",	--704
		x"fc",	--705
		x"12",	--706
		x"eb",	--707
		x"53",	--708
		x"41",	--709
		x"4b",	--710
		x"00",	--711
		x"12",	--712
		x"e5",	--713
		x"12",	--714
		x"12",	--715
		x"12",	--716
		x"fc",	--717
		x"12",	--718
		x"eb",	--719
		x"50",	--720
		x"00",	--721
		x"43",	--722
		x"53",	--723
		x"41",	--724
		x"41",	--725
		x"12",	--726
		x"fc",	--727
		x"12",	--728
		x"eb",	--729
		x"40",	--730
		x"fc",	--731
		x"00",	--732
		x"12",	--733
		x"eb",	--734
		x"4b",	--735
		x"00",	--736
		x"12",	--737
		x"fc",	--738
		x"12",	--739
		x"eb",	--740
		x"52",	--741
		x"43",	--742
		x"3f",	--743
		x"12",	--744
		x"12",	--745
		x"43",	--746
		x"00",	--747
		x"4f",	--748
		x"93",	--749
		x"24",	--750
		x"53",	--751
		x"43",	--752
		x"43",	--753
		x"3c",	--754
		x"90",	--755
		x"00",	--756
		x"2c",	--757
		x"5c",	--758
		x"5c",	--759
		x"5c",	--760
		x"5c",	--761
		x"11",	--762
		x"5d",	--763
		x"50",	--764
		x"ff",	--765
		x"43",	--766
		x"4f",	--767
		x"93",	--768
		x"24",	--769
		x"90",	--770
		x"00",	--771
		x"24",	--772
		x"4d",	--773
		x"50",	--774
		x"ff",	--775
		x"93",	--776
		x"23",	--777
		x"90",	--778
		x"00",	--779
		x"2c",	--780
		x"5c",	--781
		x"4c",	--782
		x"5b",	--783
		x"5b",	--784
		x"5b",	--785
		x"11",	--786
		x"5d",	--787
		x"50",	--788
		x"ff",	--789
		x"4f",	--790
		x"93",	--791
		x"23",	--792
		x"43",	--793
		x"00",	--794
		x"4c",	--795
		x"41",	--796
		x"41",	--797
		x"41",	--798
		x"43",	--799
		x"3f",	--800
		x"4d",	--801
		x"50",	--802
		x"ff",	--803
		x"90",	--804
		x"00",	--805
		x"2c",	--806
		x"5c",	--807
		x"5c",	--808
		x"5c",	--809
		x"5c",	--810
		x"11",	--811
		x"5d",	--812
		x"50",	--813
		x"ff",	--814
		x"43",	--815
		x"3f",	--816
		x"4d",	--817
		x"50",	--818
		x"ff",	--819
		x"90",	--820
		x"00",	--821
		x"2c",	--822
		x"5c",	--823
		x"5c",	--824
		x"5c",	--825
		x"5c",	--826
		x"11",	--827
		x"5d",	--828
		x"50",	--829
		x"ff",	--830
		x"43",	--831
		x"3f",	--832
		x"11",	--833
		x"12",	--834
		x"12",	--835
		x"fc",	--836
		x"12",	--837
		x"eb",	--838
		x"52",	--839
		x"43",	--840
		x"4c",	--841
		x"41",	--842
		x"41",	--843
		x"41",	--844
		x"43",	--845
		x"3f",	--846
		x"12",	--847
		x"12",	--848
		x"4e",	--849
		x"4c",	--850
		x"4e",	--851
		x"00",	--852
		x"4d",	--853
		x"00",	--854
		x"4c",	--855
		x"00",	--856
		x"4d",	--857
		x"43",	--858
		x"40",	--859
		x"36",	--860
		x"40",	--861
		x"01",	--862
		x"12",	--863
		x"fa",	--864
		x"4e",	--865
		x"00",	--866
		x"12",	--867
		x"c2",	--868
		x"43",	--869
		x"4a",	--870
		x"01",	--871
		x"40",	--872
		x"00",	--873
		x"01",	--874
		x"42",	--875
		x"01",	--876
		x"00",	--877
		x"41",	--878
		x"43",	--879
		x"41",	--880
		x"41",	--881
		x"41",	--882
		x"12",	--883
		x"12",	--884
		x"12",	--885
		x"43",	--886
		x"00",	--887
		x"40",	--888
		x"3f",	--889
		x"00",	--890
		x"4f",	--891
		x"4b",	--892
		x"00",	--893
		x"43",	--894
		x"12",	--895
		x"f5",	--896
		x"43",	--897
		x"40",	--898
		x"3f",	--899
		x"12",	--900
		x"f0",	--901
		x"4e",	--902
		x"4f",	--903
		x"4b",	--904
		x"00",	--905
		x"43",	--906
		x"12",	--907
		x"f5",	--908
		x"4e",	--909
		x"4f",	--910
		x"48",	--911
		x"49",	--912
		x"12",	--913
		x"f0",	--914
		x"12",	--915
		x"ed",	--916
		x"4e",	--917
		x"00",	--918
		x"43",	--919
		x"00",	--920
		x"41",	--921
		x"41",	--922
		x"41",	--923
		x"41",	--924
		x"12",	--925
		x"12",	--926
		x"12",	--927
		x"4d",	--928
		x"4e",	--929
		x"4d",	--930
		x"00",	--931
		x"4e",	--932
		x"00",	--933
		x"4f",	--934
		x"49",	--935
		x"00",	--936
		x"43",	--937
		x"12",	--938
		x"f5",	--939
		x"4e",	--940
		x"4f",	--941
		x"4a",	--942
		x"4b",	--943
		x"12",	--944
		x"f0",	--945
		x"4e",	--946
		x"4f",	--947
		x"49",	--948
		x"00",	--949
		x"43",	--950
		x"12",	--951
		x"f5",	--952
		x"4e",	--953
		x"4f",	--954
		x"4a",	--955
		x"4b",	--956
		x"12",	--957
		x"f0",	--958
		x"12",	--959
		x"ed",	--960
		x"4e",	--961
		x"00",	--962
		x"41",	--963
		x"41",	--964
		x"41",	--965
		x"41",	--966
		x"12",	--967
		x"12",	--968
		x"93",	--969
		x"02",	--970
		x"38",	--971
		x"40",	--972
		x"02",	--973
		x"43",	--974
		x"12",	--975
		x"4b",	--976
		x"ff",	--977
		x"11",	--978
		x"12",	--979
		x"12",	--980
		x"fc",	--981
		x"12",	--982
		x"eb",	--983
		x"50",	--984
		x"00",	--985
		x"53",	--986
		x"50",	--987
		x"00",	--988
		x"92",	--989
		x"02",	--990
		x"3b",	--991
		x"43",	--992
		x"41",	--993
		x"41",	--994
		x"41",	--995
		x"42",	--996
		x"02",	--997
		x"90",	--998
		x"00",	--999
		x"34",	--1000
		x"4e",	--1001
		x"5f",	--1002
		x"5e",	--1003
		x"5f",	--1004
		x"50",	--1005
		x"02",	--1006
		x"40",	--1007
		x"00",	--1008
		x"00",	--1009
		x"40",	--1010
		x"e7",	--1011
		x"00",	--1012
		x"40",	--1013
		x"02",	--1014
		x"00",	--1015
		x"53",	--1016
		x"4e",	--1017
		x"02",	--1018
		x"41",	--1019
		x"12",	--1020
		x"42",	--1021
		x"02",	--1022
		x"90",	--1023
		x"00",	--1024
		x"34",	--1025
		x"4b",	--1026
		x"5c",	--1027
		x"5b",	--1028
		x"5c",	--1029
		x"50",	--1030
		x"02",	--1031
		x"4f",	--1032
		x"00",	--1033
		x"4e",	--1034
		x"00",	--1035
		x"4d",	--1036
		x"00",	--1037
		x"53",	--1038
		x"4b",	--1039
		x"02",	--1040
		x"43",	--1041
		x"41",	--1042
		x"41",	--1043
		x"43",	--1044
		x"3f",	--1045
		x"12",	--1046
		x"50",	--1047
		x"ff",	--1048
		x"42",	--1049
		x"02",	--1050
		x"93",	--1051
		x"38",	--1052
		x"92",	--1053
		x"02",	--1054
		x"24",	--1055
		x"40",	--1056
		x"02",	--1057
		x"43",	--1058
		x"3c",	--1059
		x"50",	--1060
		x"00",	--1061
		x"9f",	--1062
		x"ff",	--1063
		x"24",	--1064
		x"53",	--1065
		x"9b",	--1066
		x"23",	--1067
		x"12",	--1068
		x"fc",	--1069
		x"12",	--1070
		x"eb",	--1071
		x"53",	--1072
		x"43",	--1073
		x"50",	--1074
		x"00",	--1075
		x"41",	--1076
		x"41",	--1077
		x"43",	--1078
		x"4e",	--1079
		x"00",	--1080
		x"4e",	--1081
		x"93",	--1082
		x"24",	--1083
		x"53",	--1084
		x"43",	--1085
		x"3c",	--1086
		x"4e",	--1087
		x"93",	--1088
		x"24",	--1089
		x"53",	--1090
		x"92",	--1091
		x"34",	--1092
		x"90",	--1093
		x"00",	--1094
		x"23",	--1095
		x"43",	--1096
		x"ff",	--1097
		x"4f",	--1098
		x"5d",	--1099
		x"51",	--1100
		x"4e",	--1101
		x"00",	--1102
		x"53",	--1103
		x"4e",	--1104
		x"93",	--1105
		x"23",	--1106
		x"4c",	--1107
		x"5e",	--1108
		x"5e",	--1109
		x"5c",	--1110
		x"50",	--1111
		x"02",	--1112
		x"41",	--1113
		x"12",	--1114
		x"00",	--1115
		x"50",	--1116
		x"00",	--1117
		x"41",	--1118
		x"41",	--1119
		x"43",	--1120
		x"3f",	--1121
		x"d0",	--1122
		x"02",	--1123
		x"01",	--1124
		x"40",	--1125
		x"0b",	--1126
		x"01",	--1127
		x"43",	--1128
		x"41",	--1129
		x"12",	--1130
		x"4f",	--1131
		x"42",	--1132
		x"02",	--1133
		x"90",	--1134
		x"00",	--1135
		x"34",	--1136
		x"4f",	--1137
		x"5c",	--1138
		x"4c",	--1139
		x"5d",	--1140
		x"5d",	--1141
		x"5d",	--1142
		x"8c",	--1143
		x"50",	--1144
		x"02",	--1145
		x"43",	--1146
		x"00",	--1147
		x"43",	--1148
		x"00",	--1149
		x"43",	--1150
		x"00",	--1151
		x"4b",	--1152
		x"00",	--1153
		x"4e",	--1154
		x"00",	--1155
		x"4f",	--1156
		x"53",	--1157
		x"4e",	--1158
		x"02",	--1159
		x"41",	--1160
		x"41",	--1161
		x"43",	--1162
		x"3f",	--1163
		x"5f",	--1164
		x"4f",	--1165
		x"5c",	--1166
		x"5c",	--1167
		x"5c",	--1168
		x"8f",	--1169
		x"50",	--1170
		x"02",	--1171
		x"43",	--1172
		x"00",	--1173
		x"4e",	--1174
		x"00",	--1175
		x"43",	--1176
		x"00",	--1177
		x"4d",	--1178
		x"00",	--1179
		x"43",	--1180
		x"00",	--1181
		x"43",	--1182
		x"41",	--1183
		x"5f",	--1184
		x"4f",	--1185
		x"5e",	--1186
		x"5e",	--1187
		x"5e",	--1188
		x"8f",	--1189
		x"43",	--1190
		x"02",	--1191
		x"43",	--1192
		x"41",	--1193
		x"12",	--1194
		x"12",	--1195
		x"12",	--1196
		x"12",	--1197
		x"12",	--1198
		x"12",	--1199
		x"12",	--1200
		x"12",	--1201
		x"12",	--1202
		x"93",	--1203
		x"02",	--1204
		x"38",	--1205
		x"40",	--1206
		x"02",	--1207
		x"4a",	--1208
		x"53",	--1209
		x"4a",	--1210
		x"52",	--1211
		x"4a",	--1212
		x"50",	--1213
		x"00",	--1214
		x"43",	--1215
		x"3c",	--1216
		x"53",	--1217
		x"4f",	--1218
		x"00",	--1219
		x"53",	--1220
		x"50",	--1221
		x"00",	--1222
		x"50",	--1223
		x"00",	--1224
		x"50",	--1225
		x"00",	--1226
		x"50",	--1227
		x"00",	--1228
		x"92",	--1229
		x"02",	--1230
		x"34",	--1231
		x"93",	--1232
		x"00",	--1233
		x"27",	--1234
		x"4b",	--1235
		x"9b",	--1236
		x"00",	--1237
		x"2b",	--1238
		x"43",	--1239
		x"00",	--1240
		x"4b",	--1241
		x"00",	--1242
		x"12",	--1243
		x"00",	--1244
		x"93",	--1245
		x"00",	--1246
		x"27",	--1247
		x"47",	--1248
		x"53",	--1249
		x"4f",	--1250
		x"00",	--1251
		x"98",	--1252
		x"2b",	--1253
		x"43",	--1254
		x"00",	--1255
		x"3f",	--1256
		x"f0",	--1257
		x"ff",	--1258
		x"01",	--1259
		x"41",	--1260
		x"41",	--1261
		x"41",	--1262
		x"41",	--1263
		x"41",	--1264
		x"41",	--1265
		x"41",	--1266
		x"41",	--1267
		x"41",	--1268
		x"13",	--1269
		x"4e",	--1270
		x"00",	--1271
		x"43",	--1272
		x"41",	--1273
		x"4f",	--1274
		x"4f",	--1275
		x"41",	--1276
		x"42",	--1277
		x"00",	--1278
		x"f2",	--1279
		x"23",	--1280
		x"4f",	--1281
		x"00",	--1282
		x"43",	--1283
		x"41",	--1284
		x"f0",	--1285
		x"00",	--1286
		x"4f",	--1287
		x"fd",	--1288
		x"11",	--1289
		x"12",	--1290
		x"e9",	--1291
		x"41",	--1292
		x"12",	--1293
		x"4f",	--1294
		x"4f",	--1295
		x"11",	--1296
		x"11",	--1297
		x"11",	--1298
		x"11",	--1299
		x"4e",	--1300
		x"12",	--1301
		x"ea",	--1302
		x"4b",	--1303
		x"12",	--1304
		x"ea",	--1305
		x"41",	--1306
		x"41",	--1307
		x"12",	--1308
		x"12",	--1309
		x"4f",	--1310
		x"40",	--1311
		x"00",	--1312
		x"4a",	--1313
		x"4b",	--1314
		x"f0",	--1315
		x"00",	--1316
		x"24",	--1317
		x"11",	--1318
		x"53",	--1319
		x"23",	--1320
		x"f3",	--1321
		x"24",	--1322
		x"40",	--1323
		x"00",	--1324
		x"12",	--1325
		x"e9",	--1326
		x"53",	--1327
		x"93",	--1328
		x"23",	--1329
		x"41",	--1330
		x"41",	--1331
		x"41",	--1332
		x"40",	--1333
		x"00",	--1334
		x"3f",	--1335
		x"12",	--1336
		x"4f",	--1337
		x"4f",	--1338
		x"10",	--1339
		x"11",	--1340
		x"4e",	--1341
		x"12",	--1342
		x"ea",	--1343
		x"4b",	--1344
		x"12",	--1345
		x"ea",	--1346
		x"41",	--1347
		x"41",	--1348
		x"12",	--1349
		x"12",	--1350
		x"4e",	--1351
		x"4f",	--1352
		x"4f",	--1353
		x"10",	--1354
		x"11",	--1355
		x"4d",	--1356
		x"12",	--1357
		x"ea",	--1358
		x"4b",	--1359
		x"12",	--1360
		x"ea",	--1361
		x"4b",	--1362
		x"4a",	--1363
		x"10",	--1364
		x"10",	--1365
		x"ec",	--1366
		x"ec",	--1367
		x"4d",	--1368
		x"12",	--1369
		x"ea",	--1370
		x"4a",	--1371
		x"12",	--1372
		x"ea",	--1373
		x"41",	--1374
		x"41",	--1375
		x"41",	--1376
		x"12",	--1377
		x"12",	--1378
		x"12",	--1379
		x"4f",	--1380
		x"93",	--1381
		x"24",	--1382
		x"4e",	--1383
		x"53",	--1384
		x"43",	--1385
		x"4a",	--1386
		x"5b",	--1387
		x"4d",	--1388
		x"11",	--1389
		x"12",	--1390
		x"ea",	--1391
		x"99",	--1392
		x"24",	--1393
		x"53",	--1394
		x"b0",	--1395
		x"00",	--1396
		x"20",	--1397
		x"40",	--1398
		x"00",	--1399
		x"12",	--1400
		x"e9",	--1401
		x"3f",	--1402
		x"40",	--1403
		x"00",	--1404
		x"12",	--1405
		x"e9",	--1406
		x"3f",	--1407
		x"41",	--1408
		x"41",	--1409
		x"41",	--1410
		x"41",	--1411
		x"12",	--1412
		x"12",	--1413
		x"12",	--1414
		x"4f",	--1415
		x"93",	--1416
		x"24",	--1417
		x"4e",	--1418
		x"53",	--1419
		x"43",	--1420
		x"4a",	--1421
		x"11",	--1422
		x"12",	--1423
		x"ea",	--1424
		x"99",	--1425
		x"24",	--1426
		x"53",	--1427
		x"b0",	--1428
		x"00",	--1429
		x"23",	--1430
		x"40",	--1431
		x"00",	--1432
		x"12",	--1433
		x"e9",	--1434
		x"4a",	--1435
		x"11",	--1436
		x"12",	--1437
		x"ea",	--1438
		x"99",	--1439
		x"23",	--1440
		x"41",	--1441
		x"41",	--1442
		x"41",	--1443
		x"41",	--1444
		x"12",	--1445
		x"12",	--1446
		x"12",	--1447
		x"50",	--1448
		x"ff",	--1449
		x"4f",	--1450
		x"93",	--1451
		x"38",	--1452
		x"90",	--1453
		x"00",	--1454
		x"38",	--1455
		x"43",	--1456
		x"41",	--1457
		x"59",	--1458
		x"40",	--1459
		x"00",	--1460
		x"4b",	--1461
		x"12",	--1462
		x"fa",	--1463
		x"50",	--1464
		x"00",	--1465
		x"4f",	--1466
		x"00",	--1467
		x"53",	--1468
		x"40",	--1469
		x"00",	--1470
		x"4b",	--1471
		x"12",	--1472
		x"fa",	--1473
		x"4f",	--1474
		x"90",	--1475
		x"00",	--1476
		x"37",	--1477
		x"49",	--1478
		x"53",	--1479
		x"51",	--1480
		x"40",	--1481
		x"00",	--1482
		x"4b",	--1483
		x"12",	--1484
		x"fa",	--1485
		x"50",	--1486
		x"00",	--1487
		x"4f",	--1488
		x"00",	--1489
		x"53",	--1490
		x"41",	--1491
		x"5a",	--1492
		x"4f",	--1493
		x"11",	--1494
		x"12",	--1495
		x"e9",	--1496
		x"93",	--1497
		x"23",	--1498
		x"50",	--1499
		x"00",	--1500
		x"41",	--1501
		x"41",	--1502
		x"41",	--1503
		x"41",	--1504
		x"40",	--1505
		x"00",	--1506
		x"12",	--1507
		x"e9",	--1508
		x"e3",	--1509
		x"53",	--1510
		x"3f",	--1511
		x"43",	--1512
		x"43",	--1513
		x"3f",	--1514
		x"12",	--1515
		x"12",	--1516
		x"12",	--1517
		x"41",	--1518
		x"52",	--1519
		x"4b",	--1520
		x"49",	--1521
		x"93",	--1522
		x"20",	--1523
		x"3c",	--1524
		x"11",	--1525
		x"12",	--1526
		x"e9",	--1527
		x"49",	--1528
		x"4a",	--1529
		x"53",	--1530
		x"4a",	--1531
		x"00",	--1532
		x"93",	--1533
		x"24",	--1534
		x"90",	--1535
		x"00",	--1536
		x"23",	--1537
		x"49",	--1538
		x"53",	--1539
		x"49",	--1540
		x"00",	--1541
		x"50",	--1542
		x"ff",	--1543
		x"90",	--1544
		x"00",	--1545
		x"2f",	--1546
		x"4f",	--1547
		x"5f",	--1548
		x"4f",	--1549
		x"fc",	--1550
		x"41",	--1551
		x"41",	--1552
		x"41",	--1553
		x"41",	--1554
		x"4b",	--1555
		x"52",	--1556
		x"4b",	--1557
		x"00",	--1558
		x"4b",	--1559
		x"12",	--1560
		x"ea",	--1561
		x"49",	--1562
		x"3f",	--1563
		x"4b",	--1564
		x"53",	--1565
		x"4b",	--1566
		x"12",	--1567
		x"ea",	--1568
		x"49",	--1569
		x"3f",	--1570
		x"4b",	--1571
		x"53",	--1572
		x"4f",	--1573
		x"49",	--1574
		x"93",	--1575
		x"27",	--1576
		x"53",	--1577
		x"11",	--1578
		x"12",	--1579
		x"e9",	--1580
		x"49",	--1581
		x"93",	--1582
		x"23",	--1583
		x"3f",	--1584
		x"4b",	--1585
		x"52",	--1586
		x"4b",	--1587
		x"00",	--1588
		x"4b",	--1589
		x"12",	--1590
		x"eb",	--1591
		x"49",	--1592
		x"3f",	--1593
		x"4b",	--1594
		x"53",	--1595
		x"4b",	--1596
		x"4e",	--1597
		x"10",	--1598
		x"11",	--1599
		x"10",	--1600
		x"11",	--1601
		x"12",	--1602
		x"ea",	--1603
		x"49",	--1604
		x"3f",	--1605
		x"4b",	--1606
		x"53",	--1607
		x"4b",	--1608
		x"12",	--1609
		x"eb",	--1610
		x"49",	--1611
		x"3f",	--1612
		x"4b",	--1613
		x"53",	--1614
		x"4b",	--1615
		x"12",	--1616
		x"e9",	--1617
		x"49",	--1618
		x"3f",	--1619
		x"4b",	--1620
		x"53",	--1621
		x"4b",	--1622
		x"12",	--1623
		x"ea",	--1624
		x"49",	--1625
		x"3f",	--1626
		x"4b",	--1627
		x"53",	--1628
		x"4b",	--1629
		x"12",	--1630
		x"ea",	--1631
		x"49",	--1632
		x"3f",	--1633
		x"40",	--1634
		x"00",	--1635
		x"12",	--1636
		x"e9",	--1637
		x"3f",	--1638
		x"12",	--1639
		x"12",	--1640
		x"42",	--1641
		x"02",	--1642
		x"42",	--1643
		x"00",	--1644
		x"04",	--1645
		x"42",	--1646
		x"02",	--1647
		x"90",	--1648
		x"00",	--1649
		x"34",	--1650
		x"53",	--1651
		x"02",	--1652
		x"42",	--1653
		x"02",	--1654
		x"42",	--1655
		x"02",	--1656
		x"9f",	--1657
		x"20",	--1658
		x"53",	--1659
		x"02",	--1660
		x"40",	--1661
		x"00",	--1662
		x"00",	--1663
		x"41",	--1664
		x"41",	--1665
		x"c0",	--1666
		x"00",	--1667
		x"00",	--1668
		x"13",	--1669
		x"43",	--1670
		x"02",	--1671
		x"3f",	--1672
		x"4e",	--1673
		x"4f",	--1674
		x"40",	--1675
		x"36",	--1676
		x"40",	--1677
		x"01",	--1678
		x"12",	--1679
		x"fa",	--1680
		x"53",	--1681
		x"4e",	--1682
		x"00",	--1683
		x"40",	--1684
		x"00",	--1685
		x"00",	--1686
		x"41",	--1687
		x"42",	--1688
		x"02",	--1689
		x"42",	--1690
		x"02",	--1691
		x"9f",	--1692
		x"38",	--1693
		x"42",	--1694
		x"02",	--1695
		x"82",	--1696
		x"02",	--1697
		x"41",	--1698
		x"42",	--1699
		x"02",	--1700
		x"42",	--1701
		x"02",	--1702
		x"40",	--1703
		x"00",	--1704
		x"8d",	--1705
		x"8e",	--1706
		x"41",	--1707
		x"42",	--1708
		x"02",	--1709
		x"4f",	--1710
		x"04",	--1711
		x"42",	--1712
		x"02",	--1713
		x"42",	--1714
		x"02",	--1715
		x"9e",	--1716
		x"24",	--1717
		x"42",	--1718
		x"02",	--1719
		x"90",	--1720
		x"00",	--1721
		x"38",	--1722
		x"43",	--1723
		x"02",	--1724
		x"41",	--1725
		x"53",	--1726
		x"02",	--1727
		x"41",	--1728
		x"43",	--1729
		x"41",	--1730
		x"12",	--1731
		x"12",	--1732
		x"4e",	--1733
		x"4f",	--1734
		x"43",	--1735
		x"40",	--1736
		x"4f",	--1737
		x"12",	--1738
		x"f4",	--1739
		x"93",	--1740
		x"34",	--1741
		x"4a",	--1742
		x"4b",	--1743
		x"12",	--1744
		x"f4",	--1745
		x"41",	--1746
		x"41",	--1747
		x"41",	--1748
		x"43",	--1749
		x"40",	--1750
		x"4f",	--1751
		x"4a",	--1752
		x"4b",	--1753
		x"12",	--1754
		x"f0",	--1755
		x"12",	--1756
		x"f4",	--1757
		x"53",	--1758
		x"60",	--1759
		x"80",	--1760
		x"41",	--1761
		x"41",	--1762
		x"41",	--1763
		x"12",	--1764
		x"12",	--1765
		x"12",	--1766
		x"12",	--1767
		x"12",	--1768
		x"12",	--1769
		x"12",	--1770
		x"12",	--1771
		x"50",	--1772
		x"ff",	--1773
		x"4d",	--1774
		x"4f",	--1775
		x"93",	--1776
		x"28",	--1777
		x"4e",	--1778
		x"93",	--1779
		x"28",	--1780
		x"92",	--1781
		x"20",	--1782
		x"40",	--1783
		x"f0",	--1784
		x"92",	--1785
		x"24",	--1786
		x"93",	--1787
		x"24",	--1788
		x"93",	--1789
		x"24",	--1790
		x"4f",	--1791
		x"00",	--1792
		x"00",	--1793
		x"4e",	--1794
		x"00",	--1795
		x"4f",	--1796
		x"00",	--1797
		x"4f",	--1798
		x"00",	--1799
		x"4e",	--1800
		x"00",	--1801
		x"4e",	--1802
		x"00",	--1803
		x"41",	--1804
		x"8b",	--1805
		x"4c",	--1806
		x"93",	--1807
		x"38",	--1808
		x"90",	--1809
		x"00",	--1810
		x"34",	--1811
		x"93",	--1812
		x"38",	--1813
		x"46",	--1814
		x"00",	--1815
		x"47",	--1816
		x"00",	--1817
		x"49",	--1818
		x"f0",	--1819
		x"00",	--1820
		x"24",	--1821
		x"46",	--1822
		x"47",	--1823
		x"c3",	--1824
		x"10",	--1825
		x"10",	--1826
		x"53",	--1827
		x"23",	--1828
		x"4a",	--1829
		x"00",	--1830
		x"4b",	--1831
		x"00",	--1832
		x"43",	--1833
		x"43",	--1834
		x"f0",	--1835
		x"00",	--1836
		x"24",	--1837
		x"5c",	--1838
		x"6d",	--1839
		x"53",	--1840
		x"23",	--1841
		x"53",	--1842
		x"63",	--1843
		x"f6",	--1844
		x"f7",	--1845
		x"43",	--1846
		x"43",	--1847
		x"93",	--1848
		x"20",	--1849
		x"93",	--1850
		x"24",	--1851
		x"41",	--1852
		x"00",	--1853
		x"41",	--1854
		x"00",	--1855
		x"da",	--1856
		x"db",	--1857
		x"4f",	--1858
		x"00",	--1859
		x"9e",	--1860
		x"00",	--1861
		x"20",	--1862
		x"4f",	--1863
		x"00",	--1864
		x"41",	--1865
		x"00",	--1866
		x"46",	--1867
		x"47",	--1868
		x"54",	--1869
		x"65",	--1870
		x"4e",	--1871
		x"00",	--1872
		x"4f",	--1873
		x"00",	--1874
		x"40",	--1875
		x"00",	--1876
		x"00",	--1877
		x"93",	--1878
		x"38",	--1879
		x"48",	--1880
		x"50",	--1881
		x"00",	--1882
		x"41",	--1883
		x"41",	--1884
		x"41",	--1885
		x"41",	--1886
		x"41",	--1887
		x"41",	--1888
		x"41",	--1889
		x"41",	--1890
		x"41",	--1891
		x"91",	--1892
		x"38",	--1893
		x"4b",	--1894
		x"00",	--1895
		x"43",	--1896
		x"43",	--1897
		x"4f",	--1898
		x"00",	--1899
		x"9e",	--1900
		x"00",	--1901
		x"27",	--1902
		x"93",	--1903
		x"24",	--1904
		x"46",	--1905
		x"47",	--1906
		x"84",	--1907
		x"75",	--1908
		x"93",	--1909
		x"38",	--1910
		x"43",	--1911
		x"00",	--1912
		x"41",	--1913
		x"00",	--1914
		x"4e",	--1915
		x"00",	--1916
		x"4f",	--1917
		x"00",	--1918
		x"4e",	--1919
		x"4f",	--1920
		x"53",	--1921
		x"63",	--1922
		x"90",	--1923
		x"3f",	--1924
		x"28",	--1925
		x"90",	--1926
		x"40",	--1927
		x"2c",	--1928
		x"93",	--1929
		x"2c",	--1930
		x"48",	--1931
		x"00",	--1932
		x"53",	--1933
		x"5e",	--1934
		x"6f",	--1935
		x"4b",	--1936
		x"53",	--1937
		x"4e",	--1938
		x"4f",	--1939
		x"53",	--1940
		x"63",	--1941
		x"90",	--1942
		x"3f",	--1943
		x"2b",	--1944
		x"24",	--1945
		x"4e",	--1946
		x"00",	--1947
		x"4f",	--1948
		x"00",	--1949
		x"4a",	--1950
		x"00",	--1951
		x"40",	--1952
		x"00",	--1953
		x"00",	--1954
		x"93",	--1955
		x"37",	--1956
		x"4e",	--1957
		x"4f",	--1958
		x"f3",	--1959
		x"f3",	--1960
		x"c3",	--1961
		x"10",	--1962
		x"10",	--1963
		x"4c",	--1964
		x"4d",	--1965
		x"de",	--1966
		x"df",	--1967
		x"4a",	--1968
		x"00",	--1969
		x"4b",	--1970
		x"00",	--1971
		x"53",	--1972
		x"00",	--1973
		x"48",	--1974
		x"3f",	--1975
		x"93",	--1976
		x"23",	--1977
		x"4f",	--1978
		x"00",	--1979
		x"4f",	--1980
		x"00",	--1981
		x"00",	--1982
		x"4f",	--1983
		x"00",	--1984
		x"00",	--1985
		x"4f",	--1986
		x"00",	--1987
		x"00",	--1988
		x"4e",	--1989
		x"00",	--1990
		x"ff",	--1991
		x"00",	--1992
		x"4e",	--1993
		x"00",	--1994
		x"4d",	--1995
		x"3f",	--1996
		x"43",	--1997
		x"43",	--1998
		x"3f",	--1999
		x"e3",	--2000
		x"53",	--2001
		x"90",	--2002
		x"00",	--2003
		x"37",	--2004
		x"3f",	--2005
		x"93",	--2006
		x"2b",	--2007
		x"3f",	--2008
		x"44",	--2009
		x"45",	--2010
		x"86",	--2011
		x"77",	--2012
		x"3f",	--2013
		x"4e",	--2014
		x"3f",	--2015
		x"43",	--2016
		x"00",	--2017
		x"41",	--2018
		x"00",	--2019
		x"e3",	--2020
		x"e3",	--2021
		x"53",	--2022
		x"63",	--2023
		x"4e",	--2024
		x"00",	--2025
		x"4f",	--2026
		x"00",	--2027
		x"3f",	--2028
		x"93",	--2029
		x"27",	--2030
		x"59",	--2031
		x"00",	--2032
		x"44",	--2033
		x"00",	--2034
		x"45",	--2035
		x"00",	--2036
		x"49",	--2037
		x"f0",	--2038
		x"00",	--2039
		x"24",	--2040
		x"4d",	--2041
		x"44",	--2042
		x"45",	--2043
		x"c3",	--2044
		x"10",	--2045
		x"10",	--2046
		x"53",	--2047
		x"23",	--2048
		x"4c",	--2049
		x"00",	--2050
		x"4d",	--2051
		x"00",	--2052
		x"43",	--2053
		x"43",	--2054
		x"f0",	--2055
		x"00",	--2056
		x"24",	--2057
		x"5c",	--2058
		x"6d",	--2059
		x"53",	--2060
		x"23",	--2061
		x"53",	--2062
		x"63",	--2063
		x"f4",	--2064
		x"f5",	--2065
		x"43",	--2066
		x"43",	--2067
		x"93",	--2068
		x"20",	--2069
		x"93",	--2070
		x"20",	--2071
		x"43",	--2072
		x"43",	--2073
		x"41",	--2074
		x"00",	--2075
		x"41",	--2076
		x"00",	--2077
		x"da",	--2078
		x"db",	--2079
		x"3f",	--2080
		x"43",	--2081
		x"43",	--2082
		x"3f",	--2083
		x"92",	--2084
		x"23",	--2085
		x"9e",	--2086
		x"00",	--2087
		x"00",	--2088
		x"27",	--2089
		x"40",	--2090
		x"fd",	--2091
		x"3f",	--2092
		x"50",	--2093
		x"ff",	--2094
		x"4e",	--2095
		x"00",	--2096
		x"4f",	--2097
		x"00",	--2098
		x"4c",	--2099
		x"00",	--2100
		x"4d",	--2101
		x"00",	--2102
		x"41",	--2103
		x"50",	--2104
		x"00",	--2105
		x"41",	--2106
		x"52",	--2107
		x"12",	--2108
		x"f8",	--2109
		x"41",	--2110
		x"50",	--2111
		x"00",	--2112
		x"41",	--2113
		x"12",	--2114
		x"f8",	--2115
		x"41",	--2116
		x"52",	--2117
		x"41",	--2118
		x"50",	--2119
		x"00",	--2120
		x"41",	--2121
		x"50",	--2122
		x"00",	--2123
		x"12",	--2124
		x"ed",	--2125
		x"12",	--2126
		x"f6",	--2127
		x"50",	--2128
		x"00",	--2129
		x"41",	--2130
		x"50",	--2131
		x"ff",	--2132
		x"4e",	--2133
		x"00",	--2134
		x"4f",	--2135
		x"00",	--2136
		x"4c",	--2137
		x"00",	--2138
		x"4d",	--2139
		x"00",	--2140
		x"41",	--2141
		x"50",	--2142
		x"00",	--2143
		x"41",	--2144
		x"52",	--2145
		x"12",	--2146
		x"f8",	--2147
		x"41",	--2148
		x"50",	--2149
		x"00",	--2150
		x"41",	--2151
		x"12",	--2152
		x"f8",	--2153
		x"e3",	--2154
		x"00",	--2155
		x"41",	--2156
		x"52",	--2157
		x"41",	--2158
		x"50",	--2159
		x"00",	--2160
		x"41",	--2161
		x"50",	--2162
		x"00",	--2163
		x"12",	--2164
		x"ed",	--2165
		x"12",	--2166
		x"f6",	--2167
		x"50",	--2168
		x"00",	--2169
		x"41",	--2170
		x"12",	--2171
		x"12",	--2172
		x"12",	--2173
		x"12",	--2174
		x"12",	--2175
		x"12",	--2176
		x"12",	--2177
		x"12",	--2178
		x"50",	--2179
		x"ff",	--2180
		x"4e",	--2181
		x"00",	--2182
		x"4f",	--2183
		x"00",	--2184
		x"4c",	--2185
		x"00",	--2186
		x"4d",	--2187
		x"00",	--2188
		x"41",	--2189
		x"50",	--2190
		x"00",	--2191
		x"41",	--2192
		x"52",	--2193
		x"12",	--2194
		x"f8",	--2195
		x"41",	--2196
		x"50",	--2197
		x"00",	--2198
		x"41",	--2199
		x"12",	--2200
		x"f8",	--2201
		x"41",	--2202
		x"00",	--2203
		x"93",	--2204
		x"28",	--2205
		x"41",	--2206
		x"00",	--2207
		x"93",	--2208
		x"28",	--2209
		x"92",	--2210
		x"24",	--2211
		x"92",	--2212
		x"24",	--2213
		x"93",	--2214
		x"24",	--2215
		x"93",	--2216
		x"24",	--2217
		x"41",	--2218
		x"00",	--2219
		x"41",	--2220
		x"00",	--2221
		x"41",	--2222
		x"00",	--2223
		x"41",	--2224
		x"00",	--2225
		x"40",	--2226
		x"00",	--2227
		x"43",	--2228
		x"43",	--2229
		x"43",	--2230
		x"43",	--2231
		x"43",	--2232
		x"00",	--2233
		x"43",	--2234
		x"00",	--2235
		x"43",	--2236
		x"43",	--2237
		x"4c",	--2238
		x"00",	--2239
		x"3c",	--2240
		x"58",	--2241
		x"69",	--2242
		x"c3",	--2243
		x"10",	--2244
		x"10",	--2245
		x"53",	--2246
		x"00",	--2247
		x"24",	--2248
		x"b3",	--2249
		x"24",	--2250
		x"58",	--2251
		x"69",	--2252
		x"56",	--2253
		x"67",	--2254
		x"43",	--2255
		x"43",	--2256
		x"99",	--2257
		x"28",	--2258
		x"24",	--2259
		x"43",	--2260
		x"43",	--2261
		x"5c",	--2262
		x"6d",	--2263
		x"56",	--2264
		x"67",	--2265
		x"93",	--2266
		x"37",	--2267
		x"d3",	--2268
		x"d3",	--2269
		x"3f",	--2270
		x"98",	--2271
		x"2b",	--2272
		x"3f",	--2273
		x"4a",	--2274
		x"00",	--2275
		x"4b",	--2276
		x"00",	--2277
		x"4f",	--2278
		x"41",	--2279
		x"00",	--2280
		x"51",	--2281
		x"00",	--2282
		x"4a",	--2283
		x"53",	--2284
		x"46",	--2285
		x"00",	--2286
		x"43",	--2287
		x"91",	--2288
		x"00",	--2289
		x"00",	--2290
		x"24",	--2291
		x"4d",	--2292
		x"00",	--2293
		x"93",	--2294
		x"38",	--2295
		x"90",	--2296
		x"40",	--2297
		x"2c",	--2298
		x"41",	--2299
		x"00",	--2300
		x"53",	--2301
		x"41",	--2302
		x"00",	--2303
		x"41",	--2304
		x"00",	--2305
		x"4d",	--2306
		x"5e",	--2307
		x"6f",	--2308
		x"93",	--2309
		x"38",	--2310
		x"5a",	--2311
		x"6b",	--2312
		x"53",	--2313
		x"90",	--2314
		x"40",	--2315
		x"2b",	--2316
		x"4a",	--2317
		x"00",	--2318
		x"4b",	--2319
		x"00",	--2320
		x"4c",	--2321
		x"00",	--2322
		x"4e",	--2323
		x"4f",	--2324
		x"f0",	--2325
		x"00",	--2326
		x"f3",	--2327
		x"90",	--2328
		x"00",	--2329
		x"24",	--2330
		x"4e",	--2331
		x"00",	--2332
		x"4f",	--2333
		x"00",	--2334
		x"40",	--2335
		x"00",	--2336
		x"00",	--2337
		x"41",	--2338
		x"52",	--2339
		x"12",	--2340
		x"f6",	--2341
		x"50",	--2342
		x"00",	--2343
		x"41",	--2344
		x"41",	--2345
		x"41",	--2346
		x"41",	--2347
		x"41",	--2348
		x"41",	--2349
		x"41",	--2350
		x"41",	--2351
		x"41",	--2352
		x"d3",	--2353
		x"d3",	--2354
		x"3f",	--2355
		x"50",	--2356
		x"00",	--2357
		x"4a",	--2358
		x"b3",	--2359
		x"24",	--2360
		x"41",	--2361
		x"00",	--2362
		x"41",	--2363
		x"00",	--2364
		x"c3",	--2365
		x"10",	--2366
		x"10",	--2367
		x"4c",	--2368
		x"4d",	--2369
		x"d3",	--2370
		x"d0",	--2371
		x"80",	--2372
		x"46",	--2373
		x"00",	--2374
		x"47",	--2375
		x"00",	--2376
		x"c3",	--2377
		x"10",	--2378
		x"10",	--2379
		x"53",	--2380
		x"93",	--2381
		x"3b",	--2382
		x"48",	--2383
		x"00",	--2384
		x"3f",	--2385
		x"93",	--2386
		x"24",	--2387
		x"43",	--2388
		x"91",	--2389
		x"00",	--2390
		x"00",	--2391
		x"24",	--2392
		x"4f",	--2393
		x"00",	--2394
		x"41",	--2395
		x"50",	--2396
		x"00",	--2397
		x"3f",	--2398
		x"93",	--2399
		x"23",	--2400
		x"4e",	--2401
		x"4f",	--2402
		x"f0",	--2403
		x"00",	--2404
		x"f3",	--2405
		x"93",	--2406
		x"23",	--2407
		x"93",	--2408
		x"23",	--2409
		x"93",	--2410
		x"00",	--2411
		x"20",	--2412
		x"93",	--2413
		x"00",	--2414
		x"27",	--2415
		x"50",	--2416
		x"00",	--2417
		x"63",	--2418
		x"f0",	--2419
		x"ff",	--2420
		x"f3",	--2421
		x"3f",	--2422
		x"43",	--2423
		x"3f",	--2424
		x"43",	--2425
		x"3f",	--2426
		x"43",	--2427
		x"91",	--2428
		x"00",	--2429
		x"00",	--2430
		x"24",	--2431
		x"4f",	--2432
		x"00",	--2433
		x"41",	--2434
		x"50",	--2435
		x"00",	--2436
		x"3f",	--2437
		x"43",	--2438
		x"3f",	--2439
		x"93",	--2440
		x"23",	--2441
		x"40",	--2442
		x"fd",	--2443
		x"3f",	--2444
		x"12",	--2445
		x"12",	--2446
		x"12",	--2447
		x"12",	--2448
		x"12",	--2449
		x"50",	--2450
		x"ff",	--2451
		x"4e",	--2452
		x"00",	--2453
		x"4f",	--2454
		x"00",	--2455
		x"4c",	--2456
		x"00",	--2457
		x"4d",	--2458
		x"00",	--2459
		x"41",	--2460
		x"50",	--2461
		x"00",	--2462
		x"41",	--2463
		x"52",	--2464
		x"12",	--2465
		x"f8",	--2466
		x"41",	--2467
		x"52",	--2468
		x"41",	--2469
		x"12",	--2470
		x"f8",	--2471
		x"41",	--2472
		x"00",	--2473
		x"93",	--2474
		x"28",	--2475
		x"41",	--2476
		x"00",	--2477
		x"93",	--2478
		x"28",	--2479
		x"e1",	--2480
		x"00",	--2481
		x"00",	--2482
		x"92",	--2483
		x"24",	--2484
		x"93",	--2485
		x"24",	--2486
		x"92",	--2487
		x"24",	--2488
		x"93",	--2489
		x"24",	--2490
		x"41",	--2491
		x"00",	--2492
		x"81",	--2493
		x"00",	--2494
		x"4d",	--2495
		x"00",	--2496
		x"41",	--2497
		x"00",	--2498
		x"41",	--2499
		x"00",	--2500
		x"41",	--2501
		x"00",	--2502
		x"41",	--2503
		x"00",	--2504
		x"99",	--2505
		x"2c",	--2506
		x"5e",	--2507
		x"6f",	--2508
		x"53",	--2509
		x"4d",	--2510
		x"00",	--2511
		x"40",	--2512
		x"00",	--2513
		x"43",	--2514
		x"40",	--2515
		x"40",	--2516
		x"43",	--2517
		x"43",	--2518
		x"3c",	--2519
		x"dc",	--2520
		x"dd",	--2521
		x"88",	--2522
		x"79",	--2523
		x"c3",	--2524
		x"10",	--2525
		x"10",	--2526
		x"5e",	--2527
		x"6f",	--2528
		x"53",	--2529
		x"24",	--2530
		x"99",	--2531
		x"2b",	--2532
		x"23",	--2533
		x"98",	--2534
		x"2b",	--2535
		x"3f",	--2536
		x"9f",	--2537
		x"2b",	--2538
		x"98",	--2539
		x"2f",	--2540
		x"3f",	--2541
		x"4a",	--2542
		x"4b",	--2543
		x"f0",	--2544
		x"00",	--2545
		x"f3",	--2546
		x"90",	--2547
		x"00",	--2548
		x"24",	--2549
		x"4a",	--2550
		x"00",	--2551
		x"4b",	--2552
		x"00",	--2553
		x"41",	--2554
		x"50",	--2555
		x"00",	--2556
		x"12",	--2557
		x"f6",	--2558
		x"50",	--2559
		x"00",	--2560
		x"41",	--2561
		x"41",	--2562
		x"41",	--2563
		x"41",	--2564
		x"41",	--2565
		x"41",	--2566
		x"42",	--2567
		x"00",	--2568
		x"41",	--2569
		x"50",	--2570
		x"00",	--2571
		x"3f",	--2572
		x"9e",	--2573
		x"23",	--2574
		x"40",	--2575
		x"fd",	--2576
		x"3f",	--2577
		x"93",	--2578
		x"23",	--2579
		x"4a",	--2580
		x"4b",	--2581
		x"f0",	--2582
		x"00",	--2583
		x"f3",	--2584
		x"93",	--2585
		x"23",	--2586
		x"93",	--2587
		x"23",	--2588
		x"93",	--2589
		x"20",	--2590
		x"93",	--2591
		x"27",	--2592
		x"50",	--2593
		x"00",	--2594
		x"63",	--2595
		x"f0",	--2596
		x"ff",	--2597
		x"f3",	--2598
		x"3f",	--2599
		x"43",	--2600
		x"00",	--2601
		x"43",	--2602
		x"00",	--2603
		x"43",	--2604
		x"00",	--2605
		x"41",	--2606
		x"50",	--2607
		x"00",	--2608
		x"3f",	--2609
		x"41",	--2610
		x"52",	--2611
		x"3f",	--2612
		x"50",	--2613
		x"ff",	--2614
		x"4e",	--2615
		x"00",	--2616
		x"4f",	--2617
		x"00",	--2618
		x"4c",	--2619
		x"00",	--2620
		x"4d",	--2621
		x"00",	--2622
		x"41",	--2623
		x"50",	--2624
		x"00",	--2625
		x"41",	--2626
		x"52",	--2627
		x"12",	--2628
		x"f8",	--2629
		x"41",	--2630
		x"52",	--2631
		x"41",	--2632
		x"12",	--2633
		x"f8",	--2634
		x"93",	--2635
		x"00",	--2636
		x"28",	--2637
		x"93",	--2638
		x"00",	--2639
		x"28",	--2640
		x"41",	--2641
		x"52",	--2642
		x"41",	--2643
		x"50",	--2644
		x"00",	--2645
		x"12",	--2646
		x"f9",	--2647
		x"50",	--2648
		x"00",	--2649
		x"41",	--2650
		x"43",	--2651
		x"3f",	--2652
		x"50",	--2653
		x"ff",	--2654
		x"4e",	--2655
		x"00",	--2656
		x"4f",	--2657
		x"00",	--2658
		x"41",	--2659
		x"52",	--2660
		x"41",	--2661
		x"12",	--2662
		x"f8",	--2663
		x"41",	--2664
		x"00",	--2665
		x"93",	--2666
		x"24",	--2667
		x"28",	--2668
		x"92",	--2669
		x"24",	--2670
		x"41",	--2671
		x"00",	--2672
		x"93",	--2673
		x"38",	--2674
		x"90",	--2675
		x"00",	--2676
		x"38",	--2677
		x"93",	--2678
		x"00",	--2679
		x"20",	--2680
		x"43",	--2681
		x"40",	--2682
		x"7f",	--2683
		x"50",	--2684
		x"00",	--2685
		x"41",	--2686
		x"41",	--2687
		x"00",	--2688
		x"41",	--2689
		x"00",	--2690
		x"40",	--2691
		x"00",	--2692
		x"8d",	--2693
		x"4c",	--2694
		x"f0",	--2695
		x"00",	--2696
		x"20",	--2697
		x"93",	--2698
		x"00",	--2699
		x"27",	--2700
		x"e3",	--2701
		x"e3",	--2702
		x"53",	--2703
		x"63",	--2704
		x"50",	--2705
		x"00",	--2706
		x"41",	--2707
		x"43",	--2708
		x"43",	--2709
		x"50",	--2710
		x"00",	--2711
		x"41",	--2712
		x"c3",	--2713
		x"10",	--2714
		x"10",	--2715
		x"53",	--2716
		x"23",	--2717
		x"3f",	--2718
		x"43",	--2719
		x"40",	--2720
		x"80",	--2721
		x"50",	--2722
		x"00",	--2723
		x"41",	--2724
		x"12",	--2725
		x"12",	--2726
		x"12",	--2727
		x"12",	--2728
		x"82",	--2729
		x"4e",	--2730
		x"4f",	--2731
		x"43",	--2732
		x"00",	--2733
		x"93",	--2734
		x"20",	--2735
		x"93",	--2736
		x"20",	--2737
		x"43",	--2738
		x"00",	--2739
		x"41",	--2740
		x"12",	--2741
		x"f6",	--2742
		x"52",	--2743
		x"41",	--2744
		x"41",	--2745
		x"41",	--2746
		x"41",	--2747
		x"41",	--2748
		x"40",	--2749
		x"00",	--2750
		x"00",	--2751
		x"40",	--2752
		x"00",	--2753
		x"00",	--2754
		x"4a",	--2755
		x"00",	--2756
		x"4b",	--2757
		x"00",	--2758
		x"4a",	--2759
		x"4b",	--2760
		x"12",	--2761
		x"f6",	--2762
		x"53",	--2763
		x"93",	--2764
		x"38",	--2765
		x"27",	--2766
		x"4a",	--2767
		x"00",	--2768
		x"4b",	--2769
		x"00",	--2770
		x"4f",	--2771
		x"f0",	--2772
		x"00",	--2773
		x"20",	--2774
		x"40",	--2775
		x"00",	--2776
		x"8f",	--2777
		x"4e",	--2778
		x"00",	--2779
		x"3f",	--2780
		x"51",	--2781
		x"00",	--2782
		x"00",	--2783
		x"61",	--2784
		x"00",	--2785
		x"00",	--2786
		x"53",	--2787
		x"23",	--2788
		x"3f",	--2789
		x"4f",	--2790
		x"e3",	--2791
		x"53",	--2792
		x"43",	--2793
		x"43",	--2794
		x"4e",	--2795
		x"f0",	--2796
		x"00",	--2797
		x"24",	--2798
		x"5c",	--2799
		x"6d",	--2800
		x"53",	--2801
		x"23",	--2802
		x"53",	--2803
		x"63",	--2804
		x"fa",	--2805
		x"fb",	--2806
		x"43",	--2807
		x"43",	--2808
		x"93",	--2809
		x"20",	--2810
		x"93",	--2811
		x"20",	--2812
		x"43",	--2813
		x"43",	--2814
		x"f0",	--2815
		x"00",	--2816
		x"20",	--2817
		x"48",	--2818
		x"49",	--2819
		x"da",	--2820
		x"db",	--2821
		x"4d",	--2822
		x"00",	--2823
		x"4e",	--2824
		x"00",	--2825
		x"40",	--2826
		x"00",	--2827
		x"8f",	--2828
		x"4e",	--2829
		x"00",	--2830
		x"3f",	--2831
		x"c3",	--2832
		x"10",	--2833
		x"10",	--2834
		x"53",	--2835
		x"23",	--2836
		x"3f",	--2837
		x"12",	--2838
		x"12",	--2839
		x"12",	--2840
		x"93",	--2841
		x"2c",	--2842
		x"90",	--2843
		x"01",	--2844
		x"28",	--2845
		x"40",	--2846
		x"00",	--2847
		x"43",	--2848
		x"42",	--2849
		x"4e",	--2850
		x"4f",	--2851
		x"49",	--2852
		x"93",	--2853
		x"20",	--2854
		x"50",	--2855
		x"fd",	--2856
		x"4c",	--2857
		x"43",	--2858
		x"8e",	--2859
		x"7f",	--2860
		x"4a",	--2861
		x"41",	--2862
		x"41",	--2863
		x"41",	--2864
		x"41",	--2865
		x"90",	--2866
		x"01",	--2867
		x"28",	--2868
		x"42",	--2869
		x"43",	--2870
		x"40",	--2871
		x"00",	--2872
		x"4e",	--2873
		x"4f",	--2874
		x"49",	--2875
		x"93",	--2876
		x"27",	--2877
		x"c3",	--2878
		x"10",	--2879
		x"10",	--2880
		x"53",	--2881
		x"23",	--2882
		x"3f",	--2883
		x"40",	--2884
		x"00",	--2885
		x"43",	--2886
		x"40",	--2887
		x"00",	--2888
		x"3f",	--2889
		x"40",	--2890
		x"00",	--2891
		x"43",	--2892
		x"43",	--2893
		x"3f",	--2894
		x"12",	--2895
		x"12",	--2896
		x"12",	--2897
		x"12",	--2898
		x"12",	--2899
		x"4f",	--2900
		x"4f",	--2901
		x"00",	--2902
		x"4f",	--2903
		x"00",	--2904
		x"4d",	--2905
		x"00",	--2906
		x"4d",	--2907
		x"93",	--2908
		x"28",	--2909
		x"92",	--2910
		x"24",	--2911
		x"93",	--2912
		x"24",	--2913
		x"93",	--2914
		x"24",	--2915
		x"4d",	--2916
		x"00",	--2917
		x"90",	--2918
		x"ff",	--2919
		x"38",	--2920
		x"90",	--2921
		x"00",	--2922
		x"34",	--2923
		x"4e",	--2924
		x"4f",	--2925
		x"f0",	--2926
		x"00",	--2927
		x"f3",	--2928
		x"90",	--2929
		x"00",	--2930
		x"24",	--2931
		x"50",	--2932
		x"00",	--2933
		x"63",	--2934
		x"93",	--2935
		x"38",	--2936
		x"4b",	--2937
		x"50",	--2938
		x"00",	--2939
		x"c3",	--2940
		x"10",	--2941
		x"10",	--2942
		x"c3",	--2943
		x"10",	--2944
		x"10",	--2945
		x"c3",	--2946
		x"10",	--2947
		x"10",	--2948
		x"c3",	--2949
		x"10",	--2950
		x"10",	--2951
		x"c3",	--2952
		x"10",	--2953
		x"10",	--2954
		x"c3",	--2955
		x"10",	--2956
		x"10",	--2957
		x"c3",	--2958
		x"10",	--2959
		x"10",	--2960
		x"f3",	--2961
		x"f0",	--2962
		x"00",	--2963
		x"4d",	--2964
		x"3c",	--2965
		x"93",	--2966
		x"23",	--2967
		x"43",	--2968
		x"43",	--2969
		x"43",	--2970
		x"4d",	--2971
		x"5d",	--2972
		x"5d",	--2973
		x"5d",	--2974
		x"5d",	--2975
		x"5d",	--2976
		x"5d",	--2977
		x"5d",	--2978
		x"4f",	--2979
		x"f0",	--2980
		x"00",	--2981
		x"dd",	--2982
		x"4a",	--2983
		x"11",	--2984
		x"43",	--2985
		x"10",	--2986
		x"4c",	--2987
		x"df",	--2988
		x"4d",	--2989
		x"41",	--2990
		x"41",	--2991
		x"41",	--2992
		x"41",	--2993
		x"41",	--2994
		x"41",	--2995
		x"93",	--2996
		x"23",	--2997
		x"4e",	--2998
		x"4f",	--2999
		x"f0",	--3000
		x"00",	--3001
		x"f3",	--3002
		x"93",	--3003
		x"20",	--3004
		x"93",	--3005
		x"27",	--3006
		x"50",	--3007
		x"00",	--3008
		x"63",	--3009
		x"3f",	--3010
		x"c3",	--3011
		x"10",	--3012
		x"10",	--3013
		x"4b",	--3014
		x"50",	--3015
		x"00",	--3016
		x"3f",	--3017
		x"43",	--3018
		x"43",	--3019
		x"43",	--3020
		x"3f",	--3021
		x"d3",	--3022
		x"d0",	--3023
		x"00",	--3024
		x"f3",	--3025
		x"f0",	--3026
		x"00",	--3027
		x"43",	--3028
		x"3f",	--3029
		x"40",	--3030
		x"ff",	--3031
		x"8b",	--3032
		x"90",	--3033
		x"00",	--3034
		x"34",	--3035
		x"4e",	--3036
		x"4f",	--3037
		x"47",	--3038
		x"f0",	--3039
		x"00",	--3040
		x"24",	--3041
		x"c3",	--3042
		x"10",	--3043
		x"10",	--3044
		x"53",	--3045
		x"23",	--3046
		x"43",	--3047
		x"43",	--3048
		x"f0",	--3049
		x"00",	--3050
		x"24",	--3051
		x"58",	--3052
		x"69",	--3053
		x"53",	--3054
		x"23",	--3055
		x"53",	--3056
		x"63",	--3057
		x"fe",	--3058
		x"ff",	--3059
		x"43",	--3060
		x"43",	--3061
		x"93",	--3062
		x"20",	--3063
		x"93",	--3064
		x"20",	--3065
		x"43",	--3066
		x"43",	--3067
		x"4e",	--3068
		x"4f",	--3069
		x"dc",	--3070
		x"dd",	--3071
		x"48",	--3072
		x"49",	--3073
		x"f0",	--3074
		x"00",	--3075
		x"f3",	--3076
		x"90",	--3077
		x"00",	--3078
		x"24",	--3079
		x"50",	--3080
		x"00",	--3081
		x"63",	--3082
		x"48",	--3083
		x"49",	--3084
		x"c3",	--3085
		x"10",	--3086
		x"10",	--3087
		x"c3",	--3088
		x"10",	--3089
		x"10",	--3090
		x"c3",	--3091
		x"10",	--3092
		x"10",	--3093
		x"c3",	--3094
		x"10",	--3095
		x"10",	--3096
		x"c3",	--3097
		x"10",	--3098
		x"10",	--3099
		x"c3",	--3100
		x"10",	--3101
		x"10",	--3102
		x"c3",	--3103
		x"10",	--3104
		x"10",	--3105
		x"f3",	--3106
		x"f0",	--3107
		x"00",	--3108
		x"43",	--3109
		x"90",	--3110
		x"40",	--3111
		x"2f",	--3112
		x"43",	--3113
		x"3f",	--3114
		x"43",	--3115
		x"43",	--3116
		x"3f",	--3117
		x"93",	--3118
		x"23",	--3119
		x"48",	--3120
		x"49",	--3121
		x"f0",	--3122
		x"00",	--3123
		x"f3",	--3124
		x"93",	--3125
		x"24",	--3126
		x"50",	--3127
		x"00",	--3128
		x"63",	--3129
		x"3f",	--3130
		x"93",	--3131
		x"27",	--3132
		x"3f",	--3133
		x"12",	--3134
		x"12",	--3135
		x"4f",	--3136
		x"4f",	--3137
		x"00",	--3138
		x"f0",	--3139
		x"00",	--3140
		x"4f",	--3141
		x"00",	--3142
		x"c3",	--3143
		x"10",	--3144
		x"c3",	--3145
		x"10",	--3146
		x"c3",	--3147
		x"10",	--3148
		x"c3",	--3149
		x"10",	--3150
		x"c3",	--3151
		x"10",	--3152
		x"c3",	--3153
		x"10",	--3154
		x"c3",	--3155
		x"10",	--3156
		x"4d",	--3157
		x"4f",	--3158
		x"00",	--3159
		x"b0",	--3160
		x"00",	--3161
		x"43",	--3162
		x"6f",	--3163
		x"4f",	--3164
		x"00",	--3165
		x"93",	--3166
		x"20",	--3167
		x"93",	--3168
		x"24",	--3169
		x"40",	--3170
		x"ff",	--3171
		x"00",	--3172
		x"4a",	--3173
		x"4b",	--3174
		x"5c",	--3175
		x"6d",	--3176
		x"5c",	--3177
		x"6d",	--3178
		x"5c",	--3179
		x"6d",	--3180
		x"5c",	--3181
		x"6d",	--3182
		x"5c",	--3183
		x"6d",	--3184
		x"5c",	--3185
		x"6d",	--3186
		x"5c",	--3187
		x"6d",	--3188
		x"40",	--3189
		x"00",	--3190
		x"00",	--3191
		x"90",	--3192
		x"40",	--3193
		x"2c",	--3194
		x"40",	--3195
		x"ff",	--3196
		x"5c",	--3197
		x"6d",	--3198
		x"4f",	--3199
		x"53",	--3200
		x"90",	--3201
		x"40",	--3202
		x"2b",	--3203
		x"4a",	--3204
		x"00",	--3205
		x"4c",	--3206
		x"00",	--3207
		x"4d",	--3208
		x"00",	--3209
		x"41",	--3210
		x"41",	--3211
		x"41",	--3212
		x"90",	--3213
		x"00",	--3214
		x"24",	--3215
		x"50",	--3216
		x"ff",	--3217
		x"4d",	--3218
		x"00",	--3219
		x"40",	--3220
		x"00",	--3221
		x"00",	--3222
		x"4a",	--3223
		x"4b",	--3224
		x"5c",	--3225
		x"6d",	--3226
		x"5c",	--3227
		x"6d",	--3228
		x"5c",	--3229
		x"6d",	--3230
		x"5c",	--3231
		x"6d",	--3232
		x"5c",	--3233
		x"6d",	--3234
		x"5c",	--3235
		x"6d",	--3236
		x"5c",	--3237
		x"6d",	--3238
		x"4c",	--3239
		x"4d",	--3240
		x"d3",	--3241
		x"d0",	--3242
		x"40",	--3243
		x"4a",	--3244
		x"00",	--3245
		x"4b",	--3246
		x"00",	--3247
		x"41",	--3248
		x"41",	--3249
		x"41",	--3250
		x"93",	--3251
		x"23",	--3252
		x"43",	--3253
		x"00",	--3254
		x"41",	--3255
		x"41",	--3256
		x"41",	--3257
		x"93",	--3258
		x"24",	--3259
		x"4a",	--3260
		x"4b",	--3261
		x"f3",	--3262
		x"f0",	--3263
		x"00",	--3264
		x"93",	--3265
		x"20",	--3266
		x"93",	--3267
		x"24",	--3268
		x"43",	--3269
		x"00",	--3270
		x"3f",	--3271
		x"93",	--3272
		x"23",	--3273
		x"42",	--3274
		x"00",	--3275
		x"3f",	--3276
		x"43",	--3277
		x"00",	--3278
		x"3f",	--3279
		x"12",	--3280
		x"4f",	--3281
		x"93",	--3282
		x"28",	--3283
		x"4e",	--3284
		x"93",	--3285
		x"28",	--3286
		x"92",	--3287
		x"24",	--3288
		x"92",	--3289
		x"24",	--3290
		x"93",	--3291
		x"24",	--3292
		x"93",	--3293
		x"24",	--3294
		x"4f",	--3295
		x"00",	--3296
		x"9e",	--3297
		x"00",	--3298
		x"24",	--3299
		x"93",	--3300
		x"20",	--3301
		x"43",	--3302
		x"4e",	--3303
		x"41",	--3304
		x"41",	--3305
		x"93",	--3306
		x"24",	--3307
		x"93",	--3308
		x"00",	--3309
		x"23",	--3310
		x"43",	--3311
		x"4e",	--3312
		x"41",	--3313
		x"41",	--3314
		x"93",	--3315
		x"00",	--3316
		x"27",	--3317
		x"43",	--3318
		x"3f",	--3319
		x"4f",	--3320
		x"00",	--3321
		x"4e",	--3322
		x"00",	--3323
		x"9b",	--3324
		x"3b",	--3325
		x"9c",	--3326
		x"38",	--3327
		x"4f",	--3328
		x"00",	--3329
		x"4f",	--3330
		x"00",	--3331
		x"4e",	--3332
		x"00",	--3333
		x"4e",	--3334
		x"00",	--3335
		x"9f",	--3336
		x"2b",	--3337
		x"9e",	--3338
		x"28",	--3339
		x"9b",	--3340
		x"2b",	--3341
		x"9e",	--3342
		x"28",	--3343
		x"9f",	--3344
		x"28",	--3345
		x"9c",	--3346
		x"28",	--3347
		x"43",	--3348
		x"3f",	--3349
		x"93",	--3350
		x"23",	--3351
		x"43",	--3352
		x"3f",	--3353
		x"92",	--3354
		x"23",	--3355
		x"4e",	--3356
		x"00",	--3357
		x"4f",	--3358
		x"00",	--3359
		x"8f",	--3360
		x"3f",	--3361
		x"43",	--3362
		x"93",	--3363
		x"34",	--3364
		x"40",	--3365
		x"00",	--3366
		x"e3",	--3367
		x"53",	--3368
		x"93",	--3369
		x"34",	--3370
		x"e3",	--3371
		x"e3",	--3372
		x"53",	--3373
		x"12",	--3374
		x"12",	--3375
		x"fb",	--3376
		x"41",	--3377
		x"b3",	--3378
		x"24",	--3379
		x"e3",	--3380
		x"53",	--3381
		x"b3",	--3382
		x"24",	--3383
		x"e3",	--3384
		x"53",	--3385
		x"41",	--3386
		x"12",	--3387
		x"fa",	--3388
		x"4e",	--3389
		x"41",	--3390
		x"12",	--3391
		x"12",	--3392
		x"12",	--3393
		x"40",	--3394
		x"00",	--3395
		x"4c",	--3396
		x"4d",	--3397
		x"43",	--3398
		x"43",	--3399
		x"5e",	--3400
		x"6f",	--3401
		x"6c",	--3402
		x"6d",	--3403
		x"9b",	--3404
		x"28",	--3405
		x"20",	--3406
		x"9a",	--3407
		x"28",	--3408
		x"8a",	--3409
		x"7b",	--3410
		x"d3",	--3411
		x"83",	--3412
		x"23",	--3413
		x"41",	--3414
		x"41",	--3415
		x"41",	--3416
		x"41",	--3417
		x"12",	--3418
		x"fa",	--3419
		x"4c",	--3420
		x"4d",	--3421
		x"41",	--3422
		x"12",	--3423
		x"43",	--3424
		x"93",	--3425
		x"34",	--3426
		x"40",	--3427
		x"00",	--3428
		x"e3",	--3429
		x"e3",	--3430
		x"53",	--3431
		x"63",	--3432
		x"93",	--3433
		x"34",	--3434
		x"e3",	--3435
		x"e3",	--3436
		x"e3",	--3437
		x"53",	--3438
		x"63",	--3439
		x"12",	--3440
		x"fa",	--3441
		x"b3",	--3442
		x"24",	--3443
		x"e3",	--3444
		x"e3",	--3445
		x"53",	--3446
		x"63",	--3447
		x"b3",	--3448
		x"24",	--3449
		x"e3",	--3450
		x"e3",	--3451
		x"53",	--3452
		x"63",	--3453
		x"41",	--3454
		x"41",	--3455
		x"12",	--3456
		x"fa",	--3457
		x"4c",	--3458
		x"4d",	--3459
		x"41",	--3460
		x"40",	--3461
		x"00",	--3462
		x"4e",	--3463
		x"43",	--3464
		x"5f",	--3465
		x"6e",	--3466
		x"9d",	--3467
		x"28",	--3468
		x"8d",	--3469
		x"d3",	--3470
		x"83",	--3471
		x"23",	--3472
		x"41",	--3473
		x"12",	--3474
		x"fb",	--3475
		x"4e",	--3476
		x"41",	--3477
		x"13",	--3478
		x"d0",	--3479
		x"00",	--3480
		x"3f",	--3481
		x"61",	--3482
		x"74",	--3483
		x"6e",	--3484
		x"20",	--3485
		x"6f",	--3486
		x"20",	--3487
		x"20",	--3488
		x"65",	--3489
		x"20",	--3490
		x"62",	--3491
		x"6e",	--3492
		x"66",	--3493
		x"6c",	--3494
		x"0d",	--3495
		x"00",	--3496
		x"65",	--3497
		x"73",	--3498
		x"6f",	--3499
		x"6c",	--3500
		x"20",	--3501
		x"6f",	--3502
		x"20",	--3503
		x"65",	--3504
		x"20",	--3505
		x"68",	--3506
		x"74",	--3507
		x"0a",	--3508
		x"53",	--3509
		x"6f",	--3510
		x"0d",	--3511
		x"00",	--3512
		x"72",	--3513
		x"6f",	--3514
		x"3a",	--3515
		x"6d",	--3516
		x"73",	--3517
		x"69",	--3518
		x"67",	--3519
		x"61",	--3520
		x"67",	--3521
		x"6d",	--3522
		x"6e",	--3523
		x"0d",	--3524
		x"00",	--3525
		x"6f",	--3526
		x"72",	--3527
		x"63",	--3528
		x"20",	--3529
		x"73",	--3530
		x"67",	--3531
		x"3a",	--3532
		x"0a",	--3533
		x"09",	--3534
		x"73",	--3535
		x"4c",	--3536
		x"46",	--3537
		x"20",	--3538
		x"49",	--3539
		x"48",	--3540
		x"20",	--3541
		x"54",	--3542
		x"4d",	--3543
		x"4f",	--3544
		x"54",	--3545
		x"0d",	--3546
		x"00",	--3547
		x"64",	--3548
		x"25",	--3549
		x"0d",	--3550
		x"00",	--3551
		x"77",	--3552
		x"25",	--3553
		x"20",	--3554
		x"77",	--3555
		x"25",	--3556
		x"0d",	--3557
		x"00",	--3558
		x"e4",	--3559
		x"e4",	--3560
		x"e4",	--3561
		x"e4",	--3562
		x"e4",	--3563
		x"e4",	--3564
		x"e4",	--3565
		x"e4",	--3566
		x"0a",	--3567
		x"3d",	--3568
		x"3d",	--3569
		x"3d",	--3570
		x"4d",	--3571
		x"72",	--3572
		x"65",	--3573
		x"20",	--3574
		x"43",	--3575
		x"20",	--3576
		x"3d",	--3577
		x"3d",	--3578
		x"3d",	--3579
		x"0a",	--3580
		x"69",	--3581
		x"74",	--3582
		x"72",	--3583
		x"63",	--3584
		x"69",	--3585
		x"65",	--3586
		x"6d",	--3587
		x"64",	--3588
		x"00",	--3589
		x"72",	--3590
		x"74",	--3591
		x"00",	--3592
		x"65",	--3593
		x"64",	--3594
		x"70",	--3595
		x"6d",	--3596
		x"65",	--3597
		x"63",	--3598
		x"64",	--3599
		x"72",	--3600
		x"62",	--3601
		x"6f",	--3602
		x"6c",	--3603
		x"61",	--3604
		x"65",	--3605
		x"00",	--3606
		x"0a",	--3607
		x"08",	--3608
		x"08",	--3609
		x"25",	--3610
		x"00",	--3611
		x"72",	--3612
		x"74",	--3613
		x"0a",	--3614
		x"00",	--3615
		x"72",	--3616
		x"6f",	--3617
		x"3a",	--3618
		x"6d",	--3619
		x"73",	--3620
		x"69",	--3621
		x"67",	--3622
		x"61",	--3623
		x"67",	--3624
		x"6d",	--3625
		x"6e",	--3626
		x"0d",	--3627
		x"00",	--3628
		x"6f",	--3629
		x"72",	--3630
		x"63",	--3631
		x"20",	--3632
		x"73",	--3633
		x"67",	--3634
		x"3a",	--3635
		x"0a",	--3636
		x"09",	--3637
		x"73",	--3638
		x"52",	--3639
		x"47",	--3640
		x"53",	--3641
		x"45",	--3642
		x"20",	--3643
		x"41",	--3644
		x"55",	--3645
		x"0d",	--3646
		x"00",	--3647
		x"3d",	--3648
		x"64",	--3649
		x"76",	--3650
		x"25",	--3651
		x"0d",	--3652
		x"00",	--3653
		x"25",	--3654
		x"20",	--3655
		x"45",	--3656
		x"49",	--3657
		x"54",	--3658
		x"52",	--3659
		x"0a",	--3660
		x"72",	--3661
		x"61",	--3662
		x"0a",	--3663
		x"00",	--3664
		x"63",	--3665
		x"69",	--3666
		x"20",	--3667
		x"6f",	--3668
		x"20",	--3669
		x"20",	--3670
		x"75",	--3671
		x"62",	--3672
		x"72",	--3673
		x"0a",	--3674
		x"25",	--3675
		x"20",	--3676
		x"73",	--3677
		x"0a",	--3678
		x"25",	--3679
		x"3a",	--3680
		x"6e",	--3681
		x"20",	--3682
		x"75",	--3683
		x"68",	--3684
		x"63",	--3685
		x"6d",	--3686
		x"61",	--3687
		x"64",	--3688
		x"0a",	--3689
		x"00",	--3690
		x"ec",	--3691
		x"eb",	--3692
		x"eb",	--3693
		x"eb",	--3694
		x"eb",	--3695
		x"eb",	--3696
		x"eb",	--3697
		x"eb",	--3698
		x"eb",	--3699
		x"eb",	--3700
		x"eb",	--3701
		x"eb",	--3702
		x"eb",	--3703
		x"eb",	--3704
		x"eb",	--3705
		x"eb",	--3706
		x"eb",	--3707
		x"eb",	--3708
		x"eb",	--3709
		x"eb",	--3710
		x"eb",	--3711
		x"eb",	--3712
		x"eb",	--3713
		x"eb",	--3714
		x"eb",	--3715
		x"eb",	--3716
		x"eb",	--3717
		x"eb",	--3718
		x"eb",	--3719
		x"ec",	--3720
		x"eb",	--3721
		x"eb",	--3722
		x"eb",	--3723
		x"eb",	--3724
		x"eb",	--3725
		x"eb",	--3726
		x"eb",	--3727
		x"eb",	--3728
		x"eb",	--3729
		x"eb",	--3730
		x"eb",	--3731
		x"eb",	--3732
		x"eb",	--3733
		x"eb",	--3734
		x"eb",	--3735
		x"eb",	--3736
		x"eb",	--3737
		x"eb",	--3738
		x"eb",	--3739
		x"eb",	--3740
		x"eb",	--3741
		x"eb",	--3742
		x"eb",	--3743
		x"eb",	--3744
		x"eb",	--3745
		x"eb",	--3746
		x"eb",	--3747
		x"eb",	--3748
		x"eb",	--3749
		x"eb",	--3750
		x"eb",	--3751
		x"ec",	--3752
		x"ec",	--3753
		x"ec",	--3754
		x"eb",	--3755
		x"eb",	--3756
		x"eb",	--3757
		x"eb",	--3758
		x"eb",	--3759
		x"eb",	--3760
		x"eb",	--3761
		x"ec",	--3762
		x"eb",	--3763
		x"ec",	--3764
		x"eb",	--3765
		x"eb",	--3766
		x"eb",	--3767
		x"eb",	--3768
		x"ec",	--3769
		x"eb",	--3770
		x"eb",	--3771
		x"eb",	--3772
		x"ec",	--3773
		x"ec",	--3774
		x"31",	--3775
		x"33",	--3776
		x"35",	--3777
		x"37",	--3778
		x"39",	--3779
		x"62",	--3780
		x"64",	--3781
		x"66",	--3782
		x"00",	--3783
		x"00",	--3784
		x"00",	--3785
		x"00",	--3786
		x"00",	--3787
		x"01",	--3788
		x"02",	--3789
		x"03",	--3790
		x"03",	--3791
		x"04",	--3792
		x"04",	--3793
		x"04",	--3794
		x"04",	--3795
		x"05",	--3796
		x"05",	--3797
		x"05",	--3798
		x"05",	--3799
		x"05",	--3800
		x"05",	--3801
		x"05",	--3802
		x"05",	--3803
		x"06",	--3804
		x"06",	--3805
		x"06",	--3806
		x"06",	--3807
		x"06",	--3808
		x"06",	--3809
		x"06",	--3810
		x"06",	--3811
		x"06",	--3812
		x"06",	--3813
		x"06",	--3814
		x"06",	--3815
		x"06",	--3816
		x"06",	--3817
		x"06",	--3818
		x"06",	--3819
		x"07",	--3820
		x"07",	--3821
		x"07",	--3822
		x"07",	--3823
		x"07",	--3824
		x"07",	--3825
		x"07",	--3826
		x"07",	--3827
		x"07",	--3828
		x"07",	--3829
		x"07",	--3830
		x"07",	--3831
		x"07",	--3832
		x"07",	--3833
		x"07",	--3834
		x"07",	--3835
		x"07",	--3836
		x"07",	--3837
		x"07",	--3838
		x"07",	--3839
		x"07",	--3840
		x"07",	--3841
		x"07",	--3842
		x"07",	--3843
		x"07",	--3844
		x"07",	--3845
		x"07",	--3846
		x"07",	--3847
		x"07",	--3848
		x"07",	--3849
		x"07",	--3850
		x"07",	--3851
		x"08",	--3852
		x"08",	--3853
		x"08",	--3854
		x"08",	--3855
		x"08",	--3856
		x"08",	--3857
		x"08",	--3858
		x"08",	--3859
		x"08",	--3860
		x"08",	--3861
		x"08",	--3862
		x"08",	--3863
		x"08",	--3864
		x"08",	--3865
		x"08",	--3866
		x"08",	--3867
		x"08",	--3868
		x"08",	--3869
		x"08",	--3870
		x"08",	--3871
		x"08",	--3872
		x"08",	--3873
		x"08",	--3874
		x"08",	--3875
		x"08",	--3876
		x"08",	--3877
		x"08",	--3878
		x"08",	--3879
		x"08",	--3880
		x"08",	--3881
		x"08",	--3882
		x"08",	--3883
		x"08",	--3884
		x"08",	--3885
		x"08",	--3886
		x"08",	--3887
		x"08",	--3888
		x"08",	--3889
		x"08",	--3890
		x"08",	--3891
		x"08",	--3892
		x"08",	--3893
		x"08",	--3894
		x"08",	--3895
		x"08",	--3896
		x"08",	--3897
		x"08",	--3898
		x"08",	--3899
		x"08",	--3900
		x"08",	--3901
		x"08",	--3902
		x"08",	--3903
		x"08",	--3904
		x"08",	--3905
		x"08",	--3906
		x"08",	--3907
		x"08",	--3908
		x"08",	--3909
		x"08",	--3910
		x"08",	--3911
		x"08",	--3912
		x"08",	--3913
		x"08",	--3914
		x"08",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"65",	--3918
		x"70",	--3919
		x"00",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"ec",	--4087
		x"e9",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
