library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"58",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"06",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"58",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"90",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"52",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"58",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"06",	--29
		x"f9",	--30
		x"31",	--31
		x"be",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"80",	--41
		x"0f",	--42
		x"b0",	--43
		x"4e",	--44
		x"b0",	--45
		x"94",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"e1",	--50
		x"b0",	--51
		x"12",	--52
		x"21",	--53
		x"3d",	--54
		x"fe",	--55
		x"3e",	--56
		x"32",	--57
		x"7f",	--58
		x"77",	--59
		x"b0",	--60
		x"c4",	--61
		x"3d",	--62
		x"04",	--63
		x"3e",	--64
		x"d2",	--65
		x"7f",	--66
		x"72",	--67
		x"b0",	--68
		x"c4",	--69
		x"3d",	--70
		x"09",	--71
		x"3e",	--72
		x"f4",	--73
		x"7f",	--74
		x"70",	--75
		x"b0",	--76
		x"c4",	--77
		x"3d",	--78
		x"0d",	--79
		x"3e",	--80
		x"b0",	--81
		x"7f",	--82
		x"65",	--83
		x"b0",	--84
		x"c4",	--85
		x"3d",	--86
		x"15",	--87
		x"3e",	--88
		x"be",	--89
		x"7f",	--90
		x"62",	--91
		x"b0",	--92
		x"c4",	--93
		x"0f",	--94
		x"b0",	--95
		x"5a",	--96
		x"2c",	--97
		x"3d",	--98
		x"20",	--99
		x"3e",	--100
		x"80",	--101
		x"0f",	--102
		x"3f",	--103
		x"0e",	--104
		x"b0",	--105
		x"6a",	--106
		x"0f",	--107
		x"3f",	--108
		x"0e",	--109
		x"b0",	--110
		x"b2",	--111
		x"2c",	--112
		x"3d",	--113
		x"20",	--114
		x"3e",	--115
		x"88",	--116
		x"0f",	--117
		x"2f",	--118
		x"b0",	--119
		x"6a",	--120
		x"0f",	--121
		x"2f",	--122
		x"b0",	--123
		x"b2",	--124
		x"0e",	--125
		x"2e",	--126
		x"0f",	--127
		x"3f",	--128
		x"0e",	--129
		x"b0",	--130
		x"ea",	--131
		x"3e",	--132
		x"98",	--133
		x"0f",	--134
		x"2f",	--135
		x"b0",	--136
		x"28",	--137
		x"3e",	--138
		x"9a",	--139
		x"0f",	--140
		x"b0",	--141
		x"28",	--142
		x"0e",	--143
		x"0f",	--144
		x"2f",	--145
		x"b0",	--146
		x"a6",	--147
		x"b0",	--148
		x"48",	--149
		x"0d",	--150
		x"3e",	--151
		x"c8",	--152
		x"3f",	--153
		x"f4",	--154
		x"b0",	--155
		x"58",	--156
		x"b0",	--157
		x"9e",	--158
		x"f2",	--159
		x"80",	--160
		x"19",	--161
		x"32",	--162
		x"0b",	--163
		x"b0",	--164
		x"5c",	--165
		x"0f",	--166
		x"fc",	--167
		x"b0",	--168
		x"84",	--169
		x"7f",	--170
		x"11",	--171
		x"7f",	--172
		x"0d",	--173
		x"17",	--174
		x"30",	--175
		x"20",	--176
		x"b0",	--177
		x"12",	--178
		x"21",	--179
		x"0e",	--180
		x"3e",	--181
		x"18",	--182
		x"5f",	--183
		x"18",	--184
		x"b0",	--185
		x"f8",	--186
		x"0b",	--187
		x"e7",	--188
		x"0b",	--189
		x"e5",	--190
		x"3b",	--191
		x"30",	--192
		x"23",	--193
		x"b0",	--194
		x"12",	--195
		x"21",	--196
		x"de",	--197
		x"3b",	--198
		x"28",	--199
		x"db",	--200
		x"4e",	--201
		x"8e",	--202
		x"0e",	--203
		x"30",	--204
		x"27",	--205
		x"81",	--206
		x"44",	--207
		x"b0",	--208
		x"12",	--209
		x"21",	--210
		x"3e",	--211
		x"18",	--212
		x"0e",	--213
		x"0e",	--214
		x"1f",	--215
		x"40",	--216
		x"ce",	--217
		x"00",	--218
		x"1b",	--219
		x"c7",	--220
		x"30",	--221
		x"58",	--222
		x"b2",	--223
		x"00",	--224
		x"92",	--225
		x"a2",	--226
		x"94",	--227
		x"b2",	--228
		x"6d",	--229
		x"96",	--230
		x"30",	--231
		x"60",	--232
		x"b0",	--233
		x"12",	--234
		x"92",	--235
		x"90",	--236
		x"b1",	--237
		x"7e",	--238
		x"00",	--239
		x"b0",	--240
		x"12",	--241
		x"21",	--242
		x"0f",	--243
		x"30",	--244
		x"82",	--245
		x"12",	--246
		x"82",	--247
		x"10",	--248
		x"30",	--249
		x"31",	--250
		x"ff",	--251
		x"20",	--252
		x"01",	--253
		x"39",	--254
		x"cf",	--255
		x"02",	--256
		x"36",	--257
		x"0d",	--258
		x"0e",	--259
		x"2e",	--260
		x"0f",	--261
		x"2f",	--262
		x"b0",	--263
		x"50",	--264
		x"81",	--265
		x"00",	--266
		x"40",	--267
		x"0d",	--268
		x"0e",	--269
		x"0f",	--270
		x"2f",	--271
		x"b0",	--272
		x"50",	--273
		x"81",	--274
		x"00",	--275
		x"37",	--276
		x"1e",	--277
		x"04",	--278
		x"0f",	--279
		x"b0",	--280
		x"76",	--281
		x"0c",	--282
		x"3d",	--283
		x"c8",	--284
		x"b0",	--285
		x"46",	--286
		x"0d",	--287
		x"0e",	--288
		x"1f",	--289
		x"12",	--290
		x"b0",	--291
		x"06",	--292
		x"1e",	--293
		x"02",	--294
		x"0f",	--295
		x"b0",	--296
		x"76",	--297
		x"0c",	--298
		x"3d",	--299
		x"c8",	--300
		x"b0",	--301
		x"46",	--302
		x"0d",	--303
		x"0e",	--304
		x"1f",	--305
		x"10",	--306
		x"b0",	--307
		x"06",	--308
		x"0f",	--309
		x"31",	--310
		x"30",	--311
		x"30",	--312
		x"97",	--313
		x"81",	--314
		x"08",	--315
		x"b0",	--316
		x"12",	--317
		x"1f",	--318
		x"08",	--319
		x"6f",	--320
		x"8f",	--321
		x"81",	--322
		x"00",	--323
		x"30",	--324
		x"a8",	--325
		x"b0",	--326
		x"12",	--327
		x"21",	--328
		x"3f",	--329
		x"31",	--330
		x"30",	--331
		x"30",	--332
		x"b9",	--333
		x"b0",	--334
		x"12",	--335
		x"21",	--336
		x"3f",	--337
		x"e3",	--338
		x"82",	--339
		x"14",	--340
		x"82",	--341
		x"16",	--342
		x"30",	--343
		x"12",	--344
		x"9a",	--345
		x"12",	--346
		x"98",	--347
		x"30",	--348
		x"d9",	--349
		x"b0",	--350
		x"12",	--351
		x"31",	--352
		x"06",	--353
		x"0f",	--354
		x"30",	--355
		x"1f",	--356
		x"06",	--357
		x"1f",	--358
		x"18",	--359
		x"2f",	--360
		x"1c",	--361
		x"09",	--362
		x"3f",	--363
		x"03",	--364
		x"0d",	--365
		x"3f",	--366
		x"03",	--367
		x"06",	--368
		x"82",	--369
		x"06",	--370
		x"30",	--371
		x"f2",	--372
		x"0c",	--373
		x"19",	--374
		x"1f",	--375
		x"82",	--376
		x"06",	--377
		x"30",	--378
		x"f2",	--379
		x"19",	--380
		x"82",	--381
		x"06",	--382
		x"30",	--383
		x"e2",	--384
		x"19",	--385
		x"1f",	--386
		x"82",	--387
		x"06",	--388
		x"30",	--389
		x"0f",	--390
		x"e6",	--391
		x"c2",	--392
		x"19",	--393
		x"1f",	--394
		x"82",	--395
		x"06",	--396
		x"30",	--397
		x"5e",	--398
		x"19",	--399
		x"4e",	--400
		x"0f",	--401
		x"03",	--402
		x"c2",	--403
		x"19",	--404
		x"30",	--405
		x"c2",	--406
		x"19",	--407
		x"30",	--408
		x"0b",	--409
		x"31",	--410
		x"fa",	--411
		x"0b",	--412
		x"30",	--413
		x"2a",	--414
		x"b0",	--415
		x"12",	--416
		x"21",	--417
		x"fb",	--418
		x"20",	--419
		x"01",	--420
		x"2a",	--421
		x"cb",	--422
		x"02",	--423
		x"27",	--424
		x"0d",	--425
		x"0e",	--426
		x"2e",	--427
		x"0f",	--428
		x"2f",	--429
		x"b0",	--430
		x"50",	--431
		x"81",	--432
		x"00",	--433
		x"2f",	--434
		x"0d",	--435
		x"0e",	--436
		x"0f",	--437
		x"2f",	--438
		x"b0",	--439
		x"50",	--440
		x"81",	--441
		x"00",	--442
		x"26",	--443
		x"11",	--444
		x"04",	--445
		x"11",	--446
		x"08",	--447
		x"30",	--448
		x"78",	--449
		x"b0",	--450
		x"12",	--451
		x"31",	--452
		x"06",	--453
		x"1f",	--454
		x"04",	--455
		x"9f",	--456
		x"02",	--457
		x"00",	--458
		x"0f",	--459
		x"31",	--460
		x"06",	--461
		x"3b",	--462
		x"30",	--463
		x"30",	--464
		x"32",	--465
		x"b0",	--466
		x"12",	--467
		x"6f",	--468
		x"8f",	--469
		x"81",	--470
		x"00",	--471
		x"30",	--472
		x"43",	--473
		x"b0",	--474
		x"12",	--475
		x"21",	--476
		x"3f",	--477
		x"31",	--478
		x"06",	--479
		x"3b",	--480
		x"30",	--481
		x"30",	--482
		x"58",	--483
		x"b0",	--484
		x"12",	--485
		x"21",	--486
		x"3f",	--487
		x"e3",	--488
		x"0b",	--489
		x"21",	--490
		x"0b",	--491
		x"30",	--492
		x"84",	--493
		x"b0",	--494
		x"12",	--495
		x"21",	--496
		x"fb",	--497
		x"20",	--498
		x"01",	--499
		x"1b",	--500
		x"cb",	--501
		x"02",	--502
		x"18",	--503
		x"0d",	--504
		x"0e",	--505
		x"2e",	--506
		x"0f",	--507
		x"2f",	--508
		x"b0",	--509
		x"50",	--510
		x"81",	--511
		x"00",	--512
		x"1f",	--513
		x"1f",	--514
		x"02",	--515
		x"2f",	--516
		x"0f",	--517
		x"30",	--518
		x"78",	--519
		x"b0",	--520
		x"12",	--521
		x"31",	--522
		x"06",	--523
		x"0f",	--524
		x"21",	--525
		x"3b",	--526
		x"30",	--527
		x"30",	--528
		x"32",	--529
		x"b0",	--530
		x"12",	--531
		x"6f",	--532
		x"8f",	--533
		x"81",	--534
		x"00",	--535
		x"30",	--536
		x"8b",	--537
		x"b0",	--538
		x"12",	--539
		x"21",	--540
		x"3f",	--541
		x"21",	--542
		x"3b",	--543
		x"30",	--544
		x"30",	--545
		x"58",	--546
		x"b0",	--547
		x"12",	--548
		x"21",	--549
		x"3f",	--550
		x"e5",	--551
		x"0b",	--552
		x"0a",	--553
		x"09",	--554
		x"08",	--555
		x"07",	--556
		x"8f",	--557
		x"00",	--558
		x"8d",	--559
		x"00",	--560
		x"6c",	--561
		x"4c",	--562
		x"5f",	--563
		x"0b",	--564
		x"1b",	--565
		x"08",	--566
		x"0a",	--567
		x"07",	--568
		x"09",	--569
		x"18",	--570
		x"7a",	--571
		x"0a",	--572
		x"35",	--573
		x"2c",	--574
		x"0c",	--575
		x"0c",	--576
		x"0c",	--577
		x"0c",	--578
		x"8f",	--579
		x"00",	--580
		x"3c",	--581
		x"d0",	--582
		x"6a",	--583
		x"8a",	--584
		x"0c",	--585
		x"8f",	--586
		x"00",	--587
		x"17",	--588
		x"19",	--589
		x"0a",	--590
		x"08",	--591
		x"7c",	--592
		x"4c",	--593
		x"40",	--594
		x"7c",	--595
		x"78",	--596
		x"1b",	--597
		x"7c",	--598
		x"20",	--599
		x"43",	--600
		x"4a",	--601
		x"7a",	--602
		x"d0",	--603
		x"07",	--604
		x"dd",	--605
		x"7a",	--606
		x"0a",	--607
		x"46",	--608
		x"2a",	--609
		x"0a",	--610
		x"0c",	--611
		x"0c",	--612
		x"0c",	--613
		x"0c",	--614
		x"8f",	--615
		x"00",	--616
		x"3c",	--617
		x"d0",	--618
		x"68",	--619
		x"88",	--620
		x"0c",	--621
		x"8f",	--622
		x"00",	--623
		x"dc",	--624
		x"17",	--625
		x"da",	--626
		x"4a",	--627
		x"7a",	--628
		x"9f",	--629
		x"7a",	--630
		x"06",	--631
		x"0a",	--632
		x"2c",	--633
		x"0c",	--634
		x"0c",	--635
		x"0c",	--636
		x"0c",	--637
		x"8f",	--638
		x"00",	--639
		x"3c",	--640
		x"a9",	--641
		x"c4",	--642
		x"4a",	--643
		x"7a",	--644
		x"bf",	--645
		x"7a",	--646
		x"06",	--647
		x"1e",	--648
		x"2c",	--649
		x"0c",	--650
		x"0c",	--651
		x"0c",	--652
		x"0c",	--653
		x"8f",	--654
		x"00",	--655
		x"3c",	--656
		x"c9",	--657
		x"b4",	--658
		x"9d",	--659
		x"00",	--660
		x"0f",	--661
		x"37",	--662
		x"38",	--663
		x"39",	--664
		x"3a",	--665
		x"3b",	--666
		x"30",	--667
		x"9d",	--668
		x"00",	--669
		x"0f",	--670
		x"1f",	--671
		x"0f",	--672
		x"37",	--673
		x"38",	--674
		x"39",	--675
		x"3a",	--676
		x"3b",	--677
		x"30",	--678
		x"8c",	--679
		x"0c",	--680
		x"30",	--681
		x"9a",	--682
		x"b0",	--683
		x"12",	--684
		x"21",	--685
		x"0f",	--686
		x"37",	--687
		x"38",	--688
		x"39",	--689
		x"3a",	--690
		x"3b",	--691
		x"30",	--692
		x"0b",	--693
		x"0a",	--694
		x"0b",	--695
		x"0a",	--696
		x"8f",	--697
		x"00",	--698
		x"8f",	--699
		x"02",	--700
		x"8f",	--701
		x"04",	--702
		x"0c",	--703
		x"0d",	--704
		x"3e",	--705
		x"00",	--706
		x"3f",	--707
		x"6e",	--708
		x"b0",	--709
		x"aa",	--710
		x"8b",	--711
		x"02",	--712
		x"02",	--713
		x"32",	--714
		x"03",	--715
		x"82",	--716
		x"32",	--717
		x"b2",	--718
		x"18",	--719
		x"38",	--720
		x"9b",	--721
		x"3a",	--722
		x"06",	--723
		x"32",	--724
		x"0f",	--725
		x"3a",	--726
		x"3b",	--727
		x"30",	--728
		x"0b",	--729
		x"09",	--730
		x"08",	--731
		x"8f",	--732
		x"06",	--733
		x"bf",	--734
		x"00",	--735
		x"08",	--736
		x"2b",	--737
		x"1e",	--738
		x"02",	--739
		x"0f",	--740
		x"b0",	--741
		x"76",	--742
		x"0c",	--743
		x"3d",	--744
		x"00",	--745
		x"b0",	--746
		x"22",	--747
		x"08",	--748
		x"09",	--749
		x"1e",	--750
		x"06",	--751
		x"0f",	--752
		x"b0",	--753
		x"76",	--754
		x"0c",	--755
		x"0d",	--756
		x"0e",	--757
		x"0f",	--758
		x"b0",	--759
		x"d2",	--760
		x"b0",	--761
		x"b2",	--762
		x"8b",	--763
		x"04",	--764
		x"9b",	--765
		x"00",	--766
		x"38",	--767
		x"39",	--768
		x"3b",	--769
		x"30",	--770
		x"0b",	--771
		x"0a",	--772
		x"09",	--773
		x"0a",	--774
		x"0b",	--775
		x"8f",	--776
		x"06",	--777
		x"8f",	--778
		x"08",	--779
		x"29",	--780
		x"1e",	--781
		x"02",	--782
		x"0f",	--783
		x"b0",	--784
		x"76",	--785
		x"0c",	--786
		x"0d",	--787
		x"0e",	--788
		x"0f",	--789
		x"b0",	--790
		x"22",	--791
		x"0a",	--792
		x"0b",	--793
		x"1e",	--794
		x"06",	--795
		x"0f",	--796
		x"b0",	--797
		x"76",	--798
		x"0c",	--799
		x"0d",	--800
		x"0e",	--801
		x"0f",	--802
		x"b0",	--803
		x"d2",	--804
		x"b0",	--805
		x"b2",	--806
		x"89",	--807
		x"04",	--808
		x"39",	--809
		x"3a",	--810
		x"3b",	--811
		x"30",	--812
		x"0b",	--813
		x"0a",	--814
		x"92",	--815
		x"08",	--816
		x"14",	--817
		x"3b",	--818
		x"1c",	--819
		x"0a",	--820
		x"2b",	--821
		x"5f",	--822
		x"fc",	--823
		x"8f",	--824
		x"0f",	--825
		x"30",	--826
		x"af",	--827
		x"b0",	--828
		x"12",	--829
		x"31",	--830
		x"06",	--831
		x"1a",	--832
		x"3b",	--833
		x"06",	--834
		x"1a",	--835
		x"08",	--836
		x"ef",	--837
		x"0f",	--838
		x"3a",	--839
		x"3b",	--840
		x"30",	--841
		x"1e",	--842
		x"08",	--843
		x"3e",	--844
		x"20",	--845
		x"12",	--846
		x"0f",	--847
		x"0f",	--848
		x"0f",	--849
		x"0f",	--850
		x"3f",	--851
		x"18",	--852
		x"ff",	--853
		x"68",	--854
		x"00",	--855
		x"bf",	--856
		x"5a",	--857
		x"02",	--858
		x"bf",	--859
		x"00",	--860
		x"04",	--861
		x"1e",	--862
		x"82",	--863
		x"08",	--864
		x"30",	--865
		x"0b",	--866
		x"1b",	--867
		x"08",	--868
		x"3b",	--869
		x"20",	--870
		x"12",	--871
		x"0c",	--872
		x"0c",	--873
		x"0c",	--874
		x"0c",	--875
		x"3c",	--876
		x"18",	--877
		x"cc",	--878
		x"00",	--879
		x"8c",	--880
		x"02",	--881
		x"8c",	--882
		x"04",	--883
		x"1b",	--884
		x"82",	--885
		x"08",	--886
		x"0f",	--887
		x"3b",	--888
		x"30",	--889
		x"3f",	--890
		x"fc",	--891
		x"0b",	--892
		x"1b",	--893
		x"08",	--894
		x"1b",	--895
		x"0f",	--896
		x"5f",	--897
		x"18",	--898
		x"14",	--899
		x"3d",	--900
		x"1e",	--901
		x"0c",	--902
		x"05",	--903
		x"3d",	--904
		x"06",	--905
		x"cd",	--906
		x"fa",	--907
		x"0c",	--908
		x"1c",	--909
		x"0c",	--910
		x"f8",	--911
		x"30",	--912
		x"b7",	--913
		x"b0",	--914
		x"12",	--915
		x"21",	--916
		x"3f",	--917
		x"3b",	--918
		x"30",	--919
		x"0c",	--920
		x"0d",	--921
		x"0d",	--922
		x"0c",	--923
		x"0c",	--924
		x"3c",	--925
		x"18",	--926
		x"0f",	--927
		x"9c",	--928
		x"02",	--929
		x"3b",	--930
		x"30",	--931
		x"b2",	--932
		x"d2",	--933
		x"60",	--934
		x"b2",	--935
		x"b8",	--936
		x"72",	--937
		x"0f",	--938
		x"30",	--939
		x"0b",	--940
		x"0a",	--941
		x"0a",	--942
		x"1f",	--943
		x"0a",	--944
		x"3f",	--945
		x"20",	--946
		x"19",	--947
		x"0b",	--948
		x"0b",	--949
		x"0c",	--950
		x"0c",	--951
		x"0c",	--952
		x"0c",	--953
		x"3c",	--954
		x"d8",	--955
		x"8c",	--956
		x"00",	--957
		x"8c",	--958
		x"02",	--959
		x"8c",	--960
		x"04",	--961
		x"8c",	--962
		x"06",	--963
		x"8c",	--964
		x"08",	--965
		x"0e",	--966
		x"1e",	--967
		x"82",	--968
		x"0a",	--969
		x"3a",	--970
		x"3b",	--971
		x"30",	--972
		x"3f",	--973
		x"fb",	--974
		x"0f",	--975
		x"0e",	--976
		x"0e",	--977
		x"0e",	--978
		x"0e",	--979
		x"9e",	--980
		x"d8",	--981
		x"0f",	--982
		x"30",	--983
		x"0f",	--984
		x"0e",	--985
		x"0e",	--986
		x"0e",	--987
		x"0e",	--988
		x"8e",	--989
		x"d8",	--990
		x"0f",	--991
		x"30",	--992
		x"0f",	--993
		x"0e",	--994
		x"0d",	--995
		x"0c",	--996
		x"0b",	--997
		x"0a",	--998
		x"92",	--999
		x"0a",	--1000
		x"20",	--1001
		x"3b",	--1002
		x"da",	--1003
		x"0a",	--1004
		x"09",	--1005
		x"1f",	--1006
		x"8b",	--1007
		x"00",	--1008
		x"1a",	--1009
		x"3b",	--1010
		x"0a",	--1011
		x"1a",	--1012
		x"0a",	--1013
		x"13",	--1014
		x"8b",	--1015
		x"fe",	--1016
		x"f7",	--1017
		x"2f",	--1018
		x"1f",	--1019
		x"02",	--1020
		x"f0",	--1021
		x"8b",	--1022
		x"00",	--1023
		x"1f",	--1024
		x"06",	--1025
		x"9b",	--1026
		x"04",	--1027
		x"1a",	--1028
		x"3b",	--1029
		x"0a",	--1030
		x"1a",	--1031
		x"0a",	--1032
		x"ed",	--1033
		x"b2",	--1034
		x"fe",	--1035
		x"60",	--1036
		x"3a",	--1037
		x"3b",	--1038
		x"3c",	--1039
		x"3d",	--1040
		x"3e",	--1041
		x"3f",	--1042
		x"00",	--1043
		x"8f",	--1044
		x"00",	--1045
		x"0f",	--1046
		x"30",	--1047
		x"2f",	--1048
		x"2f",	--1049
		x"30",	--1050
		x"5e",	--1051
		x"81",	--1052
		x"3e",	--1053
		x"fc",	--1054
		x"c2",	--1055
		x"84",	--1056
		x"0f",	--1057
		x"30",	--1058
		x"3f",	--1059
		x"0f",	--1060
		x"5f",	--1061
		x"76",	--1062
		x"8f",	--1063
		x"b0",	--1064
		x"36",	--1065
		x"30",	--1066
		x"0b",	--1067
		x"0b",	--1068
		x"0e",	--1069
		x"0e",	--1070
		x"0e",	--1071
		x"0e",	--1072
		x"0e",	--1073
		x"0f",	--1074
		x"b0",	--1075
		x"46",	--1076
		x"0f",	--1077
		x"b0",	--1078
		x"46",	--1079
		x"3b",	--1080
		x"30",	--1081
		x"0b",	--1082
		x"0a",	--1083
		x"0a",	--1084
		x"3b",	--1085
		x"07",	--1086
		x"0e",	--1087
		x"4d",	--1088
		x"7d",	--1089
		x"0f",	--1090
		x"03",	--1091
		x"0e",	--1092
		x"7d",	--1093
		x"fd",	--1094
		x"1e",	--1095
		x"0a",	--1096
		x"3f",	--1097
		x"31",	--1098
		x"b0",	--1099
		x"36",	--1100
		x"3b",	--1101
		x"3b",	--1102
		x"ef",	--1103
		x"3a",	--1104
		x"3b",	--1105
		x"30",	--1106
		x"3f",	--1107
		x"30",	--1108
		x"f5",	--1109
		x"0b",	--1110
		x"0b",	--1111
		x"0e",	--1112
		x"8e",	--1113
		x"8e",	--1114
		x"0f",	--1115
		x"b0",	--1116
		x"56",	--1117
		x"0f",	--1118
		x"b0",	--1119
		x"56",	--1120
		x"3b",	--1121
		x"30",	--1122
		x"0b",	--1123
		x"0a",	--1124
		x"0a",	--1125
		x"0b",	--1126
		x"0d",	--1127
		x"8d",	--1128
		x"8d",	--1129
		x"0f",	--1130
		x"b0",	--1131
		x"56",	--1132
		x"0f",	--1133
		x"b0",	--1134
		x"56",	--1135
		x"0c",	--1136
		x"0d",	--1137
		x"8d",	--1138
		x"8c",	--1139
		x"4d",	--1140
		x"0d",	--1141
		x"0f",	--1142
		x"b0",	--1143
		x"56",	--1144
		x"0f",	--1145
		x"b0",	--1146
		x"56",	--1147
		x"3a",	--1148
		x"3b",	--1149
		x"30",	--1150
		x"0b",	--1151
		x"0a",	--1152
		x"09",	--1153
		x"0a",	--1154
		x"0e",	--1155
		x"19",	--1156
		x"09",	--1157
		x"39",	--1158
		x"0b",	--1159
		x"0d",	--1160
		x"0d",	--1161
		x"6f",	--1162
		x"8f",	--1163
		x"b0",	--1164
		x"56",	--1165
		x"0b",	--1166
		x"0e",	--1167
		x"1b",	--1168
		x"3b",	--1169
		x"07",	--1170
		x"05",	--1171
		x"3f",	--1172
		x"20",	--1173
		x"b0",	--1174
		x"36",	--1175
		x"ef",	--1176
		x"3f",	--1177
		x"3a",	--1178
		x"b0",	--1179
		x"36",	--1180
		x"ea",	--1181
		x"39",	--1182
		x"3a",	--1183
		x"3b",	--1184
		x"30",	--1185
		x"0b",	--1186
		x"0a",	--1187
		x"09",	--1188
		x"0a",	--1189
		x"0e",	--1190
		x"17",	--1191
		x"09",	--1192
		x"39",	--1193
		x"0b",	--1194
		x"6f",	--1195
		x"8f",	--1196
		x"b0",	--1197
		x"46",	--1198
		x"0b",	--1199
		x"0e",	--1200
		x"1b",	--1201
		x"3b",	--1202
		x"07",	--1203
		x"f6",	--1204
		x"3f",	--1205
		x"20",	--1206
		x"b0",	--1207
		x"36",	--1208
		x"6f",	--1209
		x"8f",	--1210
		x"b0",	--1211
		x"46",	--1212
		x"0b",	--1213
		x"f2",	--1214
		x"39",	--1215
		x"3a",	--1216
		x"3b",	--1217
		x"30",	--1218
		x"0b",	--1219
		x"0a",	--1220
		x"09",	--1221
		x"31",	--1222
		x"ec",	--1223
		x"0b",	--1224
		x"0f",	--1225
		x"34",	--1226
		x"3b",	--1227
		x"0a",	--1228
		x"38",	--1229
		x"09",	--1230
		x"0a",	--1231
		x"0a",	--1232
		x"3e",	--1233
		x"0a",	--1234
		x"0f",	--1235
		x"b0",	--1236
		x"a2",	--1237
		x"7f",	--1238
		x"30",	--1239
		x"ca",	--1240
		x"00",	--1241
		x"19",	--1242
		x"3e",	--1243
		x"0a",	--1244
		x"0f",	--1245
		x"b0",	--1246
		x"70",	--1247
		x"0b",	--1248
		x"3f",	--1249
		x"0a",	--1250
		x"eb",	--1251
		x"0a",	--1252
		x"1a",	--1253
		x"09",	--1254
		x"3e",	--1255
		x"0a",	--1256
		x"0f",	--1257
		x"b0",	--1258
		x"a2",	--1259
		x"7f",	--1260
		x"30",	--1261
		x"c9",	--1262
		x"00",	--1263
		x"3a",	--1264
		x"0f",	--1265
		x"0f",	--1266
		x"6f",	--1267
		x"8f",	--1268
		x"b0",	--1269
		x"36",	--1270
		x"0a",	--1271
		x"f7",	--1272
		x"31",	--1273
		x"14",	--1274
		x"39",	--1275
		x"3a",	--1276
		x"3b",	--1277
		x"30",	--1278
		x"3f",	--1279
		x"2d",	--1280
		x"b0",	--1281
		x"36",	--1282
		x"3b",	--1283
		x"1b",	--1284
		x"c5",	--1285
		x"1a",	--1286
		x"09",	--1287
		x"dd",	--1288
		x"0b",	--1289
		x"0a",	--1290
		x"09",	--1291
		x"0b",	--1292
		x"3b",	--1293
		x"39",	--1294
		x"6f",	--1295
		x"4f",	--1296
		x"0b",	--1297
		x"1a",	--1298
		x"8f",	--1299
		x"b0",	--1300
		x"36",	--1301
		x"0a",	--1302
		x"09",	--1303
		x"19",	--1304
		x"5f",	--1305
		x"01",	--1306
		x"4f",	--1307
		x"10",	--1308
		x"7f",	--1309
		x"25",	--1310
		x"f3",	--1311
		x"0a",	--1312
		x"1a",	--1313
		x"5f",	--1314
		x"01",	--1315
		x"7f",	--1316
		x"db",	--1317
		x"7f",	--1318
		x"54",	--1319
		x"ee",	--1320
		x"4f",	--1321
		x"0f",	--1322
		x"10",	--1323
		x"ce",	--1324
		x"39",	--1325
		x"3a",	--1326
		x"3b",	--1327
		x"30",	--1328
		x"09",	--1329
		x"29",	--1330
		x"1e",	--1331
		x"02",	--1332
		x"2f",	--1333
		x"b0",	--1334
		x"fe",	--1335
		x"0b",	--1336
		x"dd",	--1337
		x"09",	--1338
		x"29",	--1339
		x"2f",	--1340
		x"b0",	--1341
		x"ac",	--1342
		x"0b",	--1343
		x"d6",	--1344
		x"0f",	--1345
		x"2b",	--1346
		x"29",	--1347
		x"6f",	--1348
		x"4f",	--1349
		x"d0",	--1350
		x"19",	--1351
		x"8f",	--1352
		x"b0",	--1353
		x"36",	--1354
		x"7f",	--1355
		x"4f",	--1356
		x"fa",	--1357
		x"c8",	--1358
		x"09",	--1359
		x"29",	--1360
		x"1e",	--1361
		x"02",	--1362
		x"2f",	--1363
		x"b0",	--1364
		x"44",	--1365
		x"0b",	--1366
		x"bf",	--1367
		x"09",	--1368
		x"29",	--1369
		x"2e",	--1370
		x"0f",	--1371
		x"8f",	--1372
		x"8f",	--1373
		x"8f",	--1374
		x"8f",	--1375
		x"b0",	--1376
		x"c6",	--1377
		x"0b",	--1378
		x"b3",	--1379
		x"09",	--1380
		x"29",	--1381
		x"2f",	--1382
		x"b0",	--1383
		x"86",	--1384
		x"0b",	--1385
		x"ac",	--1386
		x"09",	--1387
		x"29",	--1388
		x"2f",	--1389
		x"b0",	--1390
		x"36",	--1391
		x"0b",	--1392
		x"a5",	--1393
		x"09",	--1394
		x"29",	--1395
		x"2f",	--1396
		x"b0",	--1397
		x"56",	--1398
		x"0b",	--1399
		x"9e",	--1400
		x"09",	--1401
		x"29",	--1402
		x"2f",	--1403
		x"b0",	--1404
		x"74",	--1405
		x"0b",	--1406
		x"97",	--1407
		x"3f",	--1408
		x"25",	--1409
		x"b0",	--1410
		x"36",	--1411
		x"92",	--1412
		x"0f",	--1413
		x"0e",	--1414
		x"1f",	--1415
		x"0c",	--1416
		x"df",	--1417
		x"85",	--1418
		x"18",	--1419
		x"1f",	--1420
		x"0c",	--1421
		x"3f",	--1422
		x"3f",	--1423
		x"13",	--1424
		x"92",	--1425
		x"0c",	--1426
		x"1e",	--1427
		x"0c",	--1428
		x"1f",	--1429
		x"0e",	--1430
		x"0e",	--1431
		x"02",	--1432
		x"92",	--1433
		x"0e",	--1434
		x"f2",	--1435
		x"10",	--1436
		x"81",	--1437
		x"3e",	--1438
		x"3f",	--1439
		x"b1",	--1440
		x"f0",	--1441
		x"00",	--1442
		x"00",	--1443
		x"82",	--1444
		x"0c",	--1445
		x"ec",	--1446
		x"b2",	--1447
		x"c3",	--1448
		x"82",	--1449
		x"f2",	--1450
		x"11",	--1451
		x"80",	--1452
		x"30",	--1453
		x"1e",	--1454
		x"0c",	--1455
		x"1f",	--1456
		x"0e",	--1457
		x"0e",	--1458
		x"05",	--1459
		x"1f",	--1460
		x"0c",	--1461
		x"1f",	--1462
		x"0e",	--1463
		x"30",	--1464
		x"1d",	--1465
		x"0c",	--1466
		x"1e",	--1467
		x"0e",	--1468
		x"3f",	--1469
		x"40",	--1470
		x"0f",	--1471
		x"0f",	--1472
		x"30",	--1473
		x"1f",	--1474
		x"0e",	--1475
		x"5f",	--1476
		x"18",	--1477
		x"1d",	--1478
		x"0e",	--1479
		x"1e",	--1480
		x"0c",	--1481
		x"0d",	--1482
		x"0b",	--1483
		x"1e",	--1484
		x"0e",	--1485
		x"3e",	--1486
		x"3f",	--1487
		x"03",	--1488
		x"82",	--1489
		x"0e",	--1490
		x"30",	--1491
		x"92",	--1492
		x"0e",	--1493
		x"30",	--1494
		x"4f",	--1495
		x"30",	--1496
		x"0b",	--1497
		x"0a",	--1498
		x"0a",	--1499
		x"0b",	--1500
		x"0c",	--1501
		x"3d",	--1502
		x"00",	--1503
		x"b0",	--1504
		x"96",	--1505
		x"0f",	--1506
		x"07",	--1507
		x"0e",	--1508
		x"0f",	--1509
		x"b0",	--1510
		x"e6",	--1511
		x"3a",	--1512
		x"3b",	--1513
		x"30",	--1514
		x"0c",	--1515
		x"3d",	--1516
		x"00",	--1517
		x"0e",	--1518
		x"0f",	--1519
		x"b0",	--1520
		x"d2",	--1521
		x"b0",	--1522
		x"e6",	--1523
		x"0e",	--1524
		x"3f",	--1525
		x"00",	--1526
		x"3a",	--1527
		x"3b",	--1528
		x"30",	--1529
		x"0b",	--1530
		x"0a",	--1531
		x"09",	--1532
		x"08",	--1533
		x"07",	--1534
		x"06",	--1535
		x"05",	--1536
		x"04",	--1537
		x"31",	--1538
		x"fa",	--1539
		x"08",	--1540
		x"6b",	--1541
		x"6b",	--1542
		x"67",	--1543
		x"6c",	--1544
		x"6c",	--1545
		x"e9",	--1546
		x"6b",	--1547
		x"02",	--1548
		x"30",	--1549
		x"74",	--1550
		x"6c",	--1551
		x"e3",	--1552
		x"6c",	--1553
		x"bb",	--1554
		x"6b",	--1555
		x"df",	--1556
		x"91",	--1557
		x"02",	--1558
		x"00",	--1559
		x"1b",	--1560
		x"02",	--1561
		x"14",	--1562
		x"04",	--1563
		x"15",	--1564
		x"06",	--1565
		x"16",	--1566
		x"04",	--1567
		x"17",	--1568
		x"06",	--1569
		x"2c",	--1570
		x"0c",	--1571
		x"09",	--1572
		x"0c",	--1573
		x"bf",	--1574
		x"39",	--1575
		x"20",	--1576
		x"50",	--1577
		x"1c",	--1578
		x"d7",	--1579
		x"81",	--1580
		x"02",	--1581
		x"81",	--1582
		x"04",	--1583
		x"4c",	--1584
		x"7c",	--1585
		x"1f",	--1586
		x"0b",	--1587
		x"0a",	--1588
		x"0b",	--1589
		x"12",	--1590
		x"0b",	--1591
		x"0a",	--1592
		x"7c",	--1593
		x"fb",	--1594
		x"81",	--1595
		x"02",	--1596
		x"81",	--1597
		x"04",	--1598
		x"1c",	--1599
		x"0d",	--1600
		x"79",	--1601
		x"1f",	--1602
		x"04",	--1603
		x"0c",	--1604
		x"0d",	--1605
		x"79",	--1606
		x"fc",	--1607
		x"3c",	--1608
		x"3d",	--1609
		x"0c",	--1610
		x"0d",	--1611
		x"1a",	--1612
		x"0b",	--1613
		x"0c",	--1614
		x"02",	--1615
		x"0d",	--1616
		x"e5",	--1617
		x"16",	--1618
		x"02",	--1619
		x"17",	--1620
		x"04",	--1621
		x"06",	--1622
		x"07",	--1623
		x"5f",	--1624
		x"01",	--1625
		x"5f",	--1626
		x"01",	--1627
		x"28",	--1628
		x"c8",	--1629
		x"01",	--1630
		x"a8",	--1631
		x"02",	--1632
		x"0e",	--1633
		x"0f",	--1634
		x"0e",	--1635
		x"0f",	--1636
		x"88",	--1637
		x"04",	--1638
		x"88",	--1639
		x"06",	--1640
		x"f8",	--1641
		x"03",	--1642
		x"00",	--1643
		x"0f",	--1644
		x"4d",	--1645
		x"0f",	--1646
		x"31",	--1647
		x"06",	--1648
		x"34",	--1649
		x"35",	--1650
		x"36",	--1651
		x"37",	--1652
		x"38",	--1653
		x"39",	--1654
		x"3a",	--1655
		x"3b",	--1656
		x"30",	--1657
		x"2b",	--1658
		x"67",	--1659
		x"81",	--1660
		x"00",	--1661
		x"04",	--1662
		x"05",	--1663
		x"5f",	--1664
		x"01",	--1665
		x"5f",	--1666
		x"01",	--1667
		x"d8",	--1668
		x"4f",	--1669
		x"68",	--1670
		x"0e",	--1671
		x"0f",	--1672
		x"0e",	--1673
		x"0f",	--1674
		x"0f",	--1675
		x"69",	--1676
		x"c8",	--1677
		x"01",	--1678
		x"a8",	--1679
		x"02",	--1680
		x"88",	--1681
		x"04",	--1682
		x"88",	--1683
		x"06",	--1684
		x"0c",	--1685
		x"0d",	--1686
		x"3c",	--1687
		x"3d",	--1688
		x"3d",	--1689
		x"ff",	--1690
		x"05",	--1691
		x"3d",	--1692
		x"00",	--1693
		x"17",	--1694
		x"3c",	--1695
		x"15",	--1696
		x"1b",	--1697
		x"02",	--1698
		x"3b",	--1699
		x"0e",	--1700
		x"0f",	--1701
		x"0a",	--1702
		x"3b",	--1703
		x"0c",	--1704
		x"0d",	--1705
		x"3c",	--1706
		x"3d",	--1707
		x"3d",	--1708
		x"ff",	--1709
		x"f5",	--1710
		x"3c",	--1711
		x"88",	--1712
		x"04",	--1713
		x"88",	--1714
		x"06",	--1715
		x"88",	--1716
		x"02",	--1717
		x"f8",	--1718
		x"03",	--1719
		x"00",	--1720
		x"0f",	--1721
		x"b3",	--1722
		x"0c",	--1723
		x"0d",	--1724
		x"1c",	--1725
		x"0d",	--1726
		x"12",	--1727
		x"0f",	--1728
		x"0e",	--1729
		x"0a",	--1730
		x"0b",	--1731
		x"0a",	--1732
		x"0b",	--1733
		x"88",	--1734
		x"04",	--1735
		x"88",	--1736
		x"06",	--1737
		x"98",	--1738
		x"02",	--1739
		x"0f",	--1740
		x"a1",	--1741
		x"6b",	--1742
		x"9f",	--1743
		x"ad",	--1744
		x"00",	--1745
		x"9d",	--1746
		x"02",	--1747
		x"02",	--1748
		x"9d",	--1749
		x"04",	--1750
		x"04",	--1751
		x"9d",	--1752
		x"06",	--1753
		x"06",	--1754
		x"5e",	--1755
		x"01",	--1756
		x"5e",	--1757
		x"01",	--1758
		x"cd",	--1759
		x"01",	--1760
		x"0f",	--1761
		x"8c",	--1762
		x"06",	--1763
		x"07",	--1764
		x"9a",	--1765
		x"39",	--1766
		x"19",	--1767
		x"39",	--1768
		x"20",	--1769
		x"8f",	--1770
		x"3e",	--1771
		x"3c",	--1772
		x"b6",	--1773
		x"c1",	--1774
		x"0e",	--1775
		x"0f",	--1776
		x"0e",	--1777
		x"0f",	--1778
		x"97",	--1779
		x"0f",	--1780
		x"79",	--1781
		x"d8",	--1782
		x"01",	--1783
		x"a8",	--1784
		x"02",	--1785
		x"3e",	--1786
		x"3f",	--1787
		x"1e",	--1788
		x"0f",	--1789
		x"88",	--1790
		x"04",	--1791
		x"88",	--1792
		x"06",	--1793
		x"92",	--1794
		x"0c",	--1795
		x"7b",	--1796
		x"81",	--1797
		x"00",	--1798
		x"81",	--1799
		x"02",	--1800
		x"81",	--1801
		x"04",	--1802
		x"4d",	--1803
		x"7d",	--1804
		x"1f",	--1805
		x"0c",	--1806
		x"4b",	--1807
		x"0c",	--1808
		x"0d",	--1809
		x"12",	--1810
		x"0d",	--1811
		x"0c",	--1812
		x"7b",	--1813
		x"fb",	--1814
		x"81",	--1815
		x"02",	--1816
		x"81",	--1817
		x"04",	--1818
		x"1c",	--1819
		x"0d",	--1820
		x"79",	--1821
		x"1f",	--1822
		x"04",	--1823
		x"0c",	--1824
		x"0d",	--1825
		x"79",	--1826
		x"fc",	--1827
		x"3c",	--1828
		x"3d",	--1829
		x"0c",	--1830
		x"0d",	--1831
		x"1a",	--1832
		x"0b",	--1833
		x"0c",	--1834
		x"04",	--1835
		x"0d",	--1836
		x"02",	--1837
		x"0a",	--1838
		x"0b",	--1839
		x"14",	--1840
		x"02",	--1841
		x"15",	--1842
		x"04",	--1843
		x"04",	--1844
		x"05",	--1845
		x"49",	--1846
		x"0a",	--1847
		x"0b",	--1848
		x"18",	--1849
		x"6c",	--1850
		x"33",	--1851
		x"df",	--1852
		x"01",	--1853
		x"01",	--1854
		x"2f",	--1855
		x"3f",	--1856
		x"88",	--1857
		x"2c",	--1858
		x"31",	--1859
		x"e0",	--1860
		x"81",	--1861
		x"04",	--1862
		x"81",	--1863
		x"06",	--1864
		x"81",	--1865
		x"00",	--1866
		x"81",	--1867
		x"02",	--1868
		x"0e",	--1869
		x"3e",	--1870
		x"18",	--1871
		x"0f",	--1872
		x"2f",	--1873
		x"b0",	--1874
		x"a8",	--1875
		x"0e",	--1876
		x"3e",	--1877
		x"10",	--1878
		x"0f",	--1879
		x"b0",	--1880
		x"a8",	--1881
		x"0d",	--1882
		x"3d",	--1883
		x"0e",	--1884
		x"3e",	--1885
		x"10",	--1886
		x"0f",	--1887
		x"3f",	--1888
		x"18",	--1889
		x"b0",	--1890
		x"f4",	--1891
		x"b0",	--1892
		x"ca",	--1893
		x"31",	--1894
		x"20",	--1895
		x"30",	--1896
		x"31",	--1897
		x"e0",	--1898
		x"81",	--1899
		x"04",	--1900
		x"81",	--1901
		x"06",	--1902
		x"81",	--1903
		x"00",	--1904
		x"81",	--1905
		x"02",	--1906
		x"0e",	--1907
		x"3e",	--1908
		x"18",	--1909
		x"0f",	--1910
		x"2f",	--1911
		x"b0",	--1912
		x"a8",	--1913
		x"0e",	--1914
		x"3e",	--1915
		x"10",	--1916
		x"0f",	--1917
		x"b0",	--1918
		x"a8",	--1919
		x"d1",	--1920
		x"11",	--1921
		x"0d",	--1922
		x"3d",	--1923
		x"0e",	--1924
		x"3e",	--1925
		x"10",	--1926
		x"0f",	--1927
		x"3f",	--1928
		x"18",	--1929
		x"b0",	--1930
		x"f4",	--1931
		x"b0",	--1932
		x"ca",	--1933
		x"31",	--1934
		x"20",	--1935
		x"30",	--1936
		x"0b",	--1937
		x"0a",	--1938
		x"09",	--1939
		x"08",	--1940
		x"07",	--1941
		x"06",	--1942
		x"05",	--1943
		x"04",	--1944
		x"31",	--1945
		x"dc",	--1946
		x"81",	--1947
		x"04",	--1948
		x"81",	--1949
		x"06",	--1950
		x"81",	--1951
		x"00",	--1952
		x"81",	--1953
		x"02",	--1954
		x"0e",	--1955
		x"3e",	--1956
		x"18",	--1957
		x"0f",	--1958
		x"2f",	--1959
		x"b0",	--1960
		x"a8",	--1961
		x"0e",	--1962
		x"3e",	--1963
		x"10",	--1964
		x"0f",	--1965
		x"b0",	--1966
		x"a8",	--1967
		x"5f",	--1968
		x"18",	--1969
		x"6f",	--1970
		x"b6",	--1971
		x"5e",	--1972
		x"10",	--1973
		x"6e",	--1974
		x"d9",	--1975
		x"6f",	--1976
		x"ae",	--1977
		x"6e",	--1978
		x"e2",	--1979
		x"6f",	--1980
		x"ac",	--1981
		x"6e",	--1982
		x"d1",	--1983
		x"14",	--1984
		x"1c",	--1985
		x"15",	--1986
		x"1e",	--1987
		x"18",	--1988
		x"14",	--1989
		x"19",	--1990
		x"16",	--1991
		x"3c",	--1992
		x"20",	--1993
		x"0e",	--1994
		x"0f",	--1995
		x"06",	--1996
		x"07",	--1997
		x"81",	--1998
		x"20",	--1999
		x"81",	--2000
		x"22",	--2001
		x"0a",	--2002
		x"0b",	--2003
		x"81",	--2004
		x"20",	--2005
		x"08",	--2006
		x"08",	--2007
		x"09",	--2008
		x"12",	--2009
		x"05",	--2010
		x"04",	--2011
		x"b1",	--2012
		x"20",	--2013
		x"19",	--2014
		x"14",	--2015
		x"0d",	--2016
		x"0a",	--2017
		x"0b",	--2018
		x"0e",	--2019
		x"0f",	--2020
		x"1c",	--2021
		x"0d",	--2022
		x"0b",	--2023
		x"03",	--2024
		x"0b",	--2025
		x"0c",	--2026
		x"0d",	--2027
		x"0e",	--2028
		x"0f",	--2029
		x"06",	--2030
		x"07",	--2031
		x"09",	--2032
		x"e5",	--2033
		x"16",	--2034
		x"07",	--2035
		x"e2",	--2036
		x"0a",	--2037
		x"f5",	--2038
		x"f2",	--2039
		x"81",	--2040
		x"20",	--2041
		x"81",	--2042
		x"22",	--2043
		x"0c",	--2044
		x"1a",	--2045
		x"1a",	--2046
		x"1a",	--2047
		x"12",	--2048
		x"06",	--2049
		x"26",	--2050
		x"81",	--2051
		x"0a",	--2052
		x"5d",	--2053
		x"d1",	--2054
		x"11",	--2055
		x"19",	--2056
		x"83",	--2057
		x"c1",	--2058
		x"09",	--2059
		x"0c",	--2060
		x"3c",	--2061
		x"3f",	--2062
		x"00",	--2063
		x"18",	--2064
		x"1d",	--2065
		x"0a",	--2066
		x"3d",	--2067
		x"1a",	--2068
		x"20",	--2069
		x"1b",	--2070
		x"22",	--2071
		x"0c",	--2072
		x"0e",	--2073
		x"0f",	--2074
		x"0b",	--2075
		x"2a",	--2076
		x"0a",	--2077
		x"0b",	--2078
		x"3d",	--2079
		x"3f",	--2080
		x"00",	--2081
		x"f5",	--2082
		x"81",	--2083
		x"20",	--2084
		x"81",	--2085
		x"22",	--2086
		x"81",	--2087
		x"0a",	--2088
		x"0c",	--2089
		x"0d",	--2090
		x"3c",	--2091
		x"7f",	--2092
		x"0d",	--2093
		x"3c",	--2094
		x"40",	--2095
		x"44",	--2096
		x"81",	--2097
		x"0c",	--2098
		x"81",	--2099
		x"0e",	--2100
		x"f1",	--2101
		x"03",	--2102
		x"08",	--2103
		x"0f",	--2104
		x"3f",	--2105
		x"b0",	--2106
		x"ca",	--2107
		x"31",	--2108
		x"24",	--2109
		x"34",	--2110
		x"35",	--2111
		x"36",	--2112
		x"37",	--2113
		x"38",	--2114
		x"39",	--2115
		x"3a",	--2116
		x"3b",	--2117
		x"30",	--2118
		x"1e",	--2119
		x"0f",	--2120
		x"d3",	--2121
		x"3a",	--2122
		x"03",	--2123
		x"08",	--2124
		x"1e",	--2125
		x"10",	--2126
		x"1c",	--2127
		x"20",	--2128
		x"1d",	--2129
		x"22",	--2130
		x"12",	--2131
		x"0d",	--2132
		x"0c",	--2133
		x"06",	--2134
		x"07",	--2135
		x"06",	--2136
		x"37",	--2137
		x"00",	--2138
		x"81",	--2139
		x"20",	--2140
		x"81",	--2141
		x"22",	--2142
		x"12",	--2143
		x"0f",	--2144
		x"0e",	--2145
		x"1a",	--2146
		x"0f",	--2147
		x"e7",	--2148
		x"81",	--2149
		x"0a",	--2150
		x"a6",	--2151
		x"6e",	--2152
		x"36",	--2153
		x"5f",	--2154
		x"d1",	--2155
		x"11",	--2156
		x"19",	--2157
		x"20",	--2158
		x"c1",	--2159
		x"19",	--2160
		x"0f",	--2161
		x"3f",	--2162
		x"18",	--2163
		x"c5",	--2164
		x"0d",	--2165
		x"ba",	--2166
		x"0c",	--2167
		x"0d",	--2168
		x"3c",	--2169
		x"80",	--2170
		x"0d",	--2171
		x"0c",	--2172
		x"b3",	--2173
		x"0d",	--2174
		x"b1",	--2175
		x"81",	--2176
		x"20",	--2177
		x"03",	--2178
		x"81",	--2179
		x"22",	--2180
		x"ab",	--2181
		x"3e",	--2182
		x"40",	--2183
		x"0f",	--2184
		x"3e",	--2185
		x"80",	--2186
		x"3f",	--2187
		x"a4",	--2188
		x"4d",	--2189
		x"7b",	--2190
		x"4f",	--2191
		x"de",	--2192
		x"5f",	--2193
		x"d1",	--2194
		x"11",	--2195
		x"19",	--2196
		x"06",	--2197
		x"c1",	--2198
		x"11",	--2199
		x"0f",	--2200
		x"3f",	--2201
		x"10",	--2202
		x"9e",	--2203
		x"4f",	--2204
		x"f8",	--2205
		x"6f",	--2206
		x"f1",	--2207
		x"3f",	--2208
		x"88",	--2209
		x"97",	--2210
		x"0b",	--2211
		x"0a",	--2212
		x"09",	--2213
		x"08",	--2214
		x"07",	--2215
		x"31",	--2216
		x"e8",	--2217
		x"81",	--2218
		x"04",	--2219
		x"81",	--2220
		x"06",	--2221
		x"81",	--2222
		x"00",	--2223
		x"81",	--2224
		x"02",	--2225
		x"0e",	--2226
		x"3e",	--2227
		x"10",	--2228
		x"0f",	--2229
		x"2f",	--2230
		x"b0",	--2231
		x"a8",	--2232
		x"0e",	--2233
		x"3e",	--2234
		x"0f",	--2235
		x"b0",	--2236
		x"a8",	--2237
		x"5f",	--2238
		x"10",	--2239
		x"6f",	--2240
		x"5d",	--2241
		x"5e",	--2242
		x"08",	--2243
		x"6e",	--2244
		x"82",	--2245
		x"d1",	--2246
		x"09",	--2247
		x"11",	--2248
		x"6f",	--2249
		x"58",	--2250
		x"6f",	--2251
		x"56",	--2252
		x"6e",	--2253
		x"6f",	--2254
		x"6e",	--2255
		x"4c",	--2256
		x"1d",	--2257
		x"12",	--2258
		x"1d",	--2259
		x"0a",	--2260
		x"81",	--2261
		x"12",	--2262
		x"1e",	--2263
		x"14",	--2264
		x"1f",	--2265
		x"16",	--2266
		x"18",	--2267
		x"0c",	--2268
		x"19",	--2269
		x"0e",	--2270
		x"0f",	--2271
		x"1e",	--2272
		x"0e",	--2273
		x"0f",	--2274
		x"3d",	--2275
		x"81",	--2276
		x"12",	--2277
		x"37",	--2278
		x"1f",	--2279
		x"0c",	--2280
		x"3d",	--2281
		x"00",	--2282
		x"0a",	--2283
		x"0b",	--2284
		x"0b",	--2285
		x"0a",	--2286
		x"0b",	--2287
		x"0e",	--2288
		x"0f",	--2289
		x"12",	--2290
		x"0d",	--2291
		x"0c",	--2292
		x"0e",	--2293
		x"0f",	--2294
		x"37",	--2295
		x"0b",	--2296
		x"0f",	--2297
		x"f7",	--2298
		x"f2",	--2299
		x"0e",	--2300
		x"f4",	--2301
		x"ef",	--2302
		x"09",	--2303
		x"e5",	--2304
		x"0e",	--2305
		x"e3",	--2306
		x"dd",	--2307
		x"0c",	--2308
		x"0d",	--2309
		x"3c",	--2310
		x"7f",	--2311
		x"0d",	--2312
		x"3c",	--2313
		x"40",	--2314
		x"1c",	--2315
		x"81",	--2316
		x"14",	--2317
		x"81",	--2318
		x"16",	--2319
		x"0f",	--2320
		x"3f",	--2321
		x"10",	--2322
		x"b0",	--2323
		x"ca",	--2324
		x"31",	--2325
		x"18",	--2326
		x"37",	--2327
		x"38",	--2328
		x"39",	--2329
		x"3a",	--2330
		x"3b",	--2331
		x"30",	--2332
		x"e1",	--2333
		x"10",	--2334
		x"0f",	--2335
		x"3f",	--2336
		x"10",	--2337
		x"f0",	--2338
		x"4f",	--2339
		x"fa",	--2340
		x"3f",	--2341
		x"88",	--2342
		x"eb",	--2343
		x"0d",	--2344
		x"e2",	--2345
		x"0c",	--2346
		x"0d",	--2347
		x"3c",	--2348
		x"80",	--2349
		x"0d",	--2350
		x"0c",	--2351
		x"db",	--2352
		x"0d",	--2353
		x"d9",	--2354
		x"0e",	--2355
		x"02",	--2356
		x"0f",	--2357
		x"d5",	--2358
		x"3a",	--2359
		x"40",	--2360
		x"0b",	--2361
		x"3a",	--2362
		x"80",	--2363
		x"3b",	--2364
		x"ce",	--2365
		x"81",	--2366
		x"14",	--2367
		x"81",	--2368
		x"16",	--2369
		x"81",	--2370
		x"12",	--2371
		x"0f",	--2372
		x"3f",	--2373
		x"10",	--2374
		x"cb",	--2375
		x"0f",	--2376
		x"3f",	--2377
		x"c8",	--2378
		x"31",	--2379
		x"e8",	--2380
		x"81",	--2381
		x"04",	--2382
		x"81",	--2383
		x"06",	--2384
		x"81",	--2385
		x"00",	--2386
		x"81",	--2387
		x"02",	--2388
		x"0e",	--2389
		x"3e",	--2390
		x"10",	--2391
		x"0f",	--2392
		x"2f",	--2393
		x"b0",	--2394
		x"a8",	--2395
		x"0e",	--2396
		x"3e",	--2397
		x"0f",	--2398
		x"b0",	--2399
		x"a8",	--2400
		x"e1",	--2401
		x"10",	--2402
		x"0d",	--2403
		x"e1",	--2404
		x"08",	--2405
		x"0a",	--2406
		x"0e",	--2407
		x"3e",	--2408
		x"0f",	--2409
		x"3f",	--2410
		x"10",	--2411
		x"b0",	--2412
		x"cc",	--2413
		x"31",	--2414
		x"18",	--2415
		x"30",	--2416
		x"3f",	--2417
		x"fb",	--2418
		x"31",	--2419
		x"f4",	--2420
		x"81",	--2421
		x"00",	--2422
		x"81",	--2423
		x"02",	--2424
		x"0e",	--2425
		x"2e",	--2426
		x"0f",	--2427
		x"b0",	--2428
		x"a8",	--2429
		x"5f",	--2430
		x"04",	--2431
		x"6f",	--2432
		x"28",	--2433
		x"27",	--2434
		x"6f",	--2435
		x"07",	--2436
		x"1d",	--2437
		x"06",	--2438
		x"0d",	--2439
		x"21",	--2440
		x"3d",	--2441
		x"1f",	--2442
		x"09",	--2443
		x"c1",	--2444
		x"05",	--2445
		x"26",	--2446
		x"3e",	--2447
		x"3f",	--2448
		x"ff",	--2449
		x"31",	--2450
		x"0c",	--2451
		x"30",	--2452
		x"1e",	--2453
		x"08",	--2454
		x"1f",	--2455
		x"0a",	--2456
		x"3c",	--2457
		x"1e",	--2458
		x"4c",	--2459
		x"4d",	--2460
		x"7d",	--2461
		x"1f",	--2462
		x"0f",	--2463
		x"c1",	--2464
		x"05",	--2465
		x"ef",	--2466
		x"3e",	--2467
		x"3f",	--2468
		x"1e",	--2469
		x"0f",	--2470
		x"31",	--2471
		x"0c",	--2472
		x"30",	--2473
		x"0e",	--2474
		x"0f",	--2475
		x"31",	--2476
		x"0c",	--2477
		x"30",	--2478
		x"12",	--2479
		x"0f",	--2480
		x"0e",	--2481
		x"7d",	--2482
		x"fb",	--2483
		x"eb",	--2484
		x"0e",	--2485
		x"3f",	--2486
		x"00",	--2487
		x"31",	--2488
		x"0c",	--2489
		x"30",	--2490
		x"0b",	--2491
		x"0a",	--2492
		x"09",	--2493
		x"08",	--2494
		x"31",	--2495
		x"0a",	--2496
		x"0b",	--2497
		x"c1",	--2498
		x"01",	--2499
		x"0e",	--2500
		x"0d",	--2501
		x"0b",	--2502
		x"0b",	--2503
		x"e1",	--2504
		x"00",	--2505
		x"0f",	--2506
		x"b0",	--2507
		x"ca",	--2508
		x"31",	--2509
		x"38",	--2510
		x"39",	--2511
		x"3a",	--2512
		x"3b",	--2513
		x"30",	--2514
		x"f1",	--2515
		x"03",	--2516
		x"00",	--2517
		x"b1",	--2518
		x"1e",	--2519
		x"02",	--2520
		x"81",	--2521
		x"04",	--2522
		x"81",	--2523
		x"06",	--2524
		x"0e",	--2525
		x"0f",	--2526
		x"b0",	--2527
		x"58",	--2528
		x"3f",	--2529
		x"0f",	--2530
		x"18",	--2531
		x"e5",	--2532
		x"81",	--2533
		x"04",	--2534
		x"81",	--2535
		x"06",	--2536
		x"4e",	--2537
		x"7e",	--2538
		x"1f",	--2539
		x"06",	--2540
		x"3e",	--2541
		x"1e",	--2542
		x"0e",	--2543
		x"81",	--2544
		x"02",	--2545
		x"d7",	--2546
		x"91",	--2547
		x"04",	--2548
		x"04",	--2549
		x"91",	--2550
		x"06",	--2551
		x"06",	--2552
		x"7e",	--2553
		x"f8",	--2554
		x"f1",	--2555
		x"0e",	--2556
		x"3e",	--2557
		x"1e",	--2558
		x"1c",	--2559
		x"0d",	--2560
		x"48",	--2561
		x"78",	--2562
		x"1f",	--2563
		x"04",	--2564
		x"0c",	--2565
		x"0d",	--2566
		x"78",	--2567
		x"fc",	--2568
		x"3c",	--2569
		x"3d",	--2570
		x"0c",	--2571
		x"0d",	--2572
		x"18",	--2573
		x"09",	--2574
		x"0c",	--2575
		x"04",	--2576
		x"0d",	--2577
		x"02",	--2578
		x"08",	--2579
		x"09",	--2580
		x"7e",	--2581
		x"1f",	--2582
		x"0e",	--2583
		x"0d",	--2584
		x"0e",	--2585
		x"0d",	--2586
		x"0e",	--2587
		x"81",	--2588
		x"04",	--2589
		x"81",	--2590
		x"06",	--2591
		x"3e",	--2592
		x"1e",	--2593
		x"0e",	--2594
		x"81",	--2595
		x"02",	--2596
		x"a4",	--2597
		x"12",	--2598
		x"0b",	--2599
		x"0a",	--2600
		x"7e",	--2601
		x"fb",	--2602
		x"ec",	--2603
		x"0b",	--2604
		x"0a",	--2605
		x"09",	--2606
		x"1f",	--2607
		x"17",	--2608
		x"3e",	--2609
		x"00",	--2610
		x"2c",	--2611
		x"3a",	--2612
		x"18",	--2613
		x"0b",	--2614
		x"39",	--2615
		x"0c",	--2616
		x"0d",	--2617
		x"4f",	--2618
		x"4f",	--2619
		x"17",	--2620
		x"3c",	--2621
		x"90",	--2622
		x"6e",	--2623
		x"0f",	--2624
		x"0a",	--2625
		x"0b",	--2626
		x"0f",	--2627
		x"39",	--2628
		x"3a",	--2629
		x"3b",	--2630
		x"30",	--2631
		x"3f",	--2632
		x"00",	--2633
		x"0f",	--2634
		x"3a",	--2635
		x"0b",	--2636
		x"39",	--2637
		x"18",	--2638
		x"0c",	--2639
		x"0d",	--2640
		x"4f",	--2641
		x"4f",	--2642
		x"e9",	--2643
		x"12",	--2644
		x"0d",	--2645
		x"0c",	--2646
		x"7f",	--2647
		x"fb",	--2648
		x"e3",	--2649
		x"3a",	--2650
		x"10",	--2651
		x"0b",	--2652
		x"39",	--2653
		x"10",	--2654
		x"ef",	--2655
		x"3a",	--2656
		x"20",	--2657
		x"0b",	--2658
		x"09",	--2659
		x"ea",	--2660
		x"0b",	--2661
		x"0a",	--2662
		x"09",	--2663
		x"08",	--2664
		x"07",	--2665
		x"0d",	--2666
		x"1e",	--2667
		x"04",	--2668
		x"1f",	--2669
		x"06",	--2670
		x"5a",	--2671
		x"01",	--2672
		x"6c",	--2673
		x"6c",	--2674
		x"70",	--2675
		x"6c",	--2676
		x"6a",	--2677
		x"6c",	--2678
		x"36",	--2679
		x"0e",	--2680
		x"32",	--2681
		x"1b",	--2682
		x"02",	--2683
		x"3b",	--2684
		x"82",	--2685
		x"6d",	--2686
		x"3b",	--2687
		x"80",	--2688
		x"5e",	--2689
		x"0c",	--2690
		x"0d",	--2691
		x"3c",	--2692
		x"7f",	--2693
		x"0d",	--2694
		x"3c",	--2695
		x"40",	--2696
		x"40",	--2697
		x"3e",	--2698
		x"3f",	--2699
		x"0f",	--2700
		x"0f",	--2701
		x"4a",	--2702
		x"0d",	--2703
		x"3d",	--2704
		x"7f",	--2705
		x"12",	--2706
		x"0f",	--2707
		x"0e",	--2708
		x"12",	--2709
		x"0f",	--2710
		x"0e",	--2711
		x"12",	--2712
		x"0f",	--2713
		x"0e",	--2714
		x"12",	--2715
		x"0f",	--2716
		x"0e",	--2717
		x"12",	--2718
		x"0f",	--2719
		x"0e",	--2720
		x"12",	--2721
		x"0f",	--2722
		x"0e",	--2723
		x"12",	--2724
		x"0f",	--2725
		x"0e",	--2726
		x"3e",	--2727
		x"3f",	--2728
		x"7f",	--2729
		x"4d",	--2730
		x"05",	--2731
		x"0f",	--2732
		x"cc",	--2733
		x"4d",	--2734
		x"0e",	--2735
		x"0f",	--2736
		x"4d",	--2737
		x"0d",	--2738
		x"0d",	--2739
		x"0d",	--2740
		x"0d",	--2741
		x"0d",	--2742
		x"0d",	--2743
		x"0d",	--2744
		x"0c",	--2745
		x"3c",	--2746
		x"7f",	--2747
		x"0c",	--2748
		x"4f",	--2749
		x"0f",	--2750
		x"0f",	--2751
		x"0f",	--2752
		x"0d",	--2753
		x"0d",	--2754
		x"0f",	--2755
		x"37",	--2756
		x"38",	--2757
		x"39",	--2758
		x"3a",	--2759
		x"3b",	--2760
		x"30",	--2761
		x"0d",	--2762
		x"be",	--2763
		x"0c",	--2764
		x"0d",	--2765
		x"3c",	--2766
		x"80",	--2767
		x"0d",	--2768
		x"0c",	--2769
		x"02",	--2770
		x"0d",	--2771
		x"b8",	--2772
		x"3e",	--2773
		x"40",	--2774
		x"0f",	--2775
		x"b4",	--2776
		x"12",	--2777
		x"0f",	--2778
		x"0e",	--2779
		x"0d",	--2780
		x"3d",	--2781
		x"80",	--2782
		x"b2",	--2783
		x"7d",	--2784
		x"0e",	--2785
		x"0f",	--2786
		x"cd",	--2787
		x"0e",	--2788
		x"3f",	--2789
		x"10",	--2790
		x"3e",	--2791
		x"3f",	--2792
		x"7f",	--2793
		x"7d",	--2794
		x"c5",	--2795
		x"37",	--2796
		x"82",	--2797
		x"07",	--2798
		x"37",	--2799
		x"1a",	--2800
		x"4f",	--2801
		x"0c",	--2802
		x"0d",	--2803
		x"4b",	--2804
		x"7b",	--2805
		x"1f",	--2806
		x"05",	--2807
		x"12",	--2808
		x"0d",	--2809
		x"0c",	--2810
		x"7b",	--2811
		x"fb",	--2812
		x"18",	--2813
		x"09",	--2814
		x"77",	--2815
		x"1f",	--2816
		x"04",	--2817
		x"08",	--2818
		x"09",	--2819
		x"77",	--2820
		x"fc",	--2821
		x"38",	--2822
		x"39",	--2823
		x"08",	--2824
		x"09",	--2825
		x"1e",	--2826
		x"0f",	--2827
		x"08",	--2828
		x"04",	--2829
		x"09",	--2830
		x"02",	--2831
		x"0e",	--2832
		x"0f",	--2833
		x"08",	--2834
		x"09",	--2835
		x"08",	--2836
		x"09",	--2837
		x"0e",	--2838
		x"0f",	--2839
		x"3e",	--2840
		x"7f",	--2841
		x"0f",	--2842
		x"3e",	--2843
		x"40",	--2844
		x"26",	--2845
		x"38",	--2846
		x"3f",	--2847
		x"09",	--2848
		x"0e",	--2849
		x"0f",	--2850
		x"12",	--2851
		x"0f",	--2852
		x"0e",	--2853
		x"12",	--2854
		x"0f",	--2855
		x"0e",	--2856
		x"12",	--2857
		x"0f",	--2858
		x"0e",	--2859
		x"12",	--2860
		x"0f",	--2861
		x"0e",	--2862
		x"12",	--2863
		x"0f",	--2864
		x"0e",	--2865
		x"12",	--2866
		x"0f",	--2867
		x"0e",	--2868
		x"12",	--2869
		x"0f",	--2870
		x"0e",	--2871
		x"3e",	--2872
		x"3f",	--2873
		x"7f",	--2874
		x"5d",	--2875
		x"39",	--2876
		x"00",	--2877
		x"72",	--2878
		x"4d",	--2879
		x"70",	--2880
		x"08",	--2881
		x"09",	--2882
		x"da",	--2883
		x"0f",	--2884
		x"d8",	--2885
		x"0e",	--2886
		x"0f",	--2887
		x"3e",	--2888
		x"80",	--2889
		x"0f",	--2890
		x"0e",	--2891
		x"04",	--2892
		x"38",	--2893
		x"40",	--2894
		x"09",	--2895
		x"d0",	--2896
		x"0f",	--2897
		x"ce",	--2898
		x"f9",	--2899
		x"0b",	--2900
		x"0a",	--2901
		x"2a",	--2902
		x"5b",	--2903
		x"02",	--2904
		x"3b",	--2905
		x"7f",	--2906
		x"1d",	--2907
		x"02",	--2908
		x"12",	--2909
		x"0d",	--2910
		x"12",	--2911
		x"0d",	--2912
		x"12",	--2913
		x"0d",	--2914
		x"12",	--2915
		x"0d",	--2916
		x"12",	--2917
		x"0d",	--2918
		x"12",	--2919
		x"0d",	--2920
		x"12",	--2921
		x"0d",	--2922
		x"4d",	--2923
		x"5f",	--2924
		x"03",	--2925
		x"3f",	--2926
		x"80",	--2927
		x"0f",	--2928
		x"0f",	--2929
		x"ce",	--2930
		x"01",	--2931
		x"0d",	--2932
		x"2d",	--2933
		x"0a",	--2934
		x"51",	--2935
		x"be",	--2936
		x"82",	--2937
		x"02",	--2938
		x"0c",	--2939
		x"0d",	--2940
		x"0c",	--2941
		x"0d",	--2942
		x"0c",	--2943
		x"0d",	--2944
		x"0c",	--2945
		x"0d",	--2946
		x"0c",	--2947
		x"0d",	--2948
		x"0c",	--2949
		x"0d",	--2950
		x"0c",	--2951
		x"0d",	--2952
		x"0c",	--2953
		x"0d",	--2954
		x"fe",	--2955
		x"03",	--2956
		x"00",	--2957
		x"3d",	--2958
		x"00",	--2959
		x"0b",	--2960
		x"3f",	--2961
		x"81",	--2962
		x"0c",	--2963
		x"0d",	--2964
		x"0a",	--2965
		x"3f",	--2966
		x"3d",	--2967
		x"00",	--2968
		x"f9",	--2969
		x"8e",	--2970
		x"02",	--2971
		x"8e",	--2972
		x"04",	--2973
		x"8e",	--2974
		x"06",	--2975
		x"3a",	--2976
		x"3b",	--2977
		x"30",	--2978
		x"3d",	--2979
		x"ff",	--2980
		x"2a",	--2981
		x"3d",	--2982
		x"81",	--2983
		x"8e",	--2984
		x"02",	--2985
		x"fe",	--2986
		x"03",	--2987
		x"00",	--2988
		x"0c",	--2989
		x"0d",	--2990
		x"0c",	--2991
		x"0d",	--2992
		x"0c",	--2993
		x"0d",	--2994
		x"0c",	--2995
		x"0d",	--2996
		x"0c",	--2997
		x"0d",	--2998
		x"0c",	--2999
		x"0d",	--3000
		x"0c",	--3001
		x"0d",	--3002
		x"0c",	--3003
		x"0d",	--3004
		x"0a",	--3005
		x"0b",	--3006
		x"0a",	--3007
		x"3b",	--3008
		x"00",	--3009
		x"8e",	--3010
		x"04",	--3011
		x"8e",	--3012
		x"06",	--3013
		x"3a",	--3014
		x"3b",	--3015
		x"30",	--3016
		x"0b",	--3017
		x"ad",	--3018
		x"ee",	--3019
		x"00",	--3020
		x"3a",	--3021
		x"3b",	--3022
		x"30",	--3023
		x"0a",	--3024
		x"0c",	--3025
		x"0c",	--3026
		x"0d",	--3027
		x"0c",	--3028
		x"3d",	--3029
		x"10",	--3030
		x"0c",	--3031
		x"02",	--3032
		x"0d",	--3033
		x"08",	--3034
		x"de",	--3035
		x"00",	--3036
		x"e4",	--3037
		x"0b",	--3038
		x"f2",	--3039
		x"ee",	--3040
		x"00",	--3041
		x"e3",	--3042
		x"ce",	--3043
		x"00",	--3044
		x"dc",	--3045
		x"0b",	--3046
		x"6d",	--3047
		x"6d",	--3048
		x"12",	--3049
		x"6c",	--3050
		x"6c",	--3051
		x"0f",	--3052
		x"6d",	--3053
		x"41",	--3054
		x"6c",	--3055
		x"11",	--3056
		x"6d",	--3057
		x"0d",	--3058
		x"6c",	--3059
		x"14",	--3060
		x"5d",	--3061
		x"01",	--3062
		x"5d",	--3063
		x"01",	--3064
		x"14",	--3065
		x"4d",	--3066
		x"09",	--3067
		x"1e",	--3068
		x"0f",	--3069
		x"3b",	--3070
		x"30",	--3071
		x"6c",	--3072
		x"28",	--3073
		x"ce",	--3074
		x"01",	--3075
		x"f7",	--3076
		x"3e",	--3077
		x"0f",	--3078
		x"3b",	--3079
		x"30",	--3080
		x"cf",	--3081
		x"01",	--3082
		x"f0",	--3083
		x"3e",	--3084
		x"f8",	--3085
		x"1b",	--3086
		x"02",	--3087
		x"1c",	--3088
		x"02",	--3089
		x"0c",	--3090
		x"e6",	--3091
		x"0b",	--3092
		x"16",	--3093
		x"1b",	--3094
		x"04",	--3095
		x"1f",	--3096
		x"06",	--3097
		x"1c",	--3098
		x"04",	--3099
		x"1e",	--3100
		x"06",	--3101
		x"0e",	--3102
		x"da",	--3103
		x"0f",	--3104
		x"02",	--3105
		x"0c",	--3106
		x"d6",	--3107
		x"0f",	--3108
		x"06",	--3109
		x"0e",	--3110
		x"02",	--3111
		x"0b",	--3112
		x"02",	--3113
		x"0e",	--3114
		x"d1",	--3115
		x"4d",	--3116
		x"ce",	--3117
		x"3e",	--3118
		x"d6",	--3119
		x"6c",	--3120
		x"d7",	--3121
		x"5e",	--3122
		x"01",	--3123
		x"5f",	--3124
		x"01",	--3125
		x"0e",	--3126
		x"c5",	--3127
		x"0d",	--3128
		x"0f",	--3129
		x"04",	--3130
		x"3d",	--3131
		x"03",	--3132
		x"3f",	--3133
		x"1f",	--3134
		x"0e",	--3135
		x"03",	--3136
		x"5d",	--3137
		x"3e",	--3138
		x"1e",	--3139
		x"0d",	--3140
		x"b0",	--3141
		x"f6",	--3142
		x"3d",	--3143
		x"6d",	--3144
		x"02",	--3145
		x"3e",	--3146
		x"1e",	--3147
		x"5d",	--3148
		x"02",	--3149
		x"3f",	--3150
		x"1f",	--3151
		x"30",	--3152
		x"b0",	--3153
		x"70",	--3154
		x"0f",	--3155
		x"30",	--3156
		x"0b",	--3157
		x"0b",	--3158
		x"0f",	--3159
		x"06",	--3160
		x"3b",	--3161
		x"03",	--3162
		x"3e",	--3163
		x"3f",	--3164
		x"1e",	--3165
		x"0f",	--3166
		x"0d",	--3167
		x"05",	--3168
		x"5b",	--3169
		x"3c",	--3170
		x"3d",	--3171
		x"1c",	--3172
		x"0d",	--3173
		x"b0",	--3174
		x"18",	--3175
		x"6b",	--3176
		x"04",	--3177
		x"3c",	--3178
		x"3d",	--3179
		x"1c",	--3180
		x"0d",	--3181
		x"5b",	--3182
		x"04",	--3183
		x"3e",	--3184
		x"3f",	--3185
		x"1e",	--3186
		x"0f",	--3187
		x"3b",	--3188
		x"30",	--3189
		x"b0",	--3190
		x"aa",	--3191
		x"0e",	--3192
		x"0f",	--3193
		x"30",	--3194
		x"7c",	--3195
		x"10",	--3196
		x"0d",	--3197
		x"0e",	--3198
		x"0f",	--3199
		x"0e",	--3200
		x"0e",	--3201
		x"02",	--3202
		x"0e",	--3203
		x"1f",	--3204
		x"1c",	--3205
		x"f8",	--3206
		x"30",	--3207
		x"b0",	--3208
		x"f6",	--3209
		x"0f",	--3210
		x"30",	--3211
		x"0b",	--3212
		x"0a",	--3213
		x"09",	--3214
		x"79",	--3215
		x"20",	--3216
		x"0a",	--3217
		x"0b",	--3218
		x"0c",	--3219
		x"0d",	--3220
		x"0e",	--3221
		x"0f",	--3222
		x"0c",	--3223
		x"0d",	--3224
		x"0d",	--3225
		x"06",	--3226
		x"02",	--3227
		x"0c",	--3228
		x"03",	--3229
		x"0c",	--3230
		x"0d",	--3231
		x"1e",	--3232
		x"19",	--3233
		x"f2",	--3234
		x"39",	--3235
		x"3a",	--3236
		x"3b",	--3237
		x"30",	--3238
		x"b0",	--3239
		x"18",	--3240
		x"0e",	--3241
		x"0f",	--3242
		x"30",	--3243
		x"00",	--3244
		x"32",	--3245
		x"f0",	--3246
		x"fd",	--3247
		x"57",	--3248
		x"69",	--3249
		x"69",	--3250
		x"67",	--3251
		x"66",	--3252
		x"72",	--3253
		x"61",	--3254
		x"6e",	--3255
		x"77",	--3256
		x"2e",	--3257
		x"69",	--3258
		x"20",	--3259
		x"69",	--3260
		x"65",	--3261
		x"0a",	--3262
		x"57",	--3263
		x"20",	--3264
		x"68",	--3265
		x"75",	--3266
		x"64",	--3267
		x"6e",	--3268
		x"74",	--3269
		x"73",	--3270
		x"65",	--3271
		x"74",	--3272
		x"61",	--3273
		x"0d",	--3274
		x"00",	--3275
		x"6f",	--3276
		x"72",	--3277
		x"63",	--3278
		x"20",	--3279
		x"73",	--3280
		x"67",	--3281
		x"3a",	--3282
		x"0a",	--3283
		x"09",	--3284
		x"63",	--3285
		x"4c",	--3286
		x"46",	--3287
		x"20",	--3288
		x"49",	--3289
		x"48",	--3290
		x"0d",	--3291
		x"00",	--3292
		x"6f",	--3293
		x"65",	--3294
		x"68",	--3295
		x"6e",	--3296
		x"20",	--3297
		x"65",	--3298
		x"74",	--3299
		x"74",	--3300
		x"72",	--3301
		x"69",	--3302
		x"6c",	--3303
		x"20",	--3304
		x"72",	--3305
		x"6e",	--3306
		x"0d",	--3307
		x"00",	--3308
		x"64",	--3309
		x"25",	--3310
		x"0d",	--3311
		x"00",	--3312
		x"0a",	--3313
		x"3d",	--3314
		x"3d",	--3315
		x"3d",	--3316
		x"4d",	--3317
		x"72",	--3318
		x"65",	--3319
		x"20",	--3320
		x"43",	--3321
		x"20",	--3322
		x"3d",	--3323
		x"3d",	--3324
		x"3d",	--3325
		x"0a",	--3326
		x"77",	--3327
		x"69",	--3328
		x"65",	--3329
		x"72",	--3330
		x"61",	--3331
		x"00",	--3332
		x"77",	--3333
		x"00",	--3334
		x"6e",	--3335
		x"6f",	--3336
		x"65",	--3337
		x"00",	--3338
		x"6f",	--3339
		x"74",	--3340
		x"6f",	--3341
		x"64",	--3342
		x"72",	--3343
		x"0d",	--3344
		x"00",	--3345
		x"20",	--3346
		x"00",	--3347
		x"63",	--3348
		x"77",	--3349
		x"69",	--3350
		x"65",	--3351
		x"0d",	--3352
		x"63",	--3353
		x"72",	--3354
		x"65",	--3355
		x"74",	--3356
		x"75",	--3357
		x"61",	--3358
		x"65",	--3359
		x"0d",	--3360
		x"00",	--3361
		x"25",	--3362
		x"20",	--3363
		x"45",	--3364
		x"49",	--3365
		x"54",	--3366
		x"52",	--3367
		x"56",	--3368
		x"4c",	--3369
		x"45",	--3370
		x"0a",	--3371
		x"53",	--3372
		x"6d",	--3373
		x"74",	--3374
		x"69",	--3375
		x"67",	--3376
		x"77",	--3377
		x"6e",	--3378
		x"20",	--3379
		x"65",	--3380
		x"72",	--3381
		x"62",	--3382
		x"79",	--3383
		x"77",	--3384
		x"6f",	--3385
		x"67",	--3386
		x"0a",	--3387
		x"72",	--3388
		x"25",	--3389
		x"20",	--3390
		x"3d",	--3391
		x"64",	--3392
		x"0a",	--3393
		x"72",	--3394
		x"61",	--3395
		x"0a",	--3396
		x"00",	--3397
		x"25",	--3398
		x"20",	--3399
		x"45",	--3400
		x"49",	--3401
		x"54",	--3402
		x"52",	--3403
		x"0a",	--3404
		x"25",	--3405
		x"20",	--3406
		x"73",	--3407
		x"6e",	--3408
		x"74",	--3409
		x"61",	--3410
		x"6e",	--3411
		x"6d",	--3412
		x"65",	--3413
		x"0d",	--3414
		x"00",	--3415
		x"63",	--3416
		x"25",	--3417
		x"0d",	--3418
		x"00",	--3419
		x"63",	--3420
		x"20",	--3421
		x"6f",	--3422
		x"73",	--3423
		x"63",	--3424
		x"20",	--3425
		x"6f",	--3426
		x"6d",	--3427
		x"6e",	--3428
		x"0d",	--3429
		x"00",	--3430
		x"00",	--3431
		x"2e",	--3432
		x"2e",	--3433
		x"2e",	--3434
		x"2e",	--3435
		x"2e",	--3436
		x"2e",	--3437
		x"2e",	--3438
		x"2e",	--3439
		x"2e",	--3440
		x"2e",	--3441
		x"2e",	--3442
		x"2e",	--3443
		x"2e",	--3444
		x"2e",	--3445
		x"2e",	--3446
		x"2e",	--3447
		x"2e",	--3448
		x"2e",	--3449
		x"2e",	--3450
		x"2e",	--3451
		x"2e",	--3452
		x"2e",	--3453
		x"2e",	--3454
		x"2e",	--3455
		x"2e",	--3456
		x"2e",	--3457
		x"2e",	--3458
		x"2e",	--3459
		x"f2",	--3460
		x"2e",	--3461
		x"2e",	--3462
		x"2e",	--3463
		x"2e",	--3464
		x"2e",	--3465
		x"2e",	--3466
		x"2e",	--3467
		x"2e",	--3468
		x"2e",	--3469
		x"2e",	--3470
		x"2e",	--3471
		x"2e",	--3472
		x"2e",	--3473
		x"2e",	--3474
		x"2e",	--3475
		x"2e",	--3476
		x"2e",	--3477
		x"2e",	--3478
		x"2e",	--3479
		x"2e",	--3480
		x"2e",	--3481
		x"2e",	--3482
		x"2e",	--3483
		x"2e",	--3484
		x"2e",	--3485
		x"2e",	--3486
		x"2e",	--3487
		x"2e",	--3488
		x"2e",	--3489
		x"2e",	--3490
		x"2e",	--3491
		x"e4",	--3492
		x"d6",	--3493
		x"c8",	--3494
		x"2e",	--3495
		x"2e",	--3496
		x"2e",	--3497
		x"2e",	--3498
		x"2e",	--3499
		x"2e",	--3500
		x"2e",	--3501
		x"b0",	--3502
		x"2e",	--3503
		x"9e",	--3504
		x"2e",	--3505
		x"2e",	--3506
		x"2e",	--3507
		x"2e",	--3508
		x"82",	--3509
		x"2e",	--3510
		x"2e",	--3511
		x"2e",	--3512
		x"74",	--3513
		x"62",	--3514
		x"30",	--3515
		x"32",	--3516
		x"34",	--3517
		x"36",	--3518
		x"38",	--3519
		x"61",	--3520
		x"63",	--3521
		x"65",	--3522
		x"00",	--3523
		x"00",	--3524
		x"00",	--3525
		x"00",	--3526
		x"00",	--3527
		x"00",	--3528
		x"02",	--3529
		x"03",	--3530
		x"03",	--3531
		x"04",	--3532
		x"04",	--3533
		x"04",	--3534
		x"04",	--3535
		x"05",	--3536
		x"05",	--3537
		x"05",	--3538
		x"05",	--3539
		x"05",	--3540
		x"05",	--3541
		x"05",	--3542
		x"05",	--3543
		x"06",	--3544
		x"06",	--3545
		x"06",	--3546
		x"06",	--3547
		x"06",	--3548
		x"06",	--3549
		x"06",	--3550
		x"06",	--3551
		x"06",	--3552
		x"06",	--3553
		x"06",	--3554
		x"06",	--3555
		x"06",	--3556
		x"06",	--3557
		x"06",	--3558
		x"06",	--3559
		x"07",	--3560
		x"07",	--3561
		x"07",	--3562
		x"07",	--3563
		x"07",	--3564
		x"07",	--3565
		x"07",	--3566
		x"07",	--3567
		x"07",	--3568
		x"07",	--3569
		x"07",	--3570
		x"07",	--3571
		x"07",	--3572
		x"07",	--3573
		x"07",	--3574
		x"07",	--3575
		x"07",	--3576
		x"07",	--3577
		x"07",	--3578
		x"07",	--3579
		x"07",	--3580
		x"07",	--3581
		x"07",	--3582
		x"07",	--3583
		x"07",	--3584
		x"07",	--3585
		x"07",	--3586
		x"07",	--3587
		x"07",	--3588
		x"07",	--3589
		x"07",	--3590
		x"07",	--3591
		x"08",	--3592
		x"08",	--3593
		x"08",	--3594
		x"08",	--3595
		x"08",	--3596
		x"08",	--3597
		x"08",	--3598
		x"08",	--3599
		x"08",	--3600
		x"08",	--3601
		x"08",	--3602
		x"08",	--3603
		x"08",	--3604
		x"08",	--3605
		x"08",	--3606
		x"08",	--3607
		x"08",	--3608
		x"08",	--3609
		x"08",	--3610
		x"08",	--3611
		x"08",	--3612
		x"08",	--3613
		x"08",	--3614
		x"08",	--3615
		x"08",	--3616
		x"08",	--3617
		x"08",	--3618
		x"08",	--3619
		x"08",	--3620
		x"08",	--3621
		x"08",	--3622
		x"08",	--3623
		x"08",	--3624
		x"08",	--3625
		x"08",	--3626
		x"08",	--3627
		x"08",	--3628
		x"08",	--3629
		x"08",	--3630
		x"08",	--3631
		x"08",	--3632
		x"08",	--3633
		x"08",	--3634
		x"08",	--3635
		x"08",	--3636
		x"08",	--3637
		x"08",	--3638
		x"08",	--3639
		x"08",	--3640
		x"08",	--3641
		x"08",	--3642
		x"08",	--3643
		x"08",	--3644
		x"08",	--3645
		x"08",	--3646
		x"08",	--3647
		x"08",	--3648
		x"08",	--3649
		x"08",	--3650
		x"08",	--3651
		x"08",	--3652
		x"08",	--3653
		x"08",	--3654
		x"08",	--3655
		x"68",	--3656
		x"6c",	--3657
		x"00",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"ba",	--4080
		x"ba",	--4081
		x"ba",	--4082
		x"ba",	--4083
		x"ba",	--4084
		x"ba",	--4085
		x"ba",	--4086
		x"0a",	--4087
		x"c2",	--4088
		x"ba",	--4089
		x"ba",	--4090
		x"ba",	--4091
		x"ba",	--4092
		x"ba",	--4093
		x"ba",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"04",	--5
		x"40",	--6
		x"06",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"04",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fc",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"02",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"04",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"25",	--41
		x"43",	--42
		x"12",	--43
		x"eb",	--44
		x"12",	--45
		x"e6",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"f9",	--50
		x"12",	--51
		x"ea",	--52
		x"53",	--53
		x"40",	--54
		x"f9",	--55
		x"40",	--56
		x"e3",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"e6",	--61
		x"40",	--62
		x"fa",	--63
		x"40",	--64
		x"e3",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"e6",	--69
		x"40",	--70
		x"fa",	--71
		x"40",	--72
		x"e1",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"e6",	--77
		x"40",	--78
		x"fa",	--79
		x"40",	--80
		x"e2",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"e6",	--85
		x"40",	--86
		x"fa",	--87
		x"40",	--88
		x"e1",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"e6",	--93
		x"43",	--94
		x"12",	--95
		x"e6",	--96
		x"43",	--97
		x"40",	--98
		x"4e",	--99
		x"40",	--100
		x"01",	--101
		x"41",	--102
		x"50",	--103
		x"00",	--104
		x"12",	--105
		x"e5",	--106
		x"41",	--107
		x"50",	--108
		x"00",	--109
		x"12",	--110
		x"e5",	--111
		x"43",	--112
		x"40",	--113
		x"4e",	--114
		x"40",	--115
		x"01",	--116
		x"41",	--117
		x"52",	--118
		x"12",	--119
		x"e5",	--120
		x"41",	--121
		x"52",	--122
		x"12",	--123
		x"e5",	--124
		x"41",	--125
		x"52",	--126
		x"41",	--127
		x"50",	--128
		x"00",	--129
		x"12",	--130
		x"e1",	--131
		x"40",	--132
		x"01",	--133
		x"41",	--134
		x"53",	--135
		x"12",	--136
		x"e8",	--137
		x"40",	--138
		x"01",	--139
		x"41",	--140
		x"12",	--141
		x"e8",	--142
		x"41",	--143
		x"41",	--144
		x"53",	--145
		x"12",	--146
		x"e2",	--147
		x"12",	--148
		x"e7",	--149
		x"43",	--150
		x"40",	--151
		x"e2",	--152
		x"40",	--153
		x"01",	--154
		x"12",	--155
		x"e7",	--156
		x"12",	--157
		x"e7",	--158
		x"40",	--159
		x"ff",	--160
		x"00",	--161
		x"d2",	--162
		x"43",	--163
		x"12",	--164
		x"eb",	--165
		x"93",	--166
		x"27",	--167
		x"12",	--168
		x"eb",	--169
		x"92",	--170
		x"24",	--171
		x"90",	--172
		x"00",	--173
		x"20",	--174
		x"12",	--175
		x"fa",	--176
		x"12",	--177
		x"ea",	--178
		x"53",	--179
		x"41",	--180
		x"50",	--181
		x"00",	--182
		x"41",	--183
		x"00",	--184
		x"12",	--185
		x"e6",	--186
		x"43",	--187
		x"3f",	--188
		x"93",	--189
		x"27",	--190
		x"53",	--191
		x"12",	--192
		x"fa",	--193
		x"12",	--194
		x"ea",	--195
		x"53",	--196
		x"3f",	--197
		x"90",	--198
		x"00",	--199
		x"2f",	--200
		x"4f",	--201
		x"11",	--202
		x"12",	--203
		x"12",	--204
		x"fa",	--205
		x"4f",	--206
		x"00",	--207
		x"12",	--208
		x"ea",	--209
		x"52",	--210
		x"40",	--211
		x"00",	--212
		x"51",	--213
		x"5b",	--214
		x"41",	--215
		x"00",	--216
		x"4f",	--217
		x"00",	--218
		x"53",	--219
		x"3f",	--220
		x"40",	--221
		x"f9",	--222
		x"40",	--223
		x"e0",	--224
		x"01",	--225
		x"42",	--226
		x"01",	--227
		x"40",	--228
		x"02",	--229
		x"01",	--230
		x"12",	--231
		x"f9",	--232
		x"12",	--233
		x"ea",	--234
		x"43",	--235
		x"01",	--236
		x"40",	--237
		x"f9",	--238
		x"00",	--239
		x"12",	--240
		x"ea",	--241
		x"53",	--242
		x"43",	--243
		x"41",	--244
		x"4f",	--245
		x"02",	--246
		x"4e",	--247
		x"02",	--248
		x"41",	--249
		x"82",	--250
		x"90",	--251
		x"00",	--252
		x"00",	--253
		x"20",	--254
		x"93",	--255
		x"00",	--256
		x"24",	--257
		x"41",	--258
		x"4f",	--259
		x"53",	--260
		x"41",	--261
		x"52",	--262
		x"12",	--263
		x"e4",	--264
		x"93",	--265
		x"00",	--266
		x"24",	--267
		x"41",	--268
		x"4f",	--269
		x"41",	--270
		x"53",	--271
		x"12",	--272
		x"e4",	--273
		x"93",	--274
		x"00",	--275
		x"24",	--276
		x"41",	--277
		x"00",	--278
		x"43",	--279
		x"12",	--280
		x"f3",	--281
		x"43",	--282
		x"40",	--283
		x"42",	--284
		x"12",	--285
		x"f1",	--286
		x"4e",	--287
		x"4f",	--288
		x"42",	--289
		x"02",	--290
		x"12",	--291
		x"e6",	--292
		x"41",	--293
		x"00",	--294
		x"43",	--295
		x"12",	--296
		x"f3",	--297
		x"43",	--298
		x"40",	--299
		x"42",	--300
		x"12",	--301
		x"f1",	--302
		x"4e",	--303
		x"4f",	--304
		x"42",	--305
		x"02",	--306
		x"12",	--307
		x"e6",	--308
		x"43",	--309
		x"52",	--310
		x"41",	--311
		x"12",	--312
		x"f9",	--313
		x"4f",	--314
		x"00",	--315
		x"12",	--316
		x"ea",	--317
		x"41",	--318
		x"00",	--319
		x"4f",	--320
		x"11",	--321
		x"4f",	--322
		x"00",	--323
		x"12",	--324
		x"f9",	--325
		x"12",	--326
		x"ea",	--327
		x"52",	--328
		x"43",	--329
		x"52",	--330
		x"41",	--331
		x"12",	--332
		x"f9",	--333
		x"12",	--334
		x"ea",	--335
		x"53",	--336
		x"43",	--337
		x"3f",	--338
		x"4f",	--339
		x"02",	--340
		x"4e",	--341
		x"02",	--342
		x"41",	--343
		x"12",	--344
		x"01",	--345
		x"12",	--346
		x"01",	--347
		x"12",	--348
		x"f9",	--349
		x"12",	--350
		x"ea",	--351
		x"50",	--352
		x"00",	--353
		x"43",	--354
		x"41",	--355
		x"42",	--356
		x"02",	--357
		x"93",	--358
		x"24",	--359
		x"93",	--360
		x"38",	--361
		x"24",	--362
		x"90",	--363
		x"00",	--364
		x"24",	--365
		x"90",	--366
		x"00",	--367
		x"38",	--368
		x"43",	--369
		x"02",	--370
		x"41",	--371
		x"40",	--372
		x"00",	--373
		x"00",	--374
		x"53",	--375
		x"4f",	--376
		x"02",	--377
		x"41",	--378
		x"42",	--379
		x"00",	--380
		x"43",	--381
		x"02",	--382
		x"41",	--383
		x"42",	--384
		x"00",	--385
		x"53",	--386
		x"4f",	--387
		x"02",	--388
		x"41",	--389
		x"93",	--390
		x"23",	--391
		x"43",	--392
		x"00",	--393
		x"53",	--394
		x"4f",	--395
		x"02",	--396
		x"41",	--397
		x"42",	--398
		x"00",	--399
		x"4e",	--400
		x"be",	--401
		x"20",	--402
		x"df",	--403
		x"00",	--404
		x"41",	--405
		x"cf",	--406
		x"00",	--407
		x"41",	--408
		x"12",	--409
		x"50",	--410
		x"ff",	--411
		x"4f",	--412
		x"12",	--413
		x"fa",	--414
		x"12",	--415
		x"ea",	--416
		x"53",	--417
		x"90",	--418
		x"00",	--419
		x"00",	--420
		x"20",	--421
		x"93",	--422
		x"00",	--423
		x"24",	--424
		x"41",	--425
		x"4b",	--426
		x"53",	--427
		x"41",	--428
		x"52",	--429
		x"12",	--430
		x"e4",	--431
		x"93",	--432
		x"00",	--433
		x"24",	--434
		x"41",	--435
		x"4f",	--436
		x"41",	--437
		x"53",	--438
		x"12",	--439
		x"e4",	--440
		x"93",	--441
		x"00",	--442
		x"24",	--443
		x"12",	--444
		x"00",	--445
		x"12",	--446
		x"00",	--447
		x"12",	--448
		x"fa",	--449
		x"12",	--450
		x"ea",	--451
		x"50",	--452
		x"00",	--453
		x"41",	--454
		x"00",	--455
		x"41",	--456
		x"00",	--457
		x"00",	--458
		x"43",	--459
		x"50",	--460
		x"00",	--461
		x"41",	--462
		x"41",	--463
		x"12",	--464
		x"fa",	--465
		x"12",	--466
		x"ea",	--467
		x"4b",	--468
		x"11",	--469
		x"4f",	--470
		x"00",	--471
		x"12",	--472
		x"fa",	--473
		x"12",	--474
		x"ea",	--475
		x"52",	--476
		x"43",	--477
		x"50",	--478
		x"00",	--479
		x"41",	--480
		x"41",	--481
		x"12",	--482
		x"fa",	--483
		x"12",	--484
		x"ea",	--485
		x"53",	--486
		x"43",	--487
		x"3f",	--488
		x"12",	--489
		x"82",	--490
		x"4f",	--491
		x"12",	--492
		x"fa",	--493
		x"12",	--494
		x"ea",	--495
		x"53",	--496
		x"90",	--497
		x"00",	--498
		x"00",	--499
		x"20",	--500
		x"93",	--501
		x"00",	--502
		x"24",	--503
		x"41",	--504
		x"4b",	--505
		x"53",	--506
		x"41",	--507
		x"53",	--508
		x"12",	--509
		x"e4",	--510
		x"93",	--511
		x"00",	--512
		x"24",	--513
		x"41",	--514
		x"00",	--515
		x"12",	--516
		x"12",	--517
		x"12",	--518
		x"fa",	--519
		x"12",	--520
		x"ea",	--521
		x"50",	--522
		x"00",	--523
		x"43",	--524
		x"52",	--525
		x"41",	--526
		x"41",	--527
		x"12",	--528
		x"fa",	--529
		x"12",	--530
		x"ea",	--531
		x"4b",	--532
		x"11",	--533
		x"4f",	--534
		x"00",	--535
		x"12",	--536
		x"fa",	--537
		x"12",	--538
		x"ea",	--539
		x"52",	--540
		x"43",	--541
		x"52",	--542
		x"41",	--543
		x"41",	--544
		x"12",	--545
		x"fa",	--546
		x"12",	--547
		x"ea",	--548
		x"53",	--549
		x"43",	--550
		x"3f",	--551
		x"12",	--552
		x"12",	--553
		x"12",	--554
		x"12",	--555
		x"12",	--556
		x"43",	--557
		x"00",	--558
		x"43",	--559
		x"00",	--560
		x"4e",	--561
		x"93",	--562
		x"24",	--563
		x"4e",	--564
		x"53",	--565
		x"4e",	--566
		x"43",	--567
		x"43",	--568
		x"43",	--569
		x"3c",	--570
		x"90",	--571
		x"00",	--572
		x"2c",	--573
		x"4f",	--574
		x"5c",	--575
		x"5c",	--576
		x"5c",	--577
		x"5c",	--578
		x"4c",	--579
		x"00",	--580
		x"50",	--581
		x"ff",	--582
		x"48",	--583
		x"11",	--584
		x"5a",	--585
		x"4c",	--586
		x"00",	--587
		x"43",	--588
		x"53",	--589
		x"49",	--590
		x"4b",	--591
		x"4b",	--592
		x"93",	--593
		x"24",	--594
		x"90",	--595
		x"00",	--596
		x"24",	--597
		x"90",	--598
		x"00",	--599
		x"24",	--600
		x"4c",	--601
		x"50",	--602
		x"ff",	--603
		x"93",	--604
		x"23",	--605
		x"90",	--606
		x"00",	--607
		x"2c",	--608
		x"4f",	--609
		x"5a",	--610
		x"4a",	--611
		x"5c",	--612
		x"5c",	--613
		x"5a",	--614
		x"4c",	--615
		x"00",	--616
		x"50",	--617
		x"ff",	--618
		x"48",	--619
		x"11",	--620
		x"58",	--621
		x"4c",	--622
		x"00",	--623
		x"3f",	--624
		x"43",	--625
		x"3f",	--626
		x"4c",	--627
		x"50",	--628
		x"ff",	--629
		x"90",	--630
		x"00",	--631
		x"2c",	--632
		x"4f",	--633
		x"5c",	--634
		x"5c",	--635
		x"5c",	--636
		x"5c",	--637
		x"4c",	--638
		x"00",	--639
		x"50",	--640
		x"ff",	--641
		x"3f",	--642
		x"4c",	--643
		x"50",	--644
		x"ff",	--645
		x"90",	--646
		x"00",	--647
		x"2c",	--648
		x"4f",	--649
		x"5c",	--650
		x"5c",	--651
		x"5c",	--652
		x"5c",	--653
		x"4c",	--654
		x"00",	--655
		x"50",	--656
		x"ff",	--657
		x"3f",	--658
		x"43",	--659
		x"00",	--660
		x"43",	--661
		x"41",	--662
		x"41",	--663
		x"41",	--664
		x"41",	--665
		x"41",	--666
		x"41",	--667
		x"43",	--668
		x"00",	--669
		x"4a",	--670
		x"53",	--671
		x"5e",	--672
		x"41",	--673
		x"41",	--674
		x"41",	--675
		x"41",	--676
		x"41",	--677
		x"41",	--678
		x"11",	--679
		x"12",	--680
		x"12",	--681
		x"fa",	--682
		x"12",	--683
		x"ea",	--684
		x"52",	--685
		x"43",	--686
		x"41",	--687
		x"41",	--688
		x"41",	--689
		x"41",	--690
		x"41",	--691
		x"41",	--692
		x"12",	--693
		x"12",	--694
		x"4e",	--695
		x"4c",	--696
		x"4e",	--697
		x"00",	--698
		x"4d",	--699
		x"00",	--700
		x"4c",	--701
		x"00",	--702
		x"4d",	--703
		x"43",	--704
		x"40",	--705
		x"36",	--706
		x"40",	--707
		x"01",	--708
		x"12",	--709
		x"f8",	--710
		x"4e",	--711
		x"00",	--712
		x"12",	--713
		x"c2",	--714
		x"43",	--715
		x"4a",	--716
		x"01",	--717
		x"40",	--718
		x"00",	--719
		x"01",	--720
		x"42",	--721
		x"01",	--722
		x"00",	--723
		x"41",	--724
		x"43",	--725
		x"41",	--726
		x"41",	--727
		x"41",	--728
		x"12",	--729
		x"12",	--730
		x"12",	--731
		x"43",	--732
		x"00",	--733
		x"40",	--734
		x"3f",	--735
		x"00",	--736
		x"4f",	--737
		x"4b",	--738
		x"00",	--739
		x"43",	--740
		x"12",	--741
		x"f3",	--742
		x"43",	--743
		x"40",	--744
		x"3f",	--745
		x"12",	--746
		x"ef",	--747
		x"4e",	--748
		x"4f",	--749
		x"4b",	--750
		x"00",	--751
		x"43",	--752
		x"12",	--753
		x"f3",	--754
		x"4e",	--755
		x"4f",	--756
		x"48",	--757
		x"49",	--758
		x"12",	--759
		x"ee",	--760
		x"12",	--761
		x"eb",	--762
		x"4e",	--763
		x"00",	--764
		x"43",	--765
		x"00",	--766
		x"41",	--767
		x"41",	--768
		x"41",	--769
		x"41",	--770
		x"12",	--771
		x"12",	--772
		x"12",	--773
		x"4d",	--774
		x"4e",	--775
		x"4d",	--776
		x"00",	--777
		x"4e",	--778
		x"00",	--779
		x"4f",	--780
		x"49",	--781
		x"00",	--782
		x"43",	--783
		x"12",	--784
		x"f3",	--785
		x"4e",	--786
		x"4f",	--787
		x"4a",	--788
		x"4b",	--789
		x"12",	--790
		x"ef",	--791
		x"4e",	--792
		x"4f",	--793
		x"49",	--794
		x"00",	--795
		x"43",	--796
		x"12",	--797
		x"f3",	--798
		x"4e",	--799
		x"4f",	--800
		x"4a",	--801
		x"4b",	--802
		x"12",	--803
		x"ee",	--804
		x"12",	--805
		x"eb",	--806
		x"4e",	--807
		x"00",	--808
		x"41",	--809
		x"41",	--810
		x"41",	--811
		x"41",	--812
		x"12",	--813
		x"12",	--814
		x"93",	--815
		x"02",	--816
		x"38",	--817
		x"40",	--818
		x"02",	--819
		x"43",	--820
		x"12",	--821
		x"4b",	--822
		x"ff",	--823
		x"11",	--824
		x"12",	--825
		x"12",	--826
		x"fa",	--827
		x"12",	--828
		x"ea",	--829
		x"50",	--830
		x"00",	--831
		x"53",	--832
		x"50",	--833
		x"00",	--834
		x"92",	--835
		x"02",	--836
		x"3b",	--837
		x"43",	--838
		x"41",	--839
		x"41",	--840
		x"41",	--841
		x"42",	--842
		x"02",	--843
		x"90",	--844
		x"00",	--845
		x"34",	--846
		x"4e",	--847
		x"5f",	--848
		x"5e",	--849
		x"5f",	--850
		x"50",	--851
		x"02",	--852
		x"40",	--853
		x"00",	--854
		x"00",	--855
		x"40",	--856
		x"e6",	--857
		x"00",	--858
		x"40",	--859
		x"02",	--860
		x"00",	--861
		x"53",	--862
		x"4e",	--863
		x"02",	--864
		x"41",	--865
		x"12",	--866
		x"42",	--867
		x"02",	--868
		x"90",	--869
		x"00",	--870
		x"34",	--871
		x"4b",	--872
		x"5c",	--873
		x"5b",	--874
		x"5c",	--875
		x"50",	--876
		x"02",	--877
		x"4f",	--878
		x"00",	--879
		x"4e",	--880
		x"00",	--881
		x"4d",	--882
		x"00",	--883
		x"53",	--884
		x"4b",	--885
		x"02",	--886
		x"43",	--887
		x"41",	--888
		x"41",	--889
		x"43",	--890
		x"3f",	--891
		x"12",	--892
		x"42",	--893
		x"02",	--894
		x"93",	--895
		x"38",	--896
		x"92",	--897
		x"02",	--898
		x"24",	--899
		x"40",	--900
		x"02",	--901
		x"43",	--902
		x"3c",	--903
		x"50",	--904
		x"00",	--905
		x"9f",	--906
		x"ff",	--907
		x"24",	--908
		x"53",	--909
		x"9b",	--910
		x"23",	--911
		x"12",	--912
		x"fa",	--913
		x"12",	--914
		x"ea",	--915
		x"53",	--916
		x"43",	--917
		x"41",	--918
		x"41",	--919
		x"43",	--920
		x"4c",	--921
		x"5d",	--922
		x"5d",	--923
		x"5c",	--924
		x"50",	--925
		x"02",	--926
		x"4e",	--927
		x"12",	--928
		x"00",	--929
		x"41",	--930
		x"41",	--931
		x"d0",	--932
		x"02",	--933
		x"01",	--934
		x"40",	--935
		x"0b",	--936
		x"01",	--937
		x"43",	--938
		x"41",	--939
		x"12",	--940
		x"12",	--941
		x"4f",	--942
		x"42",	--943
		x"02",	--944
		x"90",	--945
		x"00",	--946
		x"34",	--947
		x"4f",	--948
		x"5b",	--949
		x"4b",	--950
		x"5c",	--951
		x"5c",	--952
		x"5b",	--953
		x"50",	--954
		x"02",	--955
		x"43",	--956
		x"00",	--957
		x"43",	--958
		x"00",	--959
		x"4a",	--960
		x"00",	--961
		x"4e",	--962
		x"00",	--963
		x"4d",	--964
		x"00",	--965
		x"4f",	--966
		x"53",	--967
		x"4e",	--968
		x"02",	--969
		x"41",	--970
		x"41",	--971
		x"41",	--972
		x"43",	--973
		x"3f",	--974
		x"5f",	--975
		x"4f",	--976
		x"5e",	--977
		x"5e",	--978
		x"5f",	--979
		x"43",	--980
		x"02",	--981
		x"43",	--982
		x"41",	--983
		x"5f",	--984
		x"4f",	--985
		x"5e",	--986
		x"5e",	--987
		x"5f",	--988
		x"43",	--989
		x"02",	--990
		x"43",	--991
		x"41",	--992
		x"12",	--993
		x"12",	--994
		x"12",	--995
		x"12",	--996
		x"12",	--997
		x"12",	--998
		x"93",	--999
		x"02",	--1000
		x"38",	--1001
		x"40",	--1002
		x"02",	--1003
		x"43",	--1004
		x"3c",	--1005
		x"53",	--1006
		x"4f",	--1007
		x"00",	--1008
		x"53",	--1009
		x"50",	--1010
		x"00",	--1011
		x"92",	--1012
		x"02",	--1013
		x"34",	--1014
		x"93",	--1015
		x"ff",	--1016
		x"27",	--1017
		x"4b",	--1018
		x"9b",	--1019
		x"00",	--1020
		x"2b",	--1021
		x"43",	--1022
		x"00",	--1023
		x"4b",	--1024
		x"00",	--1025
		x"12",	--1026
		x"00",	--1027
		x"53",	--1028
		x"50",	--1029
		x"00",	--1030
		x"92",	--1031
		x"02",	--1032
		x"3b",	--1033
		x"f0",	--1034
		x"ff",	--1035
		x"01",	--1036
		x"41",	--1037
		x"41",	--1038
		x"41",	--1039
		x"41",	--1040
		x"41",	--1041
		x"41",	--1042
		x"13",	--1043
		x"4e",	--1044
		x"00",	--1045
		x"43",	--1046
		x"41",	--1047
		x"4f",	--1048
		x"4f",	--1049
		x"41",	--1050
		x"42",	--1051
		x"00",	--1052
		x"f2",	--1053
		x"23",	--1054
		x"4f",	--1055
		x"00",	--1056
		x"43",	--1057
		x"41",	--1058
		x"f0",	--1059
		x"00",	--1060
		x"4f",	--1061
		x"fb",	--1062
		x"11",	--1063
		x"12",	--1064
		x"e8",	--1065
		x"41",	--1066
		x"12",	--1067
		x"4f",	--1068
		x"4f",	--1069
		x"11",	--1070
		x"11",	--1071
		x"11",	--1072
		x"11",	--1073
		x"4e",	--1074
		x"12",	--1075
		x"e8",	--1076
		x"4b",	--1077
		x"12",	--1078
		x"e8",	--1079
		x"41",	--1080
		x"41",	--1081
		x"12",	--1082
		x"12",	--1083
		x"4f",	--1084
		x"40",	--1085
		x"00",	--1086
		x"4a",	--1087
		x"4b",	--1088
		x"f0",	--1089
		x"00",	--1090
		x"24",	--1091
		x"11",	--1092
		x"53",	--1093
		x"23",	--1094
		x"f3",	--1095
		x"24",	--1096
		x"40",	--1097
		x"00",	--1098
		x"12",	--1099
		x"e8",	--1100
		x"53",	--1101
		x"93",	--1102
		x"23",	--1103
		x"41",	--1104
		x"41",	--1105
		x"41",	--1106
		x"40",	--1107
		x"00",	--1108
		x"3f",	--1109
		x"12",	--1110
		x"4f",	--1111
		x"4f",	--1112
		x"10",	--1113
		x"11",	--1114
		x"4e",	--1115
		x"12",	--1116
		x"e8",	--1117
		x"4b",	--1118
		x"12",	--1119
		x"e8",	--1120
		x"41",	--1121
		x"41",	--1122
		x"12",	--1123
		x"12",	--1124
		x"4e",	--1125
		x"4f",	--1126
		x"4f",	--1127
		x"10",	--1128
		x"11",	--1129
		x"4d",	--1130
		x"12",	--1131
		x"e8",	--1132
		x"4b",	--1133
		x"12",	--1134
		x"e8",	--1135
		x"4b",	--1136
		x"4a",	--1137
		x"10",	--1138
		x"10",	--1139
		x"ec",	--1140
		x"ec",	--1141
		x"4d",	--1142
		x"12",	--1143
		x"e8",	--1144
		x"4a",	--1145
		x"12",	--1146
		x"e8",	--1147
		x"41",	--1148
		x"41",	--1149
		x"41",	--1150
		x"12",	--1151
		x"12",	--1152
		x"12",	--1153
		x"4f",	--1154
		x"93",	--1155
		x"24",	--1156
		x"4e",	--1157
		x"53",	--1158
		x"43",	--1159
		x"4a",	--1160
		x"5b",	--1161
		x"4d",	--1162
		x"11",	--1163
		x"12",	--1164
		x"e8",	--1165
		x"99",	--1166
		x"24",	--1167
		x"53",	--1168
		x"b0",	--1169
		x"00",	--1170
		x"20",	--1171
		x"40",	--1172
		x"00",	--1173
		x"12",	--1174
		x"e8",	--1175
		x"3f",	--1176
		x"40",	--1177
		x"00",	--1178
		x"12",	--1179
		x"e8",	--1180
		x"3f",	--1181
		x"41",	--1182
		x"41",	--1183
		x"41",	--1184
		x"41",	--1185
		x"12",	--1186
		x"12",	--1187
		x"12",	--1188
		x"4f",	--1189
		x"93",	--1190
		x"24",	--1191
		x"4e",	--1192
		x"53",	--1193
		x"43",	--1194
		x"4a",	--1195
		x"11",	--1196
		x"12",	--1197
		x"e8",	--1198
		x"99",	--1199
		x"24",	--1200
		x"53",	--1201
		x"b0",	--1202
		x"00",	--1203
		x"23",	--1204
		x"40",	--1205
		x"00",	--1206
		x"12",	--1207
		x"e8",	--1208
		x"4a",	--1209
		x"11",	--1210
		x"12",	--1211
		x"e8",	--1212
		x"99",	--1213
		x"23",	--1214
		x"41",	--1215
		x"41",	--1216
		x"41",	--1217
		x"41",	--1218
		x"12",	--1219
		x"12",	--1220
		x"12",	--1221
		x"50",	--1222
		x"ff",	--1223
		x"4f",	--1224
		x"93",	--1225
		x"38",	--1226
		x"90",	--1227
		x"00",	--1228
		x"38",	--1229
		x"43",	--1230
		x"41",	--1231
		x"59",	--1232
		x"40",	--1233
		x"00",	--1234
		x"4b",	--1235
		x"12",	--1236
		x"f8",	--1237
		x"50",	--1238
		x"00",	--1239
		x"4f",	--1240
		x"00",	--1241
		x"53",	--1242
		x"40",	--1243
		x"00",	--1244
		x"4b",	--1245
		x"12",	--1246
		x"f8",	--1247
		x"4f",	--1248
		x"90",	--1249
		x"00",	--1250
		x"37",	--1251
		x"49",	--1252
		x"53",	--1253
		x"51",	--1254
		x"40",	--1255
		x"00",	--1256
		x"4b",	--1257
		x"12",	--1258
		x"f8",	--1259
		x"50",	--1260
		x"00",	--1261
		x"4f",	--1262
		x"00",	--1263
		x"53",	--1264
		x"41",	--1265
		x"5a",	--1266
		x"4f",	--1267
		x"11",	--1268
		x"12",	--1269
		x"e8",	--1270
		x"93",	--1271
		x"23",	--1272
		x"50",	--1273
		x"00",	--1274
		x"41",	--1275
		x"41",	--1276
		x"41",	--1277
		x"41",	--1278
		x"40",	--1279
		x"00",	--1280
		x"12",	--1281
		x"e8",	--1282
		x"e3",	--1283
		x"53",	--1284
		x"3f",	--1285
		x"43",	--1286
		x"43",	--1287
		x"3f",	--1288
		x"12",	--1289
		x"12",	--1290
		x"12",	--1291
		x"41",	--1292
		x"52",	--1293
		x"4b",	--1294
		x"49",	--1295
		x"93",	--1296
		x"20",	--1297
		x"3c",	--1298
		x"11",	--1299
		x"12",	--1300
		x"e8",	--1301
		x"49",	--1302
		x"4a",	--1303
		x"53",	--1304
		x"4a",	--1305
		x"00",	--1306
		x"93",	--1307
		x"24",	--1308
		x"90",	--1309
		x"00",	--1310
		x"23",	--1311
		x"49",	--1312
		x"53",	--1313
		x"49",	--1314
		x"00",	--1315
		x"50",	--1316
		x"ff",	--1317
		x"90",	--1318
		x"00",	--1319
		x"2f",	--1320
		x"4f",	--1321
		x"5f",	--1322
		x"4f",	--1323
		x"fa",	--1324
		x"41",	--1325
		x"41",	--1326
		x"41",	--1327
		x"41",	--1328
		x"4b",	--1329
		x"52",	--1330
		x"4b",	--1331
		x"00",	--1332
		x"4b",	--1333
		x"12",	--1334
		x"e8",	--1335
		x"49",	--1336
		x"3f",	--1337
		x"4b",	--1338
		x"53",	--1339
		x"4b",	--1340
		x"12",	--1341
		x"e8",	--1342
		x"49",	--1343
		x"3f",	--1344
		x"4b",	--1345
		x"53",	--1346
		x"4f",	--1347
		x"49",	--1348
		x"93",	--1349
		x"27",	--1350
		x"53",	--1351
		x"11",	--1352
		x"12",	--1353
		x"e8",	--1354
		x"49",	--1355
		x"93",	--1356
		x"23",	--1357
		x"3f",	--1358
		x"4b",	--1359
		x"52",	--1360
		x"4b",	--1361
		x"00",	--1362
		x"4b",	--1363
		x"12",	--1364
		x"e9",	--1365
		x"49",	--1366
		x"3f",	--1367
		x"4b",	--1368
		x"53",	--1369
		x"4b",	--1370
		x"4e",	--1371
		x"10",	--1372
		x"11",	--1373
		x"10",	--1374
		x"11",	--1375
		x"12",	--1376
		x"e8",	--1377
		x"49",	--1378
		x"3f",	--1379
		x"4b",	--1380
		x"53",	--1381
		x"4b",	--1382
		x"12",	--1383
		x"e9",	--1384
		x"49",	--1385
		x"3f",	--1386
		x"4b",	--1387
		x"53",	--1388
		x"4b",	--1389
		x"12",	--1390
		x"e8",	--1391
		x"49",	--1392
		x"3f",	--1393
		x"4b",	--1394
		x"53",	--1395
		x"4b",	--1396
		x"12",	--1397
		x"e8",	--1398
		x"49",	--1399
		x"3f",	--1400
		x"4b",	--1401
		x"53",	--1402
		x"4b",	--1403
		x"12",	--1404
		x"e8",	--1405
		x"49",	--1406
		x"3f",	--1407
		x"40",	--1408
		x"00",	--1409
		x"12",	--1410
		x"e8",	--1411
		x"3f",	--1412
		x"12",	--1413
		x"12",	--1414
		x"42",	--1415
		x"02",	--1416
		x"42",	--1417
		x"00",	--1418
		x"04",	--1419
		x"42",	--1420
		x"02",	--1421
		x"90",	--1422
		x"00",	--1423
		x"34",	--1424
		x"53",	--1425
		x"02",	--1426
		x"42",	--1427
		x"02",	--1428
		x"42",	--1429
		x"02",	--1430
		x"9f",	--1431
		x"20",	--1432
		x"53",	--1433
		x"02",	--1434
		x"40",	--1435
		x"00",	--1436
		x"00",	--1437
		x"41",	--1438
		x"41",	--1439
		x"c0",	--1440
		x"00",	--1441
		x"00",	--1442
		x"13",	--1443
		x"43",	--1444
		x"02",	--1445
		x"3f",	--1446
		x"40",	--1447
		x"09",	--1448
		x"00",	--1449
		x"40",	--1450
		x"00",	--1451
		x"00",	--1452
		x"41",	--1453
		x"42",	--1454
		x"02",	--1455
		x"42",	--1456
		x"02",	--1457
		x"9f",	--1458
		x"38",	--1459
		x"42",	--1460
		x"02",	--1461
		x"82",	--1462
		x"02",	--1463
		x"41",	--1464
		x"42",	--1465
		x"02",	--1466
		x"42",	--1467
		x"02",	--1468
		x"40",	--1469
		x"00",	--1470
		x"8d",	--1471
		x"8e",	--1472
		x"41",	--1473
		x"42",	--1474
		x"02",	--1475
		x"4f",	--1476
		x"04",	--1477
		x"42",	--1478
		x"02",	--1479
		x"42",	--1480
		x"02",	--1481
		x"9e",	--1482
		x"24",	--1483
		x"42",	--1484
		x"02",	--1485
		x"90",	--1486
		x"00",	--1487
		x"38",	--1488
		x"43",	--1489
		x"02",	--1490
		x"41",	--1491
		x"53",	--1492
		x"02",	--1493
		x"41",	--1494
		x"43",	--1495
		x"41",	--1496
		x"12",	--1497
		x"12",	--1498
		x"4e",	--1499
		x"4f",	--1500
		x"43",	--1501
		x"40",	--1502
		x"4f",	--1503
		x"12",	--1504
		x"f2",	--1505
		x"93",	--1506
		x"34",	--1507
		x"4a",	--1508
		x"4b",	--1509
		x"12",	--1510
		x"f2",	--1511
		x"41",	--1512
		x"41",	--1513
		x"41",	--1514
		x"43",	--1515
		x"40",	--1516
		x"4f",	--1517
		x"4a",	--1518
		x"4b",	--1519
		x"12",	--1520
		x"ee",	--1521
		x"12",	--1522
		x"f2",	--1523
		x"53",	--1524
		x"60",	--1525
		x"80",	--1526
		x"41",	--1527
		x"41",	--1528
		x"41",	--1529
		x"12",	--1530
		x"12",	--1531
		x"12",	--1532
		x"12",	--1533
		x"12",	--1534
		x"12",	--1535
		x"12",	--1536
		x"12",	--1537
		x"50",	--1538
		x"ff",	--1539
		x"4d",	--1540
		x"4f",	--1541
		x"93",	--1542
		x"28",	--1543
		x"4e",	--1544
		x"93",	--1545
		x"28",	--1546
		x"92",	--1547
		x"20",	--1548
		x"40",	--1549
		x"ee",	--1550
		x"92",	--1551
		x"24",	--1552
		x"93",	--1553
		x"24",	--1554
		x"93",	--1555
		x"24",	--1556
		x"4f",	--1557
		x"00",	--1558
		x"00",	--1559
		x"4e",	--1560
		x"00",	--1561
		x"4f",	--1562
		x"00",	--1563
		x"4f",	--1564
		x"00",	--1565
		x"4e",	--1566
		x"00",	--1567
		x"4e",	--1568
		x"00",	--1569
		x"41",	--1570
		x"8b",	--1571
		x"4c",	--1572
		x"93",	--1573
		x"38",	--1574
		x"90",	--1575
		x"00",	--1576
		x"34",	--1577
		x"93",	--1578
		x"38",	--1579
		x"46",	--1580
		x"00",	--1581
		x"47",	--1582
		x"00",	--1583
		x"49",	--1584
		x"f0",	--1585
		x"00",	--1586
		x"24",	--1587
		x"46",	--1588
		x"47",	--1589
		x"c3",	--1590
		x"10",	--1591
		x"10",	--1592
		x"53",	--1593
		x"23",	--1594
		x"4a",	--1595
		x"00",	--1596
		x"4b",	--1597
		x"00",	--1598
		x"43",	--1599
		x"43",	--1600
		x"f0",	--1601
		x"00",	--1602
		x"24",	--1603
		x"5c",	--1604
		x"6d",	--1605
		x"53",	--1606
		x"23",	--1607
		x"53",	--1608
		x"63",	--1609
		x"f6",	--1610
		x"f7",	--1611
		x"43",	--1612
		x"43",	--1613
		x"93",	--1614
		x"20",	--1615
		x"93",	--1616
		x"24",	--1617
		x"41",	--1618
		x"00",	--1619
		x"41",	--1620
		x"00",	--1621
		x"da",	--1622
		x"db",	--1623
		x"4f",	--1624
		x"00",	--1625
		x"9e",	--1626
		x"00",	--1627
		x"20",	--1628
		x"4f",	--1629
		x"00",	--1630
		x"41",	--1631
		x"00",	--1632
		x"46",	--1633
		x"47",	--1634
		x"54",	--1635
		x"65",	--1636
		x"4e",	--1637
		x"00",	--1638
		x"4f",	--1639
		x"00",	--1640
		x"40",	--1641
		x"00",	--1642
		x"00",	--1643
		x"93",	--1644
		x"38",	--1645
		x"48",	--1646
		x"50",	--1647
		x"00",	--1648
		x"41",	--1649
		x"41",	--1650
		x"41",	--1651
		x"41",	--1652
		x"41",	--1653
		x"41",	--1654
		x"41",	--1655
		x"41",	--1656
		x"41",	--1657
		x"91",	--1658
		x"38",	--1659
		x"4b",	--1660
		x"00",	--1661
		x"43",	--1662
		x"43",	--1663
		x"4f",	--1664
		x"00",	--1665
		x"9e",	--1666
		x"00",	--1667
		x"27",	--1668
		x"93",	--1669
		x"24",	--1670
		x"46",	--1671
		x"47",	--1672
		x"84",	--1673
		x"75",	--1674
		x"93",	--1675
		x"38",	--1676
		x"43",	--1677
		x"00",	--1678
		x"41",	--1679
		x"00",	--1680
		x"4e",	--1681
		x"00",	--1682
		x"4f",	--1683
		x"00",	--1684
		x"4e",	--1685
		x"4f",	--1686
		x"53",	--1687
		x"63",	--1688
		x"90",	--1689
		x"3f",	--1690
		x"28",	--1691
		x"90",	--1692
		x"40",	--1693
		x"2c",	--1694
		x"93",	--1695
		x"2c",	--1696
		x"48",	--1697
		x"00",	--1698
		x"53",	--1699
		x"5e",	--1700
		x"6f",	--1701
		x"4b",	--1702
		x"53",	--1703
		x"4e",	--1704
		x"4f",	--1705
		x"53",	--1706
		x"63",	--1707
		x"90",	--1708
		x"3f",	--1709
		x"2b",	--1710
		x"24",	--1711
		x"4e",	--1712
		x"00",	--1713
		x"4f",	--1714
		x"00",	--1715
		x"4a",	--1716
		x"00",	--1717
		x"40",	--1718
		x"00",	--1719
		x"00",	--1720
		x"93",	--1721
		x"37",	--1722
		x"4e",	--1723
		x"4f",	--1724
		x"f3",	--1725
		x"f3",	--1726
		x"c3",	--1727
		x"10",	--1728
		x"10",	--1729
		x"4c",	--1730
		x"4d",	--1731
		x"de",	--1732
		x"df",	--1733
		x"4a",	--1734
		x"00",	--1735
		x"4b",	--1736
		x"00",	--1737
		x"53",	--1738
		x"00",	--1739
		x"48",	--1740
		x"3f",	--1741
		x"93",	--1742
		x"23",	--1743
		x"4f",	--1744
		x"00",	--1745
		x"4f",	--1746
		x"00",	--1747
		x"00",	--1748
		x"4f",	--1749
		x"00",	--1750
		x"00",	--1751
		x"4f",	--1752
		x"00",	--1753
		x"00",	--1754
		x"4e",	--1755
		x"00",	--1756
		x"ff",	--1757
		x"00",	--1758
		x"4e",	--1759
		x"00",	--1760
		x"4d",	--1761
		x"3f",	--1762
		x"43",	--1763
		x"43",	--1764
		x"3f",	--1765
		x"e3",	--1766
		x"53",	--1767
		x"90",	--1768
		x"00",	--1769
		x"37",	--1770
		x"3f",	--1771
		x"93",	--1772
		x"2b",	--1773
		x"3f",	--1774
		x"44",	--1775
		x"45",	--1776
		x"86",	--1777
		x"77",	--1778
		x"3f",	--1779
		x"4e",	--1780
		x"3f",	--1781
		x"43",	--1782
		x"00",	--1783
		x"41",	--1784
		x"00",	--1785
		x"e3",	--1786
		x"e3",	--1787
		x"53",	--1788
		x"63",	--1789
		x"4e",	--1790
		x"00",	--1791
		x"4f",	--1792
		x"00",	--1793
		x"3f",	--1794
		x"93",	--1795
		x"27",	--1796
		x"59",	--1797
		x"00",	--1798
		x"44",	--1799
		x"00",	--1800
		x"45",	--1801
		x"00",	--1802
		x"49",	--1803
		x"f0",	--1804
		x"00",	--1805
		x"24",	--1806
		x"4d",	--1807
		x"44",	--1808
		x"45",	--1809
		x"c3",	--1810
		x"10",	--1811
		x"10",	--1812
		x"53",	--1813
		x"23",	--1814
		x"4c",	--1815
		x"00",	--1816
		x"4d",	--1817
		x"00",	--1818
		x"43",	--1819
		x"43",	--1820
		x"f0",	--1821
		x"00",	--1822
		x"24",	--1823
		x"5c",	--1824
		x"6d",	--1825
		x"53",	--1826
		x"23",	--1827
		x"53",	--1828
		x"63",	--1829
		x"f4",	--1830
		x"f5",	--1831
		x"43",	--1832
		x"43",	--1833
		x"93",	--1834
		x"20",	--1835
		x"93",	--1836
		x"20",	--1837
		x"43",	--1838
		x"43",	--1839
		x"41",	--1840
		x"00",	--1841
		x"41",	--1842
		x"00",	--1843
		x"da",	--1844
		x"db",	--1845
		x"3f",	--1846
		x"43",	--1847
		x"43",	--1848
		x"3f",	--1849
		x"92",	--1850
		x"23",	--1851
		x"9e",	--1852
		x"00",	--1853
		x"00",	--1854
		x"27",	--1855
		x"40",	--1856
		x"fb",	--1857
		x"3f",	--1858
		x"50",	--1859
		x"ff",	--1860
		x"4e",	--1861
		x"00",	--1862
		x"4f",	--1863
		x"00",	--1864
		x"4c",	--1865
		x"00",	--1866
		x"4d",	--1867
		x"00",	--1868
		x"41",	--1869
		x"50",	--1870
		x"00",	--1871
		x"41",	--1872
		x"52",	--1873
		x"12",	--1874
		x"f6",	--1875
		x"41",	--1876
		x"50",	--1877
		x"00",	--1878
		x"41",	--1879
		x"12",	--1880
		x"f6",	--1881
		x"41",	--1882
		x"52",	--1883
		x"41",	--1884
		x"50",	--1885
		x"00",	--1886
		x"41",	--1887
		x"50",	--1888
		x"00",	--1889
		x"12",	--1890
		x"eb",	--1891
		x"12",	--1892
		x"f4",	--1893
		x"50",	--1894
		x"00",	--1895
		x"41",	--1896
		x"50",	--1897
		x"ff",	--1898
		x"4e",	--1899
		x"00",	--1900
		x"4f",	--1901
		x"00",	--1902
		x"4c",	--1903
		x"00",	--1904
		x"4d",	--1905
		x"00",	--1906
		x"41",	--1907
		x"50",	--1908
		x"00",	--1909
		x"41",	--1910
		x"52",	--1911
		x"12",	--1912
		x"f6",	--1913
		x"41",	--1914
		x"50",	--1915
		x"00",	--1916
		x"41",	--1917
		x"12",	--1918
		x"f6",	--1919
		x"e3",	--1920
		x"00",	--1921
		x"41",	--1922
		x"52",	--1923
		x"41",	--1924
		x"50",	--1925
		x"00",	--1926
		x"41",	--1927
		x"50",	--1928
		x"00",	--1929
		x"12",	--1930
		x"eb",	--1931
		x"12",	--1932
		x"f4",	--1933
		x"50",	--1934
		x"00",	--1935
		x"41",	--1936
		x"12",	--1937
		x"12",	--1938
		x"12",	--1939
		x"12",	--1940
		x"12",	--1941
		x"12",	--1942
		x"12",	--1943
		x"12",	--1944
		x"50",	--1945
		x"ff",	--1946
		x"4e",	--1947
		x"00",	--1948
		x"4f",	--1949
		x"00",	--1950
		x"4c",	--1951
		x"00",	--1952
		x"4d",	--1953
		x"00",	--1954
		x"41",	--1955
		x"50",	--1956
		x"00",	--1957
		x"41",	--1958
		x"52",	--1959
		x"12",	--1960
		x"f6",	--1961
		x"41",	--1962
		x"50",	--1963
		x"00",	--1964
		x"41",	--1965
		x"12",	--1966
		x"f6",	--1967
		x"41",	--1968
		x"00",	--1969
		x"93",	--1970
		x"28",	--1971
		x"41",	--1972
		x"00",	--1973
		x"93",	--1974
		x"28",	--1975
		x"92",	--1976
		x"24",	--1977
		x"92",	--1978
		x"24",	--1979
		x"93",	--1980
		x"24",	--1981
		x"93",	--1982
		x"24",	--1983
		x"41",	--1984
		x"00",	--1985
		x"41",	--1986
		x"00",	--1987
		x"41",	--1988
		x"00",	--1989
		x"41",	--1990
		x"00",	--1991
		x"40",	--1992
		x"00",	--1993
		x"43",	--1994
		x"43",	--1995
		x"43",	--1996
		x"43",	--1997
		x"43",	--1998
		x"00",	--1999
		x"43",	--2000
		x"00",	--2001
		x"43",	--2002
		x"43",	--2003
		x"4c",	--2004
		x"00",	--2005
		x"3c",	--2006
		x"58",	--2007
		x"69",	--2008
		x"c3",	--2009
		x"10",	--2010
		x"10",	--2011
		x"53",	--2012
		x"00",	--2013
		x"24",	--2014
		x"b3",	--2015
		x"24",	--2016
		x"58",	--2017
		x"69",	--2018
		x"56",	--2019
		x"67",	--2020
		x"43",	--2021
		x"43",	--2022
		x"99",	--2023
		x"28",	--2024
		x"24",	--2025
		x"43",	--2026
		x"43",	--2027
		x"5c",	--2028
		x"6d",	--2029
		x"56",	--2030
		x"67",	--2031
		x"93",	--2032
		x"37",	--2033
		x"d3",	--2034
		x"d3",	--2035
		x"3f",	--2036
		x"98",	--2037
		x"2b",	--2038
		x"3f",	--2039
		x"4a",	--2040
		x"00",	--2041
		x"4b",	--2042
		x"00",	--2043
		x"4f",	--2044
		x"41",	--2045
		x"00",	--2046
		x"51",	--2047
		x"00",	--2048
		x"4a",	--2049
		x"53",	--2050
		x"46",	--2051
		x"00",	--2052
		x"43",	--2053
		x"91",	--2054
		x"00",	--2055
		x"00",	--2056
		x"24",	--2057
		x"4d",	--2058
		x"00",	--2059
		x"93",	--2060
		x"38",	--2061
		x"90",	--2062
		x"40",	--2063
		x"2c",	--2064
		x"41",	--2065
		x"00",	--2066
		x"53",	--2067
		x"41",	--2068
		x"00",	--2069
		x"41",	--2070
		x"00",	--2071
		x"4d",	--2072
		x"5e",	--2073
		x"6f",	--2074
		x"93",	--2075
		x"38",	--2076
		x"5a",	--2077
		x"6b",	--2078
		x"53",	--2079
		x"90",	--2080
		x"40",	--2081
		x"2b",	--2082
		x"4a",	--2083
		x"00",	--2084
		x"4b",	--2085
		x"00",	--2086
		x"4c",	--2087
		x"00",	--2088
		x"4e",	--2089
		x"4f",	--2090
		x"f0",	--2091
		x"00",	--2092
		x"f3",	--2093
		x"90",	--2094
		x"00",	--2095
		x"24",	--2096
		x"4e",	--2097
		x"00",	--2098
		x"4f",	--2099
		x"00",	--2100
		x"40",	--2101
		x"00",	--2102
		x"00",	--2103
		x"41",	--2104
		x"52",	--2105
		x"12",	--2106
		x"f4",	--2107
		x"50",	--2108
		x"00",	--2109
		x"41",	--2110
		x"41",	--2111
		x"41",	--2112
		x"41",	--2113
		x"41",	--2114
		x"41",	--2115
		x"41",	--2116
		x"41",	--2117
		x"41",	--2118
		x"d3",	--2119
		x"d3",	--2120
		x"3f",	--2121
		x"50",	--2122
		x"00",	--2123
		x"4a",	--2124
		x"b3",	--2125
		x"24",	--2126
		x"41",	--2127
		x"00",	--2128
		x"41",	--2129
		x"00",	--2130
		x"c3",	--2131
		x"10",	--2132
		x"10",	--2133
		x"4c",	--2134
		x"4d",	--2135
		x"d3",	--2136
		x"d0",	--2137
		x"80",	--2138
		x"46",	--2139
		x"00",	--2140
		x"47",	--2141
		x"00",	--2142
		x"c3",	--2143
		x"10",	--2144
		x"10",	--2145
		x"53",	--2146
		x"93",	--2147
		x"3b",	--2148
		x"48",	--2149
		x"00",	--2150
		x"3f",	--2151
		x"93",	--2152
		x"24",	--2153
		x"43",	--2154
		x"91",	--2155
		x"00",	--2156
		x"00",	--2157
		x"24",	--2158
		x"4f",	--2159
		x"00",	--2160
		x"41",	--2161
		x"50",	--2162
		x"00",	--2163
		x"3f",	--2164
		x"93",	--2165
		x"23",	--2166
		x"4e",	--2167
		x"4f",	--2168
		x"f0",	--2169
		x"00",	--2170
		x"f3",	--2171
		x"93",	--2172
		x"23",	--2173
		x"93",	--2174
		x"23",	--2175
		x"93",	--2176
		x"00",	--2177
		x"20",	--2178
		x"93",	--2179
		x"00",	--2180
		x"27",	--2181
		x"50",	--2182
		x"00",	--2183
		x"63",	--2184
		x"f0",	--2185
		x"ff",	--2186
		x"f3",	--2187
		x"3f",	--2188
		x"43",	--2189
		x"3f",	--2190
		x"43",	--2191
		x"3f",	--2192
		x"43",	--2193
		x"91",	--2194
		x"00",	--2195
		x"00",	--2196
		x"24",	--2197
		x"4f",	--2198
		x"00",	--2199
		x"41",	--2200
		x"50",	--2201
		x"00",	--2202
		x"3f",	--2203
		x"43",	--2204
		x"3f",	--2205
		x"93",	--2206
		x"23",	--2207
		x"40",	--2208
		x"fb",	--2209
		x"3f",	--2210
		x"12",	--2211
		x"12",	--2212
		x"12",	--2213
		x"12",	--2214
		x"12",	--2215
		x"50",	--2216
		x"ff",	--2217
		x"4e",	--2218
		x"00",	--2219
		x"4f",	--2220
		x"00",	--2221
		x"4c",	--2222
		x"00",	--2223
		x"4d",	--2224
		x"00",	--2225
		x"41",	--2226
		x"50",	--2227
		x"00",	--2228
		x"41",	--2229
		x"52",	--2230
		x"12",	--2231
		x"f6",	--2232
		x"41",	--2233
		x"52",	--2234
		x"41",	--2235
		x"12",	--2236
		x"f6",	--2237
		x"41",	--2238
		x"00",	--2239
		x"93",	--2240
		x"28",	--2241
		x"41",	--2242
		x"00",	--2243
		x"93",	--2244
		x"28",	--2245
		x"e1",	--2246
		x"00",	--2247
		x"00",	--2248
		x"92",	--2249
		x"24",	--2250
		x"93",	--2251
		x"24",	--2252
		x"92",	--2253
		x"24",	--2254
		x"93",	--2255
		x"24",	--2256
		x"41",	--2257
		x"00",	--2258
		x"81",	--2259
		x"00",	--2260
		x"4d",	--2261
		x"00",	--2262
		x"41",	--2263
		x"00",	--2264
		x"41",	--2265
		x"00",	--2266
		x"41",	--2267
		x"00",	--2268
		x"41",	--2269
		x"00",	--2270
		x"99",	--2271
		x"2c",	--2272
		x"5e",	--2273
		x"6f",	--2274
		x"53",	--2275
		x"4d",	--2276
		x"00",	--2277
		x"40",	--2278
		x"00",	--2279
		x"43",	--2280
		x"40",	--2281
		x"40",	--2282
		x"43",	--2283
		x"43",	--2284
		x"3c",	--2285
		x"dc",	--2286
		x"dd",	--2287
		x"88",	--2288
		x"79",	--2289
		x"c3",	--2290
		x"10",	--2291
		x"10",	--2292
		x"5e",	--2293
		x"6f",	--2294
		x"53",	--2295
		x"24",	--2296
		x"99",	--2297
		x"2b",	--2298
		x"23",	--2299
		x"98",	--2300
		x"2b",	--2301
		x"3f",	--2302
		x"9f",	--2303
		x"2b",	--2304
		x"98",	--2305
		x"2f",	--2306
		x"3f",	--2307
		x"4a",	--2308
		x"4b",	--2309
		x"f0",	--2310
		x"00",	--2311
		x"f3",	--2312
		x"90",	--2313
		x"00",	--2314
		x"24",	--2315
		x"4a",	--2316
		x"00",	--2317
		x"4b",	--2318
		x"00",	--2319
		x"41",	--2320
		x"50",	--2321
		x"00",	--2322
		x"12",	--2323
		x"f4",	--2324
		x"50",	--2325
		x"00",	--2326
		x"41",	--2327
		x"41",	--2328
		x"41",	--2329
		x"41",	--2330
		x"41",	--2331
		x"41",	--2332
		x"42",	--2333
		x"00",	--2334
		x"41",	--2335
		x"50",	--2336
		x"00",	--2337
		x"3f",	--2338
		x"9e",	--2339
		x"23",	--2340
		x"40",	--2341
		x"fb",	--2342
		x"3f",	--2343
		x"93",	--2344
		x"23",	--2345
		x"4a",	--2346
		x"4b",	--2347
		x"f0",	--2348
		x"00",	--2349
		x"f3",	--2350
		x"93",	--2351
		x"23",	--2352
		x"93",	--2353
		x"23",	--2354
		x"93",	--2355
		x"20",	--2356
		x"93",	--2357
		x"27",	--2358
		x"50",	--2359
		x"00",	--2360
		x"63",	--2361
		x"f0",	--2362
		x"ff",	--2363
		x"f3",	--2364
		x"3f",	--2365
		x"43",	--2366
		x"00",	--2367
		x"43",	--2368
		x"00",	--2369
		x"43",	--2370
		x"00",	--2371
		x"41",	--2372
		x"50",	--2373
		x"00",	--2374
		x"3f",	--2375
		x"41",	--2376
		x"52",	--2377
		x"3f",	--2378
		x"50",	--2379
		x"ff",	--2380
		x"4e",	--2381
		x"00",	--2382
		x"4f",	--2383
		x"00",	--2384
		x"4c",	--2385
		x"00",	--2386
		x"4d",	--2387
		x"00",	--2388
		x"41",	--2389
		x"50",	--2390
		x"00",	--2391
		x"41",	--2392
		x"52",	--2393
		x"12",	--2394
		x"f6",	--2395
		x"41",	--2396
		x"52",	--2397
		x"41",	--2398
		x"12",	--2399
		x"f6",	--2400
		x"93",	--2401
		x"00",	--2402
		x"28",	--2403
		x"93",	--2404
		x"00",	--2405
		x"28",	--2406
		x"41",	--2407
		x"52",	--2408
		x"41",	--2409
		x"50",	--2410
		x"00",	--2411
		x"12",	--2412
		x"f7",	--2413
		x"50",	--2414
		x"00",	--2415
		x"41",	--2416
		x"43",	--2417
		x"3f",	--2418
		x"50",	--2419
		x"ff",	--2420
		x"4e",	--2421
		x"00",	--2422
		x"4f",	--2423
		x"00",	--2424
		x"41",	--2425
		x"52",	--2426
		x"41",	--2427
		x"12",	--2428
		x"f6",	--2429
		x"41",	--2430
		x"00",	--2431
		x"93",	--2432
		x"24",	--2433
		x"28",	--2434
		x"92",	--2435
		x"24",	--2436
		x"41",	--2437
		x"00",	--2438
		x"93",	--2439
		x"38",	--2440
		x"90",	--2441
		x"00",	--2442
		x"38",	--2443
		x"93",	--2444
		x"00",	--2445
		x"20",	--2446
		x"43",	--2447
		x"40",	--2448
		x"7f",	--2449
		x"50",	--2450
		x"00",	--2451
		x"41",	--2452
		x"41",	--2453
		x"00",	--2454
		x"41",	--2455
		x"00",	--2456
		x"40",	--2457
		x"00",	--2458
		x"8d",	--2459
		x"4c",	--2460
		x"f0",	--2461
		x"00",	--2462
		x"20",	--2463
		x"93",	--2464
		x"00",	--2465
		x"27",	--2466
		x"e3",	--2467
		x"e3",	--2468
		x"53",	--2469
		x"63",	--2470
		x"50",	--2471
		x"00",	--2472
		x"41",	--2473
		x"43",	--2474
		x"43",	--2475
		x"50",	--2476
		x"00",	--2477
		x"41",	--2478
		x"c3",	--2479
		x"10",	--2480
		x"10",	--2481
		x"53",	--2482
		x"23",	--2483
		x"3f",	--2484
		x"43",	--2485
		x"40",	--2486
		x"80",	--2487
		x"50",	--2488
		x"00",	--2489
		x"41",	--2490
		x"12",	--2491
		x"12",	--2492
		x"12",	--2493
		x"12",	--2494
		x"82",	--2495
		x"4e",	--2496
		x"4f",	--2497
		x"43",	--2498
		x"00",	--2499
		x"93",	--2500
		x"20",	--2501
		x"93",	--2502
		x"20",	--2503
		x"43",	--2504
		x"00",	--2505
		x"41",	--2506
		x"12",	--2507
		x"f4",	--2508
		x"52",	--2509
		x"41",	--2510
		x"41",	--2511
		x"41",	--2512
		x"41",	--2513
		x"41",	--2514
		x"40",	--2515
		x"00",	--2516
		x"00",	--2517
		x"40",	--2518
		x"00",	--2519
		x"00",	--2520
		x"4a",	--2521
		x"00",	--2522
		x"4b",	--2523
		x"00",	--2524
		x"4a",	--2525
		x"4b",	--2526
		x"12",	--2527
		x"f4",	--2528
		x"53",	--2529
		x"93",	--2530
		x"38",	--2531
		x"27",	--2532
		x"4a",	--2533
		x"00",	--2534
		x"4b",	--2535
		x"00",	--2536
		x"4f",	--2537
		x"f0",	--2538
		x"00",	--2539
		x"20",	--2540
		x"40",	--2541
		x"00",	--2542
		x"8f",	--2543
		x"4e",	--2544
		x"00",	--2545
		x"3f",	--2546
		x"51",	--2547
		x"00",	--2548
		x"00",	--2549
		x"61",	--2550
		x"00",	--2551
		x"00",	--2552
		x"53",	--2553
		x"23",	--2554
		x"3f",	--2555
		x"4f",	--2556
		x"e3",	--2557
		x"53",	--2558
		x"43",	--2559
		x"43",	--2560
		x"4e",	--2561
		x"f0",	--2562
		x"00",	--2563
		x"24",	--2564
		x"5c",	--2565
		x"6d",	--2566
		x"53",	--2567
		x"23",	--2568
		x"53",	--2569
		x"63",	--2570
		x"fa",	--2571
		x"fb",	--2572
		x"43",	--2573
		x"43",	--2574
		x"93",	--2575
		x"20",	--2576
		x"93",	--2577
		x"20",	--2578
		x"43",	--2579
		x"43",	--2580
		x"f0",	--2581
		x"00",	--2582
		x"20",	--2583
		x"48",	--2584
		x"49",	--2585
		x"da",	--2586
		x"db",	--2587
		x"4d",	--2588
		x"00",	--2589
		x"4e",	--2590
		x"00",	--2591
		x"40",	--2592
		x"00",	--2593
		x"8f",	--2594
		x"4e",	--2595
		x"00",	--2596
		x"3f",	--2597
		x"c3",	--2598
		x"10",	--2599
		x"10",	--2600
		x"53",	--2601
		x"23",	--2602
		x"3f",	--2603
		x"12",	--2604
		x"12",	--2605
		x"12",	--2606
		x"93",	--2607
		x"2c",	--2608
		x"90",	--2609
		x"01",	--2610
		x"28",	--2611
		x"40",	--2612
		x"00",	--2613
		x"43",	--2614
		x"42",	--2615
		x"4e",	--2616
		x"4f",	--2617
		x"49",	--2618
		x"93",	--2619
		x"20",	--2620
		x"50",	--2621
		x"fb",	--2622
		x"4c",	--2623
		x"43",	--2624
		x"8e",	--2625
		x"7f",	--2626
		x"4a",	--2627
		x"41",	--2628
		x"41",	--2629
		x"41",	--2630
		x"41",	--2631
		x"90",	--2632
		x"01",	--2633
		x"28",	--2634
		x"42",	--2635
		x"43",	--2636
		x"40",	--2637
		x"00",	--2638
		x"4e",	--2639
		x"4f",	--2640
		x"49",	--2641
		x"93",	--2642
		x"27",	--2643
		x"c3",	--2644
		x"10",	--2645
		x"10",	--2646
		x"53",	--2647
		x"23",	--2648
		x"3f",	--2649
		x"40",	--2650
		x"00",	--2651
		x"43",	--2652
		x"40",	--2653
		x"00",	--2654
		x"3f",	--2655
		x"40",	--2656
		x"00",	--2657
		x"43",	--2658
		x"43",	--2659
		x"3f",	--2660
		x"12",	--2661
		x"12",	--2662
		x"12",	--2663
		x"12",	--2664
		x"12",	--2665
		x"4f",	--2666
		x"4f",	--2667
		x"00",	--2668
		x"4f",	--2669
		x"00",	--2670
		x"4d",	--2671
		x"00",	--2672
		x"4d",	--2673
		x"93",	--2674
		x"28",	--2675
		x"92",	--2676
		x"24",	--2677
		x"93",	--2678
		x"24",	--2679
		x"93",	--2680
		x"24",	--2681
		x"4d",	--2682
		x"00",	--2683
		x"90",	--2684
		x"ff",	--2685
		x"38",	--2686
		x"90",	--2687
		x"00",	--2688
		x"34",	--2689
		x"4e",	--2690
		x"4f",	--2691
		x"f0",	--2692
		x"00",	--2693
		x"f3",	--2694
		x"90",	--2695
		x"00",	--2696
		x"24",	--2697
		x"50",	--2698
		x"00",	--2699
		x"63",	--2700
		x"93",	--2701
		x"38",	--2702
		x"4b",	--2703
		x"50",	--2704
		x"00",	--2705
		x"c3",	--2706
		x"10",	--2707
		x"10",	--2708
		x"c3",	--2709
		x"10",	--2710
		x"10",	--2711
		x"c3",	--2712
		x"10",	--2713
		x"10",	--2714
		x"c3",	--2715
		x"10",	--2716
		x"10",	--2717
		x"c3",	--2718
		x"10",	--2719
		x"10",	--2720
		x"c3",	--2721
		x"10",	--2722
		x"10",	--2723
		x"c3",	--2724
		x"10",	--2725
		x"10",	--2726
		x"f3",	--2727
		x"f0",	--2728
		x"00",	--2729
		x"4d",	--2730
		x"3c",	--2731
		x"93",	--2732
		x"23",	--2733
		x"43",	--2734
		x"43",	--2735
		x"43",	--2736
		x"4d",	--2737
		x"5d",	--2738
		x"5d",	--2739
		x"5d",	--2740
		x"5d",	--2741
		x"5d",	--2742
		x"5d",	--2743
		x"5d",	--2744
		x"4f",	--2745
		x"f0",	--2746
		x"00",	--2747
		x"dd",	--2748
		x"4a",	--2749
		x"11",	--2750
		x"43",	--2751
		x"10",	--2752
		x"4c",	--2753
		x"df",	--2754
		x"4d",	--2755
		x"41",	--2756
		x"41",	--2757
		x"41",	--2758
		x"41",	--2759
		x"41",	--2760
		x"41",	--2761
		x"93",	--2762
		x"23",	--2763
		x"4e",	--2764
		x"4f",	--2765
		x"f0",	--2766
		x"00",	--2767
		x"f3",	--2768
		x"93",	--2769
		x"20",	--2770
		x"93",	--2771
		x"27",	--2772
		x"50",	--2773
		x"00",	--2774
		x"63",	--2775
		x"3f",	--2776
		x"c3",	--2777
		x"10",	--2778
		x"10",	--2779
		x"4b",	--2780
		x"50",	--2781
		x"00",	--2782
		x"3f",	--2783
		x"43",	--2784
		x"43",	--2785
		x"43",	--2786
		x"3f",	--2787
		x"d3",	--2788
		x"d0",	--2789
		x"00",	--2790
		x"f3",	--2791
		x"f0",	--2792
		x"00",	--2793
		x"43",	--2794
		x"3f",	--2795
		x"40",	--2796
		x"ff",	--2797
		x"8b",	--2798
		x"90",	--2799
		x"00",	--2800
		x"34",	--2801
		x"4e",	--2802
		x"4f",	--2803
		x"47",	--2804
		x"f0",	--2805
		x"00",	--2806
		x"24",	--2807
		x"c3",	--2808
		x"10",	--2809
		x"10",	--2810
		x"53",	--2811
		x"23",	--2812
		x"43",	--2813
		x"43",	--2814
		x"f0",	--2815
		x"00",	--2816
		x"24",	--2817
		x"58",	--2818
		x"69",	--2819
		x"53",	--2820
		x"23",	--2821
		x"53",	--2822
		x"63",	--2823
		x"fe",	--2824
		x"ff",	--2825
		x"43",	--2826
		x"43",	--2827
		x"93",	--2828
		x"20",	--2829
		x"93",	--2830
		x"20",	--2831
		x"43",	--2832
		x"43",	--2833
		x"4e",	--2834
		x"4f",	--2835
		x"dc",	--2836
		x"dd",	--2837
		x"48",	--2838
		x"49",	--2839
		x"f0",	--2840
		x"00",	--2841
		x"f3",	--2842
		x"90",	--2843
		x"00",	--2844
		x"24",	--2845
		x"50",	--2846
		x"00",	--2847
		x"63",	--2848
		x"48",	--2849
		x"49",	--2850
		x"c3",	--2851
		x"10",	--2852
		x"10",	--2853
		x"c3",	--2854
		x"10",	--2855
		x"10",	--2856
		x"c3",	--2857
		x"10",	--2858
		x"10",	--2859
		x"c3",	--2860
		x"10",	--2861
		x"10",	--2862
		x"c3",	--2863
		x"10",	--2864
		x"10",	--2865
		x"c3",	--2866
		x"10",	--2867
		x"10",	--2868
		x"c3",	--2869
		x"10",	--2870
		x"10",	--2871
		x"f3",	--2872
		x"f0",	--2873
		x"00",	--2874
		x"43",	--2875
		x"90",	--2876
		x"40",	--2877
		x"2f",	--2878
		x"43",	--2879
		x"3f",	--2880
		x"43",	--2881
		x"43",	--2882
		x"3f",	--2883
		x"93",	--2884
		x"23",	--2885
		x"48",	--2886
		x"49",	--2887
		x"f0",	--2888
		x"00",	--2889
		x"f3",	--2890
		x"93",	--2891
		x"24",	--2892
		x"50",	--2893
		x"00",	--2894
		x"63",	--2895
		x"3f",	--2896
		x"93",	--2897
		x"27",	--2898
		x"3f",	--2899
		x"12",	--2900
		x"12",	--2901
		x"4f",	--2902
		x"4f",	--2903
		x"00",	--2904
		x"f0",	--2905
		x"00",	--2906
		x"4f",	--2907
		x"00",	--2908
		x"c3",	--2909
		x"10",	--2910
		x"c3",	--2911
		x"10",	--2912
		x"c3",	--2913
		x"10",	--2914
		x"c3",	--2915
		x"10",	--2916
		x"c3",	--2917
		x"10",	--2918
		x"c3",	--2919
		x"10",	--2920
		x"c3",	--2921
		x"10",	--2922
		x"4d",	--2923
		x"4f",	--2924
		x"00",	--2925
		x"b0",	--2926
		x"00",	--2927
		x"43",	--2928
		x"6f",	--2929
		x"4f",	--2930
		x"00",	--2931
		x"93",	--2932
		x"20",	--2933
		x"93",	--2934
		x"24",	--2935
		x"40",	--2936
		x"ff",	--2937
		x"00",	--2938
		x"4a",	--2939
		x"4b",	--2940
		x"5c",	--2941
		x"6d",	--2942
		x"5c",	--2943
		x"6d",	--2944
		x"5c",	--2945
		x"6d",	--2946
		x"5c",	--2947
		x"6d",	--2948
		x"5c",	--2949
		x"6d",	--2950
		x"5c",	--2951
		x"6d",	--2952
		x"5c",	--2953
		x"6d",	--2954
		x"40",	--2955
		x"00",	--2956
		x"00",	--2957
		x"90",	--2958
		x"40",	--2959
		x"2c",	--2960
		x"40",	--2961
		x"ff",	--2962
		x"5c",	--2963
		x"6d",	--2964
		x"4f",	--2965
		x"53",	--2966
		x"90",	--2967
		x"40",	--2968
		x"2b",	--2969
		x"4a",	--2970
		x"00",	--2971
		x"4c",	--2972
		x"00",	--2973
		x"4d",	--2974
		x"00",	--2975
		x"41",	--2976
		x"41",	--2977
		x"41",	--2978
		x"90",	--2979
		x"00",	--2980
		x"24",	--2981
		x"50",	--2982
		x"ff",	--2983
		x"4d",	--2984
		x"00",	--2985
		x"40",	--2986
		x"00",	--2987
		x"00",	--2988
		x"4a",	--2989
		x"4b",	--2990
		x"5c",	--2991
		x"6d",	--2992
		x"5c",	--2993
		x"6d",	--2994
		x"5c",	--2995
		x"6d",	--2996
		x"5c",	--2997
		x"6d",	--2998
		x"5c",	--2999
		x"6d",	--3000
		x"5c",	--3001
		x"6d",	--3002
		x"5c",	--3003
		x"6d",	--3004
		x"4c",	--3005
		x"4d",	--3006
		x"d3",	--3007
		x"d0",	--3008
		x"40",	--3009
		x"4a",	--3010
		x"00",	--3011
		x"4b",	--3012
		x"00",	--3013
		x"41",	--3014
		x"41",	--3015
		x"41",	--3016
		x"93",	--3017
		x"23",	--3018
		x"43",	--3019
		x"00",	--3020
		x"41",	--3021
		x"41",	--3022
		x"41",	--3023
		x"93",	--3024
		x"24",	--3025
		x"4a",	--3026
		x"4b",	--3027
		x"f3",	--3028
		x"f0",	--3029
		x"00",	--3030
		x"93",	--3031
		x"20",	--3032
		x"93",	--3033
		x"24",	--3034
		x"43",	--3035
		x"00",	--3036
		x"3f",	--3037
		x"93",	--3038
		x"23",	--3039
		x"42",	--3040
		x"00",	--3041
		x"3f",	--3042
		x"43",	--3043
		x"00",	--3044
		x"3f",	--3045
		x"12",	--3046
		x"4f",	--3047
		x"93",	--3048
		x"28",	--3049
		x"4e",	--3050
		x"93",	--3051
		x"28",	--3052
		x"92",	--3053
		x"24",	--3054
		x"92",	--3055
		x"24",	--3056
		x"93",	--3057
		x"24",	--3058
		x"93",	--3059
		x"24",	--3060
		x"4f",	--3061
		x"00",	--3062
		x"9e",	--3063
		x"00",	--3064
		x"24",	--3065
		x"93",	--3066
		x"20",	--3067
		x"43",	--3068
		x"4e",	--3069
		x"41",	--3070
		x"41",	--3071
		x"93",	--3072
		x"24",	--3073
		x"93",	--3074
		x"00",	--3075
		x"23",	--3076
		x"43",	--3077
		x"4e",	--3078
		x"41",	--3079
		x"41",	--3080
		x"93",	--3081
		x"00",	--3082
		x"27",	--3083
		x"43",	--3084
		x"3f",	--3085
		x"4f",	--3086
		x"00",	--3087
		x"4e",	--3088
		x"00",	--3089
		x"9b",	--3090
		x"3b",	--3091
		x"9c",	--3092
		x"38",	--3093
		x"4f",	--3094
		x"00",	--3095
		x"4f",	--3096
		x"00",	--3097
		x"4e",	--3098
		x"00",	--3099
		x"4e",	--3100
		x"00",	--3101
		x"9f",	--3102
		x"2b",	--3103
		x"9e",	--3104
		x"28",	--3105
		x"9b",	--3106
		x"2b",	--3107
		x"9e",	--3108
		x"28",	--3109
		x"9f",	--3110
		x"28",	--3111
		x"9c",	--3112
		x"28",	--3113
		x"43",	--3114
		x"3f",	--3115
		x"93",	--3116
		x"23",	--3117
		x"43",	--3118
		x"3f",	--3119
		x"92",	--3120
		x"23",	--3121
		x"4e",	--3122
		x"00",	--3123
		x"4f",	--3124
		x"00",	--3125
		x"8f",	--3126
		x"3f",	--3127
		x"43",	--3128
		x"93",	--3129
		x"34",	--3130
		x"40",	--3131
		x"00",	--3132
		x"e3",	--3133
		x"53",	--3134
		x"93",	--3135
		x"34",	--3136
		x"e3",	--3137
		x"e3",	--3138
		x"53",	--3139
		x"12",	--3140
		x"12",	--3141
		x"f8",	--3142
		x"41",	--3143
		x"b3",	--3144
		x"24",	--3145
		x"e3",	--3146
		x"53",	--3147
		x"b3",	--3148
		x"24",	--3149
		x"e3",	--3150
		x"53",	--3151
		x"41",	--3152
		x"12",	--3153
		x"f8",	--3154
		x"4e",	--3155
		x"41",	--3156
		x"12",	--3157
		x"43",	--3158
		x"93",	--3159
		x"34",	--3160
		x"40",	--3161
		x"00",	--3162
		x"e3",	--3163
		x"e3",	--3164
		x"53",	--3165
		x"63",	--3166
		x"93",	--3167
		x"34",	--3168
		x"e3",	--3169
		x"e3",	--3170
		x"e3",	--3171
		x"53",	--3172
		x"63",	--3173
		x"12",	--3174
		x"f9",	--3175
		x"b3",	--3176
		x"24",	--3177
		x"e3",	--3178
		x"e3",	--3179
		x"53",	--3180
		x"63",	--3181
		x"b3",	--3182
		x"24",	--3183
		x"e3",	--3184
		x"e3",	--3185
		x"53",	--3186
		x"63",	--3187
		x"41",	--3188
		x"41",	--3189
		x"12",	--3190
		x"f8",	--3191
		x"4c",	--3192
		x"4d",	--3193
		x"41",	--3194
		x"40",	--3195
		x"00",	--3196
		x"4e",	--3197
		x"43",	--3198
		x"5f",	--3199
		x"6e",	--3200
		x"9d",	--3201
		x"28",	--3202
		x"8d",	--3203
		x"d3",	--3204
		x"83",	--3205
		x"23",	--3206
		x"41",	--3207
		x"12",	--3208
		x"f8",	--3209
		x"4e",	--3210
		x"41",	--3211
		x"12",	--3212
		x"12",	--3213
		x"12",	--3214
		x"40",	--3215
		x"00",	--3216
		x"4c",	--3217
		x"4d",	--3218
		x"43",	--3219
		x"43",	--3220
		x"5e",	--3221
		x"6f",	--3222
		x"6c",	--3223
		x"6d",	--3224
		x"9b",	--3225
		x"28",	--3226
		x"20",	--3227
		x"9a",	--3228
		x"28",	--3229
		x"8a",	--3230
		x"7b",	--3231
		x"d3",	--3232
		x"83",	--3233
		x"23",	--3234
		x"41",	--3235
		x"41",	--3236
		x"41",	--3237
		x"41",	--3238
		x"12",	--3239
		x"f9",	--3240
		x"4c",	--3241
		x"4d",	--3242
		x"41",	--3243
		x"13",	--3244
		x"d0",	--3245
		x"00",	--3246
		x"3f",	--3247
		x"61",	--3248
		x"74",	--3249
		x"6e",	--3250
		x"20",	--3251
		x"6f",	--3252
		x"20",	--3253
		x"20",	--3254
		x"65",	--3255
		x"20",	--3256
		x"62",	--3257
		x"6e",	--3258
		x"66",	--3259
		x"6c",	--3260
		x"0d",	--3261
		x"00",	--3262
		x"65",	--3263
		x"73",	--3264
		x"6f",	--3265
		x"6c",	--3266
		x"20",	--3267
		x"6f",	--3268
		x"20",	--3269
		x"65",	--3270
		x"20",	--3271
		x"68",	--3272
		x"74",	--3273
		x"0a",	--3274
		x"63",	--3275
		x"72",	--3276
		x"65",	--3277
		x"74",	--3278
		x"75",	--3279
		x"61",	--3280
		x"65",	--3281
		x"0d",	--3282
		x"00",	--3283
		x"25",	--3284
		x"20",	--3285
		x"45",	--3286
		x"54",	--3287
		x"52",	--3288
		x"47",	--3289
		x"54",	--3290
		x"0a",	--3291
		x"53",	--3292
		x"6d",	--3293
		x"74",	--3294
		x"69",	--3295
		x"67",	--3296
		x"77",	--3297
		x"6e",	--3298
		x"20",	--3299
		x"65",	--3300
		x"72",	--3301
		x"62",	--3302
		x"79",	--3303
		x"77",	--3304
		x"6f",	--3305
		x"67",	--3306
		x"0a",	--3307
		x"25",	--3308
		x"20",	--3309
		x"64",	--3310
		x"0a",	--3311
		x"0d",	--3312
		x"3d",	--3313
		x"3d",	--3314
		x"3d",	--3315
		x"20",	--3316
		x"61",	--3317
		x"63",	--3318
		x"6c",	--3319
		x"4d",	--3320
		x"55",	--3321
		x"3d",	--3322
		x"3d",	--3323
		x"3d",	--3324
		x"0d",	--3325
		x"00",	--3326
		x"72",	--3327
		x"74",	--3328
		x"00",	--3329
		x"65",	--3330
		x"64",	--3331
		x"70",	--3332
		x"6d",	--3333
		x"65",	--3334
		x"63",	--3335
		x"64",	--3336
		x"72",	--3337
		x"62",	--3338
		x"6f",	--3339
		x"6c",	--3340
		x"61",	--3341
		x"65",	--3342
		x"00",	--3343
		x"0a",	--3344
		x"08",	--3345
		x"08",	--3346
		x"25",	--3347
		x"00",	--3348
		x"72",	--3349
		x"74",	--3350
		x"0a",	--3351
		x"00",	--3352
		x"6f",	--3353
		x"72",	--3354
		x"63",	--3355
		x"20",	--3356
		x"73",	--3357
		x"67",	--3358
		x"3a",	--3359
		x"0a",	--3360
		x"09",	--3361
		x"63",	--3362
		x"52",	--3363
		x"47",	--3364
		x"53",	--3365
		x"45",	--3366
		x"20",	--3367
		x"41",	--3368
		x"55",	--3369
		x"0d",	--3370
		x"00",	--3371
		x"6f",	--3372
		x"65",	--3373
		x"68",	--3374
		x"6e",	--3375
		x"20",	--3376
		x"65",	--3377
		x"74",	--3378
		x"74",	--3379
		x"72",	--3380
		x"69",	--3381
		x"6c",	--3382
		x"20",	--3383
		x"72",	--3384
		x"6e",	--3385
		x"0d",	--3386
		x"00",	--3387
		x"3d",	--3388
		x"64",	--3389
		x"76",	--3390
		x"25",	--3391
		x"0d",	--3392
		x"00",	--3393
		x"65",	--3394
		x"64",	--3395
		x"0d",	--3396
		x"09",	--3397
		x"63",	--3398
		x"52",	--3399
		x"47",	--3400
		x"53",	--3401
		x"45",	--3402
		x"0d",	--3403
		x"00",	--3404
		x"63",	--3405
		x"69",	--3406
		x"20",	--3407
		x"6f",	--3408
		x"20",	--3409
		x"20",	--3410
		x"75",	--3411
		x"62",	--3412
		x"72",	--3413
		x"0a",	--3414
		x"25",	--3415
		x"20",	--3416
		x"73",	--3417
		x"0a",	--3418
		x"25",	--3419
		x"3a",	--3420
		x"6e",	--3421
		x"20",	--3422
		x"75",	--3423
		x"68",	--3424
		x"63",	--3425
		x"6d",	--3426
		x"61",	--3427
		x"64",	--3428
		x"0a",	--3429
		x"00",	--3430
		x"eb",	--3431
		x"ea",	--3432
		x"ea",	--3433
		x"ea",	--3434
		x"ea",	--3435
		x"ea",	--3436
		x"ea",	--3437
		x"ea",	--3438
		x"ea",	--3439
		x"ea",	--3440
		x"ea",	--3441
		x"ea",	--3442
		x"ea",	--3443
		x"ea",	--3444
		x"ea",	--3445
		x"ea",	--3446
		x"ea",	--3447
		x"ea",	--3448
		x"ea",	--3449
		x"ea",	--3450
		x"ea",	--3451
		x"ea",	--3452
		x"ea",	--3453
		x"ea",	--3454
		x"ea",	--3455
		x"ea",	--3456
		x"ea",	--3457
		x"ea",	--3458
		x"ea",	--3459
		x"ea",	--3460
		x"ea",	--3461
		x"ea",	--3462
		x"ea",	--3463
		x"ea",	--3464
		x"ea",	--3465
		x"ea",	--3466
		x"ea",	--3467
		x"ea",	--3468
		x"ea",	--3469
		x"ea",	--3470
		x"ea",	--3471
		x"ea",	--3472
		x"ea",	--3473
		x"ea",	--3474
		x"ea",	--3475
		x"ea",	--3476
		x"ea",	--3477
		x"ea",	--3478
		x"ea",	--3479
		x"ea",	--3480
		x"ea",	--3481
		x"ea",	--3482
		x"ea",	--3483
		x"ea",	--3484
		x"ea",	--3485
		x"ea",	--3486
		x"ea",	--3487
		x"ea",	--3488
		x"ea",	--3489
		x"ea",	--3490
		x"ea",	--3491
		x"ea",	--3492
		x"ea",	--3493
		x"ea",	--3494
		x"ea",	--3495
		x"ea",	--3496
		x"ea",	--3497
		x"ea",	--3498
		x"ea",	--3499
		x"ea",	--3500
		x"ea",	--3501
		x"ea",	--3502
		x"ea",	--3503
		x"ea",	--3504
		x"ea",	--3505
		x"ea",	--3506
		x"ea",	--3507
		x"ea",	--3508
		x"ea",	--3509
		x"ea",	--3510
		x"ea",	--3511
		x"ea",	--3512
		x"ea",	--3513
		x"ea",	--3514
		x"31",	--3515
		x"33",	--3516
		x"35",	--3517
		x"37",	--3518
		x"39",	--3519
		x"62",	--3520
		x"64",	--3521
		x"66",	--3522
		x"00",	--3523
		x"00",	--3524
		x"00",	--3525
		x"00",	--3526
		x"00",	--3527
		x"01",	--3528
		x"02",	--3529
		x"03",	--3530
		x"03",	--3531
		x"04",	--3532
		x"04",	--3533
		x"04",	--3534
		x"04",	--3535
		x"05",	--3536
		x"05",	--3537
		x"05",	--3538
		x"05",	--3539
		x"05",	--3540
		x"05",	--3541
		x"05",	--3542
		x"05",	--3543
		x"06",	--3544
		x"06",	--3545
		x"06",	--3546
		x"06",	--3547
		x"06",	--3548
		x"06",	--3549
		x"06",	--3550
		x"06",	--3551
		x"06",	--3552
		x"06",	--3553
		x"06",	--3554
		x"06",	--3555
		x"06",	--3556
		x"06",	--3557
		x"06",	--3558
		x"06",	--3559
		x"07",	--3560
		x"07",	--3561
		x"07",	--3562
		x"07",	--3563
		x"07",	--3564
		x"07",	--3565
		x"07",	--3566
		x"07",	--3567
		x"07",	--3568
		x"07",	--3569
		x"07",	--3570
		x"07",	--3571
		x"07",	--3572
		x"07",	--3573
		x"07",	--3574
		x"07",	--3575
		x"07",	--3576
		x"07",	--3577
		x"07",	--3578
		x"07",	--3579
		x"07",	--3580
		x"07",	--3581
		x"07",	--3582
		x"07",	--3583
		x"07",	--3584
		x"07",	--3585
		x"07",	--3586
		x"07",	--3587
		x"07",	--3588
		x"07",	--3589
		x"07",	--3590
		x"07",	--3591
		x"08",	--3592
		x"08",	--3593
		x"08",	--3594
		x"08",	--3595
		x"08",	--3596
		x"08",	--3597
		x"08",	--3598
		x"08",	--3599
		x"08",	--3600
		x"08",	--3601
		x"08",	--3602
		x"08",	--3603
		x"08",	--3604
		x"08",	--3605
		x"08",	--3606
		x"08",	--3607
		x"08",	--3608
		x"08",	--3609
		x"08",	--3610
		x"08",	--3611
		x"08",	--3612
		x"08",	--3613
		x"08",	--3614
		x"08",	--3615
		x"08",	--3616
		x"08",	--3617
		x"08",	--3618
		x"08",	--3619
		x"08",	--3620
		x"08",	--3621
		x"08",	--3622
		x"08",	--3623
		x"08",	--3624
		x"08",	--3625
		x"08",	--3626
		x"08",	--3627
		x"08",	--3628
		x"08",	--3629
		x"08",	--3630
		x"08",	--3631
		x"08",	--3632
		x"08",	--3633
		x"08",	--3634
		x"08",	--3635
		x"08",	--3636
		x"08",	--3637
		x"08",	--3638
		x"08",	--3639
		x"08",	--3640
		x"08",	--3641
		x"08",	--3642
		x"08",	--3643
		x"08",	--3644
		x"08",	--3645
		x"08",	--3646
		x"08",	--3647
		x"08",	--3648
		x"08",	--3649
		x"08",	--3650
		x"08",	--3651
		x"08",	--3652
		x"08",	--3653
		x"08",	--3654
		x"08",	--3655
		x"65",	--3656
		x"70",	--3657
		x"00",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"eb",	--4087
		x"e7",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
