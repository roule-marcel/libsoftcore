library ieee;
use ieee.std_logic_1164.all;

library work;
use work.log2_pkg.all;

package ram16_pkg is
	type ram8_t is array (natural range <>) of std_logic_vector(7 downto 0);
	type position_t is ('h', 'l');

	component ram16 is
		generic (
			DEPTH : positive := 2048;
			INIT_FILE : string := "none"
		);
		port (
			clk : in std_logic;                                      -- Memory clock
			cen : in std_logic;                                      -- Memory chip enable (low active)
			addr : in std_logic_vector(log2ceil(DEPTH)-1 downto 0);  -- Memory address
			din : in std_logic_vector(15 downto 0);                  -- Memory data input
			wen : in std_logic_vector(1 downto 0);                   -- Memory write enable (low active)
			dout : out std_logic_vector(15 downto 0)                 -- Memory data output
		);
	end component ram16;
end package ram16_pkg;
