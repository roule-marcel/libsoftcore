library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"58",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"06",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"58",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"c0",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"52",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"58",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"06",	--29
		x"f9",	--30
		x"31",	--31
		x"be",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"80",	--41
		x"0f",	--42
		x"b0",	--43
		x"66",	--44
		x"b0",	--45
		x"ac",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"10",	--50
		x"b0",	--51
		x"2a",	--52
		x"21",	--53
		x"3d",	--54
		x"2d",	--55
		x"3e",	--56
		x"4a",	--57
		x"7f",	--58
		x"77",	--59
		x"b0",	--60
		x"dc",	--61
		x"3d",	--62
		x"33",	--63
		x"3e",	--64
		x"ea",	--65
		x"7f",	--66
		x"72",	--67
		x"b0",	--68
		x"dc",	--69
		x"3d",	--70
		x"38",	--71
		x"3e",	--72
		x"f2",	--73
		x"7f",	--74
		x"70",	--75
		x"b0",	--76
		x"dc",	--77
		x"3d",	--78
		x"3c",	--79
		x"3e",	--80
		x"ae",	--81
		x"7f",	--82
		x"65",	--83
		x"b0",	--84
		x"dc",	--85
		x"3d",	--86
		x"44",	--87
		x"3e",	--88
		x"bc",	--89
		x"7f",	--90
		x"62",	--91
		x"b0",	--92
		x"dc",	--93
		x"0f",	--94
		x"b0",	--95
		x"72",	--96
		x"2c",	--97
		x"3d",	--98
		x"20",	--99
		x"3e",	--100
		x"80",	--101
		x"0f",	--102
		x"3f",	--103
		x"0e",	--104
		x"b0",	--105
		x"82",	--106
		x"0f",	--107
		x"3f",	--108
		x"0e",	--109
		x"b0",	--110
		x"ca",	--111
		x"2c",	--112
		x"3d",	--113
		x"20",	--114
		x"3e",	--115
		x"88",	--116
		x"0f",	--117
		x"2f",	--118
		x"b0",	--119
		x"82",	--120
		x"0f",	--121
		x"2f",	--122
		x"b0",	--123
		x"ca",	--124
		x"0e",	--125
		x"2e",	--126
		x"0f",	--127
		x"3f",	--128
		x"0e",	--129
		x"b0",	--130
		x"e8",	--131
		x"3e",	--132
		x"98",	--133
		x"0f",	--134
		x"2f",	--135
		x"b0",	--136
		x"40",	--137
		x"3e",	--138
		x"9c",	--139
		x"0f",	--140
		x"b0",	--141
		x"40",	--142
		x"0e",	--143
		x"0f",	--144
		x"2f",	--145
		x"b0",	--146
		x"a4",	--147
		x"b0",	--148
		x"60",	--149
		x"0d",	--150
		x"3e",	--151
		x"d6",	--152
		x"1f",	--153
		x"b0",	--154
		x"70",	--155
		x"b0",	--156
		x"b6",	--157
		x"f2",	--158
		x"80",	--159
		x"19",	--160
		x"32",	--161
		x"0b",	--162
		x"b0",	--163
		x"74",	--164
		x"0f",	--165
		x"fc",	--166
		x"b0",	--167
		x"9c",	--168
		x"7f",	--169
		x"11",	--170
		x"7f",	--171
		x"0d",	--172
		x"17",	--173
		x"30",	--174
		x"4f",	--175
		x"b0",	--176
		x"2a",	--177
		x"21",	--178
		x"0e",	--179
		x"3e",	--180
		x"18",	--181
		x"5f",	--182
		x"18",	--183
		x"b0",	--184
		x"10",	--185
		x"0b",	--186
		x"e7",	--187
		x"0b",	--188
		x"e5",	--189
		x"3b",	--190
		x"30",	--191
		x"52",	--192
		x"b0",	--193
		x"2a",	--194
		x"21",	--195
		x"de",	--196
		x"3b",	--197
		x"28",	--198
		x"db",	--199
		x"4e",	--200
		x"8e",	--201
		x"0e",	--202
		x"30",	--203
		x"56",	--204
		x"81",	--205
		x"44",	--206
		x"b0",	--207
		x"2a",	--208
		x"21",	--209
		x"3e",	--210
		x"18",	--211
		x"0e",	--212
		x"0e",	--213
		x"1f",	--214
		x"40",	--215
		x"ce",	--216
		x"00",	--217
		x"1b",	--218
		x"c7",	--219
		x"30",	--220
		x"70",	--221
		x"b2",	--222
		x"00",	--223
		x"92",	--224
		x"a2",	--225
		x"94",	--226
		x"b2",	--227
		x"6d",	--228
		x"96",	--229
		x"30",	--230
		x"78",	--231
		x"b0",	--232
		x"2a",	--233
		x"92",	--234
		x"90",	--235
		x"b1",	--236
		x"96",	--237
		x"00",	--238
		x"b0",	--239
		x"2a",	--240
		x"21",	--241
		x"0f",	--242
		x"30",	--243
		x"82",	--244
		x"12",	--245
		x"82",	--246
		x"10",	--247
		x"30",	--248
		x"31",	--249
		x"ff",	--250
		x"20",	--251
		x"01",	--252
		x"39",	--253
		x"cf",	--254
		x"02",	--255
		x"36",	--256
		x"0d",	--257
		x"0e",	--258
		x"2e",	--259
		x"0f",	--260
		x"2f",	--261
		x"b0",	--262
		x"68",	--263
		x"81",	--264
		x"00",	--265
		x"40",	--266
		x"0d",	--267
		x"0e",	--268
		x"0f",	--269
		x"2f",	--270
		x"b0",	--271
		x"68",	--272
		x"81",	--273
		x"00",	--274
		x"37",	--275
		x"1e",	--276
		x"04",	--277
		x"0f",	--278
		x"b0",	--279
		x"8e",	--280
		x"0c",	--281
		x"3d",	--282
		x"c8",	--283
		x"b0",	--284
		x"5e",	--285
		x"0d",	--286
		x"0e",	--287
		x"1f",	--288
		x"12",	--289
		x"b0",	--290
		x"1e",	--291
		x"1e",	--292
		x"02",	--293
		x"0f",	--294
		x"b0",	--295
		x"8e",	--296
		x"0c",	--297
		x"3d",	--298
		x"c8",	--299
		x"b0",	--300
		x"5e",	--301
		x"0d",	--302
		x"0e",	--303
		x"1f",	--304
		x"10",	--305
		x"b0",	--306
		x"1e",	--307
		x"0f",	--308
		x"31",	--309
		x"30",	--310
		x"30",	--311
		x"af",	--312
		x"81",	--313
		x"08",	--314
		x"b0",	--315
		x"2a",	--316
		x"1f",	--317
		x"08",	--318
		x"6f",	--319
		x"8f",	--320
		x"81",	--321
		x"00",	--322
		x"30",	--323
		x"c0",	--324
		x"b0",	--325
		x"2a",	--326
		x"21",	--327
		x"3f",	--328
		x"31",	--329
		x"30",	--330
		x"30",	--331
		x"d1",	--332
		x"b0",	--333
		x"2a",	--334
		x"21",	--335
		x"3f",	--336
		x"e3",	--337
		x"82",	--338
		x"14",	--339
		x"82",	--340
		x"16",	--341
		x"30",	--342
		x"1f",	--343
		x"16",	--344
		x"2e",	--345
		x"1f",	--346
		x"14",	--347
		x"2f",	--348
		x"2e",	--349
		x"1e",	--350
		x"02",	--351
		x"2f",	--352
		x"1f",	--353
		x"02",	--354
		x"30",	--355
		x"f1",	--356
		x"b0",	--357
		x"2a",	--358
		x"31",	--359
		x"0a",	--360
		x"0f",	--361
		x"30",	--362
		x"1e",	--363
		x"06",	--364
		x"3e",	--365
		x"06",	--366
		x"0f",	--367
		x"0f",	--368
		x"10",	--369
		x"00",	--370
		x"c2",	--371
		x"19",	--372
		x"3e",	--373
		x"07",	--374
		x"03",	--375
		x"82",	--376
		x"06",	--377
		x"30",	--378
		x"1e",	--379
		x"82",	--380
		x"06",	--381
		x"30",	--382
		x"f2",	--383
		x"0e",	--384
		x"19",	--385
		x"f2",	--386
		x"f2",	--387
		x"0a",	--388
		x"19",	--389
		x"ee",	--390
		x"e2",	--391
		x"19",	--392
		x"eb",	--393
		x"f2",	--394
		x"0d",	--395
		x"19",	--396
		x"e7",	--397
		x"f2",	--398
		x"09",	--399
		x"19",	--400
		x"e3",	--401
		x"f2",	--402
		x"03",	--403
		x"19",	--404
		x"df",	--405
		x"f2",	--406
		x"07",	--407
		x"19",	--408
		x"db",	--409
		x"5e",	--410
		x"19",	--411
		x"4e",	--412
		x"0f",	--413
		x"03",	--414
		x"c2",	--415
		x"19",	--416
		x"30",	--417
		x"c2",	--418
		x"19",	--419
		x"30",	--420
		x"0b",	--421
		x"31",	--422
		x"fa",	--423
		x"0b",	--424
		x"30",	--425
		x"5a",	--426
		x"b0",	--427
		x"2a",	--428
		x"21",	--429
		x"fb",	--430
		x"20",	--431
		x"01",	--432
		x"2a",	--433
		x"cb",	--434
		x"02",	--435
		x"27",	--436
		x"0d",	--437
		x"0e",	--438
		x"2e",	--439
		x"0f",	--440
		x"2f",	--441
		x"b0",	--442
		x"68",	--443
		x"81",	--444
		x"00",	--445
		x"2f",	--446
		x"0d",	--447
		x"0e",	--448
		x"0f",	--449
		x"2f",	--450
		x"b0",	--451
		x"68",	--452
		x"81",	--453
		x"00",	--454
		x"26",	--455
		x"11",	--456
		x"04",	--457
		x"11",	--458
		x"08",	--459
		x"30",	--460
		x"a8",	--461
		x"b0",	--462
		x"2a",	--463
		x"31",	--464
		x"06",	--465
		x"1f",	--466
		x"04",	--467
		x"9f",	--468
		x"02",	--469
		x"00",	--470
		x"0f",	--471
		x"31",	--472
		x"06",	--473
		x"3b",	--474
		x"30",	--475
		x"30",	--476
		x"62",	--477
		x"b0",	--478
		x"2a",	--479
		x"6f",	--480
		x"8f",	--481
		x"81",	--482
		x"00",	--483
		x"30",	--484
		x"73",	--485
		x"b0",	--486
		x"2a",	--487
		x"21",	--488
		x"3f",	--489
		x"31",	--490
		x"06",	--491
		x"3b",	--492
		x"30",	--493
		x"30",	--494
		x"88",	--495
		x"b0",	--496
		x"2a",	--497
		x"21",	--498
		x"3f",	--499
		x"e3",	--500
		x"0b",	--501
		x"21",	--502
		x"0b",	--503
		x"30",	--504
		x"b4",	--505
		x"b0",	--506
		x"2a",	--507
		x"21",	--508
		x"fb",	--509
		x"20",	--510
		x"01",	--511
		x"1b",	--512
		x"cb",	--513
		x"02",	--514
		x"18",	--515
		x"0d",	--516
		x"0e",	--517
		x"2e",	--518
		x"0f",	--519
		x"2f",	--520
		x"b0",	--521
		x"68",	--522
		x"81",	--523
		x"00",	--524
		x"1f",	--525
		x"1f",	--526
		x"02",	--527
		x"2f",	--528
		x"0f",	--529
		x"30",	--530
		x"a8",	--531
		x"b0",	--532
		x"2a",	--533
		x"31",	--534
		x"06",	--535
		x"0f",	--536
		x"21",	--537
		x"3b",	--538
		x"30",	--539
		x"30",	--540
		x"62",	--541
		x"b0",	--542
		x"2a",	--543
		x"6f",	--544
		x"8f",	--545
		x"81",	--546
		x"00",	--547
		x"30",	--548
		x"bb",	--549
		x"b0",	--550
		x"2a",	--551
		x"21",	--552
		x"3f",	--553
		x"21",	--554
		x"3b",	--555
		x"30",	--556
		x"30",	--557
		x"88",	--558
		x"b0",	--559
		x"2a",	--560
		x"21",	--561
		x"3f",	--562
		x"e5",	--563
		x"0b",	--564
		x"0a",	--565
		x"09",	--566
		x"08",	--567
		x"07",	--568
		x"8f",	--569
		x"00",	--570
		x"8d",	--571
		x"00",	--572
		x"6c",	--573
		x"4c",	--574
		x"5f",	--575
		x"0b",	--576
		x"1b",	--577
		x"08",	--578
		x"0a",	--579
		x"07",	--580
		x"09",	--581
		x"18",	--582
		x"7a",	--583
		x"0a",	--584
		x"35",	--585
		x"2c",	--586
		x"0c",	--587
		x"0c",	--588
		x"0c",	--589
		x"0c",	--590
		x"8f",	--591
		x"00",	--592
		x"3c",	--593
		x"d0",	--594
		x"6a",	--595
		x"8a",	--596
		x"0c",	--597
		x"8f",	--598
		x"00",	--599
		x"17",	--600
		x"19",	--601
		x"0a",	--602
		x"08",	--603
		x"7c",	--604
		x"4c",	--605
		x"40",	--606
		x"7c",	--607
		x"78",	--608
		x"1b",	--609
		x"7c",	--610
		x"20",	--611
		x"43",	--612
		x"4a",	--613
		x"7a",	--614
		x"d0",	--615
		x"07",	--616
		x"dd",	--617
		x"7a",	--618
		x"0a",	--619
		x"46",	--620
		x"2a",	--621
		x"0a",	--622
		x"0c",	--623
		x"0c",	--624
		x"0c",	--625
		x"0c",	--626
		x"8f",	--627
		x"00",	--628
		x"3c",	--629
		x"d0",	--630
		x"68",	--631
		x"88",	--632
		x"0c",	--633
		x"8f",	--634
		x"00",	--635
		x"dc",	--636
		x"17",	--637
		x"da",	--638
		x"4a",	--639
		x"7a",	--640
		x"9f",	--641
		x"7a",	--642
		x"06",	--643
		x"0a",	--644
		x"2c",	--645
		x"0c",	--646
		x"0c",	--647
		x"0c",	--648
		x"0c",	--649
		x"8f",	--650
		x"00",	--651
		x"3c",	--652
		x"a9",	--653
		x"c4",	--654
		x"4a",	--655
		x"7a",	--656
		x"bf",	--657
		x"7a",	--658
		x"06",	--659
		x"1e",	--660
		x"2c",	--661
		x"0c",	--662
		x"0c",	--663
		x"0c",	--664
		x"0c",	--665
		x"8f",	--666
		x"00",	--667
		x"3c",	--668
		x"c9",	--669
		x"b4",	--670
		x"9d",	--671
		x"00",	--672
		x"0f",	--673
		x"37",	--674
		x"38",	--675
		x"39",	--676
		x"3a",	--677
		x"3b",	--678
		x"30",	--679
		x"9d",	--680
		x"00",	--681
		x"0f",	--682
		x"1f",	--683
		x"0f",	--684
		x"37",	--685
		x"38",	--686
		x"39",	--687
		x"3a",	--688
		x"3b",	--689
		x"30",	--690
		x"8c",	--691
		x"0c",	--692
		x"30",	--693
		x"ca",	--694
		x"b0",	--695
		x"2a",	--696
		x"21",	--697
		x"0f",	--698
		x"37",	--699
		x"38",	--700
		x"39",	--701
		x"3a",	--702
		x"3b",	--703
		x"30",	--704
		x"0b",	--705
		x"0a",	--706
		x"0b",	--707
		x"0a",	--708
		x"8f",	--709
		x"00",	--710
		x"8f",	--711
		x"02",	--712
		x"8f",	--713
		x"04",	--714
		x"0c",	--715
		x"0d",	--716
		x"3e",	--717
		x"00",	--718
		x"3f",	--719
		x"6e",	--720
		x"b0",	--721
		x"c2",	--722
		x"8b",	--723
		x"02",	--724
		x"02",	--725
		x"32",	--726
		x"03",	--727
		x"82",	--728
		x"32",	--729
		x"b2",	--730
		x"18",	--731
		x"38",	--732
		x"9b",	--733
		x"3a",	--734
		x"06",	--735
		x"32",	--736
		x"0f",	--737
		x"3a",	--738
		x"3b",	--739
		x"30",	--740
		x"0b",	--741
		x"09",	--742
		x"08",	--743
		x"8f",	--744
		x"06",	--745
		x"bf",	--746
		x"00",	--747
		x"08",	--748
		x"2b",	--749
		x"1e",	--750
		x"02",	--751
		x"0f",	--752
		x"b0",	--753
		x"8e",	--754
		x"0c",	--755
		x"3d",	--756
		x"00",	--757
		x"b0",	--758
		x"3a",	--759
		x"08",	--760
		x"09",	--761
		x"1e",	--762
		x"06",	--763
		x"0f",	--764
		x"b0",	--765
		x"8e",	--766
		x"0c",	--767
		x"0d",	--768
		x"0e",	--769
		x"0f",	--770
		x"b0",	--771
		x"ea",	--772
		x"b0",	--773
		x"ca",	--774
		x"8b",	--775
		x"04",	--776
		x"9b",	--777
		x"00",	--778
		x"38",	--779
		x"39",	--780
		x"3b",	--781
		x"30",	--782
		x"0b",	--783
		x"0a",	--784
		x"09",	--785
		x"0a",	--786
		x"0b",	--787
		x"8f",	--788
		x"06",	--789
		x"8f",	--790
		x"08",	--791
		x"29",	--792
		x"1e",	--793
		x"02",	--794
		x"0f",	--795
		x"b0",	--796
		x"8e",	--797
		x"0c",	--798
		x"0d",	--799
		x"0e",	--800
		x"0f",	--801
		x"b0",	--802
		x"3a",	--803
		x"0a",	--804
		x"0b",	--805
		x"1e",	--806
		x"06",	--807
		x"0f",	--808
		x"b0",	--809
		x"8e",	--810
		x"0c",	--811
		x"0d",	--812
		x"0e",	--813
		x"0f",	--814
		x"b0",	--815
		x"ea",	--816
		x"b0",	--817
		x"ca",	--818
		x"89",	--819
		x"04",	--820
		x"39",	--821
		x"3a",	--822
		x"3b",	--823
		x"30",	--824
		x"0b",	--825
		x"0a",	--826
		x"92",	--827
		x"08",	--828
		x"14",	--829
		x"3b",	--830
		x"1c",	--831
		x"0a",	--832
		x"2b",	--833
		x"5f",	--834
		x"fc",	--835
		x"8f",	--836
		x"0f",	--837
		x"30",	--838
		x"df",	--839
		x"b0",	--840
		x"2a",	--841
		x"31",	--842
		x"06",	--843
		x"1a",	--844
		x"3b",	--845
		x"06",	--846
		x"1a",	--847
		x"08",	--848
		x"ef",	--849
		x"0f",	--850
		x"3a",	--851
		x"3b",	--852
		x"30",	--853
		x"1e",	--854
		x"08",	--855
		x"3e",	--856
		x"20",	--857
		x"12",	--858
		x"0f",	--859
		x"0f",	--860
		x"0f",	--861
		x"0f",	--862
		x"3f",	--863
		x"18",	--864
		x"ff",	--865
		x"68",	--866
		x"00",	--867
		x"bf",	--868
		x"72",	--869
		x"02",	--870
		x"bf",	--871
		x"00",	--872
		x"04",	--873
		x"1e",	--874
		x"82",	--875
		x"08",	--876
		x"30",	--877
		x"0b",	--878
		x"1b",	--879
		x"08",	--880
		x"3b",	--881
		x"20",	--882
		x"12",	--883
		x"0c",	--884
		x"0c",	--885
		x"0c",	--886
		x"0c",	--887
		x"3c",	--888
		x"18",	--889
		x"cc",	--890
		x"00",	--891
		x"8c",	--892
		x"02",	--893
		x"8c",	--894
		x"04",	--895
		x"1b",	--896
		x"82",	--897
		x"08",	--898
		x"0f",	--899
		x"3b",	--900
		x"30",	--901
		x"3f",	--902
		x"fc",	--903
		x"0b",	--904
		x"1b",	--905
		x"08",	--906
		x"1b",	--907
		x"0f",	--908
		x"5f",	--909
		x"18",	--910
		x"14",	--911
		x"3d",	--912
		x"1e",	--913
		x"0c",	--914
		x"05",	--915
		x"3d",	--916
		x"06",	--917
		x"cd",	--918
		x"fa",	--919
		x"0c",	--920
		x"1c",	--921
		x"0c",	--922
		x"f8",	--923
		x"30",	--924
		x"e7",	--925
		x"b0",	--926
		x"2a",	--927
		x"21",	--928
		x"3f",	--929
		x"3b",	--930
		x"30",	--931
		x"0c",	--932
		x"0d",	--933
		x"0d",	--934
		x"0c",	--935
		x"0c",	--936
		x"3c",	--937
		x"18",	--938
		x"0f",	--939
		x"9c",	--940
		x"02",	--941
		x"3b",	--942
		x"30",	--943
		x"b2",	--944
		x"d2",	--945
		x"60",	--946
		x"b2",	--947
		x"b8",	--948
		x"72",	--949
		x"0f",	--950
		x"30",	--951
		x"0b",	--952
		x"0a",	--953
		x"0a",	--954
		x"1f",	--955
		x"0a",	--956
		x"3f",	--957
		x"20",	--958
		x"19",	--959
		x"0b",	--960
		x"0b",	--961
		x"0c",	--962
		x"0c",	--963
		x"0c",	--964
		x"0c",	--965
		x"3c",	--966
		x"d8",	--967
		x"8c",	--968
		x"00",	--969
		x"8c",	--970
		x"02",	--971
		x"8c",	--972
		x"04",	--973
		x"8c",	--974
		x"06",	--975
		x"8c",	--976
		x"08",	--977
		x"0e",	--978
		x"1e",	--979
		x"82",	--980
		x"0a",	--981
		x"3a",	--982
		x"3b",	--983
		x"30",	--984
		x"3f",	--985
		x"fb",	--986
		x"0f",	--987
		x"0e",	--988
		x"0e",	--989
		x"0e",	--990
		x"0e",	--991
		x"9e",	--992
		x"d8",	--993
		x"0f",	--994
		x"30",	--995
		x"0f",	--996
		x"0e",	--997
		x"0e",	--998
		x"0e",	--999
		x"0e",	--1000
		x"8e",	--1001
		x"d8",	--1002
		x"0f",	--1003
		x"30",	--1004
		x"0f",	--1005
		x"0e",	--1006
		x"0d",	--1007
		x"0c",	--1008
		x"0b",	--1009
		x"0a",	--1010
		x"92",	--1011
		x"0a",	--1012
		x"20",	--1013
		x"3b",	--1014
		x"da",	--1015
		x"0a",	--1016
		x"09",	--1017
		x"1f",	--1018
		x"8b",	--1019
		x"00",	--1020
		x"1a",	--1021
		x"3b",	--1022
		x"0a",	--1023
		x"1a",	--1024
		x"0a",	--1025
		x"13",	--1026
		x"8b",	--1027
		x"fe",	--1028
		x"f7",	--1029
		x"2f",	--1030
		x"1f",	--1031
		x"02",	--1032
		x"f0",	--1033
		x"8b",	--1034
		x"00",	--1035
		x"1f",	--1036
		x"06",	--1037
		x"9b",	--1038
		x"04",	--1039
		x"1a",	--1040
		x"3b",	--1041
		x"0a",	--1042
		x"1a",	--1043
		x"0a",	--1044
		x"ed",	--1045
		x"b2",	--1046
		x"fe",	--1047
		x"60",	--1048
		x"3a",	--1049
		x"3b",	--1050
		x"3c",	--1051
		x"3d",	--1052
		x"3e",	--1053
		x"3f",	--1054
		x"00",	--1055
		x"8f",	--1056
		x"00",	--1057
		x"0f",	--1058
		x"30",	--1059
		x"2f",	--1060
		x"2f",	--1061
		x"30",	--1062
		x"5e",	--1063
		x"81",	--1064
		x"3e",	--1065
		x"fc",	--1066
		x"c2",	--1067
		x"84",	--1068
		x"0f",	--1069
		x"30",	--1070
		x"3f",	--1071
		x"0f",	--1072
		x"5f",	--1073
		x"a6",	--1074
		x"8f",	--1075
		x"b0",	--1076
		x"4e",	--1077
		x"30",	--1078
		x"0b",	--1079
		x"0b",	--1080
		x"0e",	--1081
		x"0e",	--1082
		x"0e",	--1083
		x"0e",	--1084
		x"0e",	--1085
		x"0f",	--1086
		x"b0",	--1087
		x"5e",	--1088
		x"0f",	--1089
		x"b0",	--1090
		x"5e",	--1091
		x"3b",	--1092
		x"30",	--1093
		x"0b",	--1094
		x"0a",	--1095
		x"0a",	--1096
		x"3b",	--1097
		x"07",	--1098
		x"0e",	--1099
		x"4d",	--1100
		x"7d",	--1101
		x"0f",	--1102
		x"03",	--1103
		x"0e",	--1104
		x"7d",	--1105
		x"fd",	--1106
		x"1e",	--1107
		x"0a",	--1108
		x"3f",	--1109
		x"31",	--1110
		x"b0",	--1111
		x"4e",	--1112
		x"3b",	--1113
		x"3b",	--1114
		x"ef",	--1115
		x"3a",	--1116
		x"3b",	--1117
		x"30",	--1118
		x"3f",	--1119
		x"30",	--1120
		x"f5",	--1121
		x"0b",	--1122
		x"0b",	--1123
		x"0e",	--1124
		x"8e",	--1125
		x"8e",	--1126
		x"0f",	--1127
		x"b0",	--1128
		x"6e",	--1129
		x"0f",	--1130
		x"b0",	--1131
		x"6e",	--1132
		x"3b",	--1133
		x"30",	--1134
		x"0b",	--1135
		x"0a",	--1136
		x"0a",	--1137
		x"0b",	--1138
		x"0d",	--1139
		x"8d",	--1140
		x"8d",	--1141
		x"0f",	--1142
		x"b0",	--1143
		x"6e",	--1144
		x"0f",	--1145
		x"b0",	--1146
		x"6e",	--1147
		x"0c",	--1148
		x"0d",	--1149
		x"8d",	--1150
		x"8c",	--1151
		x"4d",	--1152
		x"0d",	--1153
		x"0f",	--1154
		x"b0",	--1155
		x"6e",	--1156
		x"0f",	--1157
		x"b0",	--1158
		x"6e",	--1159
		x"3a",	--1160
		x"3b",	--1161
		x"30",	--1162
		x"0b",	--1163
		x"0a",	--1164
		x"09",	--1165
		x"0a",	--1166
		x"0e",	--1167
		x"19",	--1168
		x"09",	--1169
		x"39",	--1170
		x"0b",	--1171
		x"0d",	--1172
		x"0d",	--1173
		x"6f",	--1174
		x"8f",	--1175
		x"b0",	--1176
		x"6e",	--1177
		x"0b",	--1178
		x"0e",	--1179
		x"1b",	--1180
		x"3b",	--1181
		x"07",	--1182
		x"05",	--1183
		x"3f",	--1184
		x"20",	--1185
		x"b0",	--1186
		x"4e",	--1187
		x"ef",	--1188
		x"3f",	--1189
		x"3a",	--1190
		x"b0",	--1191
		x"4e",	--1192
		x"ea",	--1193
		x"39",	--1194
		x"3a",	--1195
		x"3b",	--1196
		x"30",	--1197
		x"0b",	--1198
		x"0a",	--1199
		x"09",	--1200
		x"0a",	--1201
		x"0e",	--1202
		x"17",	--1203
		x"09",	--1204
		x"39",	--1205
		x"0b",	--1206
		x"6f",	--1207
		x"8f",	--1208
		x"b0",	--1209
		x"5e",	--1210
		x"0b",	--1211
		x"0e",	--1212
		x"1b",	--1213
		x"3b",	--1214
		x"07",	--1215
		x"f6",	--1216
		x"3f",	--1217
		x"20",	--1218
		x"b0",	--1219
		x"4e",	--1220
		x"6f",	--1221
		x"8f",	--1222
		x"b0",	--1223
		x"5e",	--1224
		x"0b",	--1225
		x"f2",	--1226
		x"39",	--1227
		x"3a",	--1228
		x"3b",	--1229
		x"30",	--1230
		x"0b",	--1231
		x"0a",	--1232
		x"09",	--1233
		x"31",	--1234
		x"ec",	--1235
		x"0b",	--1236
		x"0f",	--1237
		x"34",	--1238
		x"3b",	--1239
		x"0a",	--1240
		x"38",	--1241
		x"09",	--1242
		x"0a",	--1243
		x"0a",	--1244
		x"3e",	--1245
		x"0a",	--1246
		x"0f",	--1247
		x"b0",	--1248
		x"ba",	--1249
		x"7f",	--1250
		x"30",	--1251
		x"ca",	--1252
		x"00",	--1253
		x"19",	--1254
		x"3e",	--1255
		x"0a",	--1256
		x"0f",	--1257
		x"b0",	--1258
		x"88",	--1259
		x"0b",	--1260
		x"3f",	--1261
		x"0a",	--1262
		x"eb",	--1263
		x"0a",	--1264
		x"1a",	--1265
		x"09",	--1266
		x"3e",	--1267
		x"0a",	--1268
		x"0f",	--1269
		x"b0",	--1270
		x"ba",	--1271
		x"7f",	--1272
		x"30",	--1273
		x"c9",	--1274
		x"00",	--1275
		x"3a",	--1276
		x"0f",	--1277
		x"0f",	--1278
		x"6f",	--1279
		x"8f",	--1280
		x"b0",	--1281
		x"4e",	--1282
		x"0a",	--1283
		x"f7",	--1284
		x"31",	--1285
		x"14",	--1286
		x"39",	--1287
		x"3a",	--1288
		x"3b",	--1289
		x"30",	--1290
		x"3f",	--1291
		x"2d",	--1292
		x"b0",	--1293
		x"4e",	--1294
		x"3b",	--1295
		x"1b",	--1296
		x"c5",	--1297
		x"1a",	--1298
		x"09",	--1299
		x"dd",	--1300
		x"0b",	--1301
		x"0a",	--1302
		x"09",	--1303
		x"0b",	--1304
		x"3b",	--1305
		x"39",	--1306
		x"6f",	--1307
		x"4f",	--1308
		x"0b",	--1309
		x"1a",	--1310
		x"8f",	--1311
		x"b0",	--1312
		x"4e",	--1313
		x"0a",	--1314
		x"09",	--1315
		x"19",	--1316
		x"5f",	--1317
		x"01",	--1318
		x"4f",	--1319
		x"10",	--1320
		x"7f",	--1321
		x"25",	--1322
		x"f3",	--1323
		x"0a",	--1324
		x"1a",	--1325
		x"5f",	--1326
		x"01",	--1327
		x"7f",	--1328
		x"db",	--1329
		x"7f",	--1330
		x"54",	--1331
		x"ee",	--1332
		x"4f",	--1333
		x"0f",	--1334
		x"10",	--1335
		x"fe",	--1336
		x"39",	--1337
		x"3a",	--1338
		x"3b",	--1339
		x"30",	--1340
		x"09",	--1341
		x"29",	--1342
		x"1e",	--1343
		x"02",	--1344
		x"2f",	--1345
		x"b0",	--1346
		x"16",	--1347
		x"0b",	--1348
		x"dd",	--1349
		x"09",	--1350
		x"29",	--1351
		x"2f",	--1352
		x"b0",	--1353
		x"c4",	--1354
		x"0b",	--1355
		x"d6",	--1356
		x"0f",	--1357
		x"2b",	--1358
		x"29",	--1359
		x"6f",	--1360
		x"4f",	--1361
		x"d0",	--1362
		x"19",	--1363
		x"8f",	--1364
		x"b0",	--1365
		x"4e",	--1366
		x"7f",	--1367
		x"4f",	--1368
		x"fa",	--1369
		x"c8",	--1370
		x"09",	--1371
		x"29",	--1372
		x"1e",	--1373
		x"02",	--1374
		x"2f",	--1375
		x"b0",	--1376
		x"5c",	--1377
		x"0b",	--1378
		x"bf",	--1379
		x"09",	--1380
		x"29",	--1381
		x"2e",	--1382
		x"0f",	--1383
		x"8f",	--1384
		x"8f",	--1385
		x"8f",	--1386
		x"8f",	--1387
		x"b0",	--1388
		x"de",	--1389
		x"0b",	--1390
		x"b3",	--1391
		x"09",	--1392
		x"29",	--1393
		x"2f",	--1394
		x"b0",	--1395
		x"9e",	--1396
		x"0b",	--1397
		x"ac",	--1398
		x"09",	--1399
		x"29",	--1400
		x"2f",	--1401
		x"b0",	--1402
		x"4e",	--1403
		x"0b",	--1404
		x"a5",	--1405
		x"09",	--1406
		x"29",	--1407
		x"2f",	--1408
		x"b0",	--1409
		x"6e",	--1410
		x"0b",	--1411
		x"9e",	--1412
		x"09",	--1413
		x"29",	--1414
		x"2f",	--1415
		x"b0",	--1416
		x"8c",	--1417
		x"0b",	--1418
		x"97",	--1419
		x"3f",	--1420
		x"25",	--1421
		x"b0",	--1422
		x"4e",	--1423
		x"92",	--1424
		x"0f",	--1425
		x"0e",	--1426
		x"1f",	--1427
		x"0c",	--1428
		x"df",	--1429
		x"85",	--1430
		x"18",	--1431
		x"1f",	--1432
		x"0c",	--1433
		x"3f",	--1434
		x"3f",	--1435
		x"13",	--1436
		x"92",	--1437
		x"0c",	--1438
		x"1e",	--1439
		x"0c",	--1440
		x"1f",	--1441
		x"0e",	--1442
		x"0e",	--1443
		x"02",	--1444
		x"92",	--1445
		x"0e",	--1446
		x"f2",	--1447
		x"10",	--1448
		x"81",	--1449
		x"3e",	--1450
		x"3f",	--1451
		x"b1",	--1452
		x"f0",	--1453
		x"00",	--1454
		x"00",	--1455
		x"82",	--1456
		x"0c",	--1457
		x"ec",	--1458
		x"b2",	--1459
		x"c3",	--1460
		x"82",	--1461
		x"f2",	--1462
		x"11",	--1463
		x"80",	--1464
		x"30",	--1465
		x"1e",	--1466
		x"0c",	--1467
		x"1f",	--1468
		x"0e",	--1469
		x"0e",	--1470
		x"05",	--1471
		x"1f",	--1472
		x"0c",	--1473
		x"1f",	--1474
		x"0e",	--1475
		x"30",	--1476
		x"1d",	--1477
		x"0c",	--1478
		x"1e",	--1479
		x"0e",	--1480
		x"3f",	--1481
		x"40",	--1482
		x"0f",	--1483
		x"0f",	--1484
		x"30",	--1485
		x"1f",	--1486
		x"0e",	--1487
		x"5f",	--1488
		x"18",	--1489
		x"1d",	--1490
		x"0e",	--1491
		x"1e",	--1492
		x"0c",	--1493
		x"0d",	--1494
		x"0b",	--1495
		x"1e",	--1496
		x"0e",	--1497
		x"3e",	--1498
		x"3f",	--1499
		x"03",	--1500
		x"82",	--1501
		x"0e",	--1502
		x"30",	--1503
		x"92",	--1504
		x"0e",	--1505
		x"30",	--1506
		x"4f",	--1507
		x"30",	--1508
		x"0b",	--1509
		x"0a",	--1510
		x"0a",	--1511
		x"0b",	--1512
		x"0c",	--1513
		x"3d",	--1514
		x"00",	--1515
		x"b0",	--1516
		x"ae",	--1517
		x"0f",	--1518
		x"07",	--1519
		x"0e",	--1520
		x"0f",	--1521
		x"b0",	--1522
		x"fe",	--1523
		x"3a",	--1524
		x"3b",	--1525
		x"30",	--1526
		x"0c",	--1527
		x"3d",	--1528
		x"00",	--1529
		x"0e",	--1530
		x"0f",	--1531
		x"b0",	--1532
		x"ea",	--1533
		x"b0",	--1534
		x"fe",	--1535
		x"0e",	--1536
		x"3f",	--1537
		x"00",	--1538
		x"3a",	--1539
		x"3b",	--1540
		x"30",	--1541
		x"0b",	--1542
		x"0a",	--1543
		x"09",	--1544
		x"08",	--1545
		x"07",	--1546
		x"06",	--1547
		x"05",	--1548
		x"04",	--1549
		x"31",	--1550
		x"fa",	--1551
		x"08",	--1552
		x"6b",	--1553
		x"6b",	--1554
		x"67",	--1555
		x"6c",	--1556
		x"6c",	--1557
		x"e9",	--1558
		x"6b",	--1559
		x"02",	--1560
		x"30",	--1561
		x"8c",	--1562
		x"6c",	--1563
		x"e3",	--1564
		x"6c",	--1565
		x"bb",	--1566
		x"6b",	--1567
		x"df",	--1568
		x"91",	--1569
		x"02",	--1570
		x"00",	--1571
		x"1b",	--1572
		x"02",	--1573
		x"14",	--1574
		x"04",	--1575
		x"15",	--1576
		x"06",	--1577
		x"16",	--1578
		x"04",	--1579
		x"17",	--1580
		x"06",	--1581
		x"2c",	--1582
		x"0c",	--1583
		x"09",	--1584
		x"0c",	--1585
		x"bf",	--1586
		x"39",	--1587
		x"20",	--1588
		x"50",	--1589
		x"1c",	--1590
		x"d7",	--1591
		x"81",	--1592
		x"02",	--1593
		x"81",	--1594
		x"04",	--1595
		x"4c",	--1596
		x"7c",	--1597
		x"1f",	--1598
		x"0b",	--1599
		x"0a",	--1600
		x"0b",	--1601
		x"12",	--1602
		x"0b",	--1603
		x"0a",	--1604
		x"7c",	--1605
		x"fb",	--1606
		x"81",	--1607
		x"02",	--1608
		x"81",	--1609
		x"04",	--1610
		x"1c",	--1611
		x"0d",	--1612
		x"79",	--1613
		x"1f",	--1614
		x"04",	--1615
		x"0c",	--1616
		x"0d",	--1617
		x"79",	--1618
		x"fc",	--1619
		x"3c",	--1620
		x"3d",	--1621
		x"0c",	--1622
		x"0d",	--1623
		x"1a",	--1624
		x"0b",	--1625
		x"0c",	--1626
		x"02",	--1627
		x"0d",	--1628
		x"e5",	--1629
		x"16",	--1630
		x"02",	--1631
		x"17",	--1632
		x"04",	--1633
		x"06",	--1634
		x"07",	--1635
		x"5f",	--1636
		x"01",	--1637
		x"5f",	--1638
		x"01",	--1639
		x"28",	--1640
		x"c8",	--1641
		x"01",	--1642
		x"a8",	--1643
		x"02",	--1644
		x"0e",	--1645
		x"0f",	--1646
		x"0e",	--1647
		x"0f",	--1648
		x"88",	--1649
		x"04",	--1650
		x"88",	--1651
		x"06",	--1652
		x"f8",	--1653
		x"03",	--1654
		x"00",	--1655
		x"0f",	--1656
		x"4d",	--1657
		x"0f",	--1658
		x"31",	--1659
		x"06",	--1660
		x"34",	--1661
		x"35",	--1662
		x"36",	--1663
		x"37",	--1664
		x"38",	--1665
		x"39",	--1666
		x"3a",	--1667
		x"3b",	--1668
		x"30",	--1669
		x"2b",	--1670
		x"67",	--1671
		x"81",	--1672
		x"00",	--1673
		x"04",	--1674
		x"05",	--1675
		x"5f",	--1676
		x"01",	--1677
		x"5f",	--1678
		x"01",	--1679
		x"d8",	--1680
		x"4f",	--1681
		x"68",	--1682
		x"0e",	--1683
		x"0f",	--1684
		x"0e",	--1685
		x"0f",	--1686
		x"0f",	--1687
		x"69",	--1688
		x"c8",	--1689
		x"01",	--1690
		x"a8",	--1691
		x"02",	--1692
		x"88",	--1693
		x"04",	--1694
		x"88",	--1695
		x"06",	--1696
		x"0c",	--1697
		x"0d",	--1698
		x"3c",	--1699
		x"3d",	--1700
		x"3d",	--1701
		x"ff",	--1702
		x"05",	--1703
		x"3d",	--1704
		x"00",	--1705
		x"17",	--1706
		x"3c",	--1707
		x"15",	--1708
		x"1b",	--1709
		x"02",	--1710
		x"3b",	--1711
		x"0e",	--1712
		x"0f",	--1713
		x"0a",	--1714
		x"3b",	--1715
		x"0c",	--1716
		x"0d",	--1717
		x"3c",	--1718
		x"3d",	--1719
		x"3d",	--1720
		x"ff",	--1721
		x"f5",	--1722
		x"3c",	--1723
		x"88",	--1724
		x"04",	--1725
		x"88",	--1726
		x"06",	--1727
		x"88",	--1728
		x"02",	--1729
		x"f8",	--1730
		x"03",	--1731
		x"00",	--1732
		x"0f",	--1733
		x"b3",	--1734
		x"0c",	--1735
		x"0d",	--1736
		x"1c",	--1737
		x"0d",	--1738
		x"12",	--1739
		x"0f",	--1740
		x"0e",	--1741
		x"0a",	--1742
		x"0b",	--1743
		x"0a",	--1744
		x"0b",	--1745
		x"88",	--1746
		x"04",	--1747
		x"88",	--1748
		x"06",	--1749
		x"98",	--1750
		x"02",	--1751
		x"0f",	--1752
		x"a1",	--1753
		x"6b",	--1754
		x"9f",	--1755
		x"ad",	--1756
		x"00",	--1757
		x"9d",	--1758
		x"02",	--1759
		x"02",	--1760
		x"9d",	--1761
		x"04",	--1762
		x"04",	--1763
		x"9d",	--1764
		x"06",	--1765
		x"06",	--1766
		x"5e",	--1767
		x"01",	--1768
		x"5e",	--1769
		x"01",	--1770
		x"cd",	--1771
		x"01",	--1772
		x"0f",	--1773
		x"8c",	--1774
		x"06",	--1775
		x"07",	--1776
		x"9a",	--1777
		x"39",	--1778
		x"19",	--1779
		x"39",	--1780
		x"20",	--1781
		x"8f",	--1782
		x"3e",	--1783
		x"3c",	--1784
		x"b6",	--1785
		x"c1",	--1786
		x"0e",	--1787
		x"0f",	--1788
		x"0e",	--1789
		x"0f",	--1790
		x"97",	--1791
		x"0f",	--1792
		x"79",	--1793
		x"d8",	--1794
		x"01",	--1795
		x"a8",	--1796
		x"02",	--1797
		x"3e",	--1798
		x"3f",	--1799
		x"1e",	--1800
		x"0f",	--1801
		x"88",	--1802
		x"04",	--1803
		x"88",	--1804
		x"06",	--1805
		x"92",	--1806
		x"0c",	--1807
		x"7b",	--1808
		x"81",	--1809
		x"00",	--1810
		x"81",	--1811
		x"02",	--1812
		x"81",	--1813
		x"04",	--1814
		x"4d",	--1815
		x"7d",	--1816
		x"1f",	--1817
		x"0c",	--1818
		x"4b",	--1819
		x"0c",	--1820
		x"0d",	--1821
		x"12",	--1822
		x"0d",	--1823
		x"0c",	--1824
		x"7b",	--1825
		x"fb",	--1826
		x"81",	--1827
		x"02",	--1828
		x"81",	--1829
		x"04",	--1830
		x"1c",	--1831
		x"0d",	--1832
		x"79",	--1833
		x"1f",	--1834
		x"04",	--1835
		x"0c",	--1836
		x"0d",	--1837
		x"79",	--1838
		x"fc",	--1839
		x"3c",	--1840
		x"3d",	--1841
		x"0c",	--1842
		x"0d",	--1843
		x"1a",	--1844
		x"0b",	--1845
		x"0c",	--1846
		x"04",	--1847
		x"0d",	--1848
		x"02",	--1849
		x"0a",	--1850
		x"0b",	--1851
		x"14",	--1852
		x"02",	--1853
		x"15",	--1854
		x"04",	--1855
		x"04",	--1856
		x"05",	--1857
		x"49",	--1858
		x"0a",	--1859
		x"0b",	--1860
		x"18",	--1861
		x"6c",	--1862
		x"33",	--1863
		x"df",	--1864
		x"01",	--1865
		x"01",	--1866
		x"2f",	--1867
		x"3f",	--1868
		x"b8",	--1869
		x"2c",	--1870
		x"31",	--1871
		x"e0",	--1872
		x"81",	--1873
		x"04",	--1874
		x"81",	--1875
		x"06",	--1876
		x"81",	--1877
		x"00",	--1878
		x"81",	--1879
		x"02",	--1880
		x"0e",	--1881
		x"3e",	--1882
		x"18",	--1883
		x"0f",	--1884
		x"2f",	--1885
		x"b0",	--1886
		x"c0",	--1887
		x"0e",	--1888
		x"3e",	--1889
		x"10",	--1890
		x"0f",	--1891
		x"b0",	--1892
		x"c0",	--1893
		x"0d",	--1894
		x"3d",	--1895
		x"0e",	--1896
		x"3e",	--1897
		x"10",	--1898
		x"0f",	--1899
		x"3f",	--1900
		x"18",	--1901
		x"b0",	--1902
		x"0c",	--1903
		x"b0",	--1904
		x"e2",	--1905
		x"31",	--1906
		x"20",	--1907
		x"30",	--1908
		x"31",	--1909
		x"e0",	--1910
		x"81",	--1911
		x"04",	--1912
		x"81",	--1913
		x"06",	--1914
		x"81",	--1915
		x"00",	--1916
		x"81",	--1917
		x"02",	--1918
		x"0e",	--1919
		x"3e",	--1920
		x"18",	--1921
		x"0f",	--1922
		x"2f",	--1923
		x"b0",	--1924
		x"c0",	--1925
		x"0e",	--1926
		x"3e",	--1927
		x"10",	--1928
		x"0f",	--1929
		x"b0",	--1930
		x"c0",	--1931
		x"d1",	--1932
		x"11",	--1933
		x"0d",	--1934
		x"3d",	--1935
		x"0e",	--1936
		x"3e",	--1937
		x"10",	--1938
		x"0f",	--1939
		x"3f",	--1940
		x"18",	--1941
		x"b0",	--1942
		x"0c",	--1943
		x"b0",	--1944
		x"e2",	--1945
		x"31",	--1946
		x"20",	--1947
		x"30",	--1948
		x"0b",	--1949
		x"0a",	--1950
		x"09",	--1951
		x"08",	--1952
		x"07",	--1953
		x"06",	--1954
		x"05",	--1955
		x"04",	--1956
		x"31",	--1957
		x"dc",	--1958
		x"81",	--1959
		x"04",	--1960
		x"81",	--1961
		x"06",	--1962
		x"81",	--1963
		x"00",	--1964
		x"81",	--1965
		x"02",	--1966
		x"0e",	--1967
		x"3e",	--1968
		x"18",	--1969
		x"0f",	--1970
		x"2f",	--1971
		x"b0",	--1972
		x"c0",	--1973
		x"0e",	--1974
		x"3e",	--1975
		x"10",	--1976
		x"0f",	--1977
		x"b0",	--1978
		x"c0",	--1979
		x"5f",	--1980
		x"18",	--1981
		x"6f",	--1982
		x"b6",	--1983
		x"5e",	--1984
		x"10",	--1985
		x"6e",	--1986
		x"d9",	--1987
		x"6f",	--1988
		x"ae",	--1989
		x"6e",	--1990
		x"e2",	--1991
		x"6f",	--1992
		x"ac",	--1993
		x"6e",	--1994
		x"d1",	--1995
		x"14",	--1996
		x"1c",	--1997
		x"15",	--1998
		x"1e",	--1999
		x"18",	--2000
		x"14",	--2001
		x"19",	--2002
		x"16",	--2003
		x"3c",	--2004
		x"20",	--2005
		x"0e",	--2006
		x"0f",	--2007
		x"06",	--2008
		x"07",	--2009
		x"81",	--2010
		x"20",	--2011
		x"81",	--2012
		x"22",	--2013
		x"0a",	--2014
		x"0b",	--2015
		x"81",	--2016
		x"20",	--2017
		x"08",	--2018
		x"08",	--2019
		x"09",	--2020
		x"12",	--2021
		x"05",	--2022
		x"04",	--2023
		x"b1",	--2024
		x"20",	--2025
		x"19",	--2026
		x"14",	--2027
		x"0d",	--2028
		x"0a",	--2029
		x"0b",	--2030
		x"0e",	--2031
		x"0f",	--2032
		x"1c",	--2033
		x"0d",	--2034
		x"0b",	--2035
		x"03",	--2036
		x"0b",	--2037
		x"0c",	--2038
		x"0d",	--2039
		x"0e",	--2040
		x"0f",	--2041
		x"06",	--2042
		x"07",	--2043
		x"09",	--2044
		x"e5",	--2045
		x"16",	--2046
		x"07",	--2047
		x"e2",	--2048
		x"0a",	--2049
		x"f5",	--2050
		x"f2",	--2051
		x"81",	--2052
		x"20",	--2053
		x"81",	--2054
		x"22",	--2055
		x"0c",	--2056
		x"1a",	--2057
		x"1a",	--2058
		x"1a",	--2059
		x"12",	--2060
		x"06",	--2061
		x"26",	--2062
		x"81",	--2063
		x"0a",	--2064
		x"5d",	--2065
		x"d1",	--2066
		x"11",	--2067
		x"19",	--2068
		x"83",	--2069
		x"c1",	--2070
		x"09",	--2071
		x"0c",	--2072
		x"3c",	--2073
		x"3f",	--2074
		x"00",	--2075
		x"18",	--2076
		x"1d",	--2077
		x"0a",	--2078
		x"3d",	--2079
		x"1a",	--2080
		x"20",	--2081
		x"1b",	--2082
		x"22",	--2083
		x"0c",	--2084
		x"0e",	--2085
		x"0f",	--2086
		x"0b",	--2087
		x"2a",	--2088
		x"0a",	--2089
		x"0b",	--2090
		x"3d",	--2091
		x"3f",	--2092
		x"00",	--2093
		x"f5",	--2094
		x"81",	--2095
		x"20",	--2096
		x"81",	--2097
		x"22",	--2098
		x"81",	--2099
		x"0a",	--2100
		x"0c",	--2101
		x"0d",	--2102
		x"3c",	--2103
		x"7f",	--2104
		x"0d",	--2105
		x"3c",	--2106
		x"40",	--2107
		x"44",	--2108
		x"81",	--2109
		x"0c",	--2110
		x"81",	--2111
		x"0e",	--2112
		x"f1",	--2113
		x"03",	--2114
		x"08",	--2115
		x"0f",	--2116
		x"3f",	--2117
		x"b0",	--2118
		x"e2",	--2119
		x"31",	--2120
		x"24",	--2121
		x"34",	--2122
		x"35",	--2123
		x"36",	--2124
		x"37",	--2125
		x"38",	--2126
		x"39",	--2127
		x"3a",	--2128
		x"3b",	--2129
		x"30",	--2130
		x"1e",	--2131
		x"0f",	--2132
		x"d3",	--2133
		x"3a",	--2134
		x"03",	--2135
		x"08",	--2136
		x"1e",	--2137
		x"10",	--2138
		x"1c",	--2139
		x"20",	--2140
		x"1d",	--2141
		x"22",	--2142
		x"12",	--2143
		x"0d",	--2144
		x"0c",	--2145
		x"06",	--2146
		x"07",	--2147
		x"06",	--2148
		x"37",	--2149
		x"00",	--2150
		x"81",	--2151
		x"20",	--2152
		x"81",	--2153
		x"22",	--2154
		x"12",	--2155
		x"0f",	--2156
		x"0e",	--2157
		x"1a",	--2158
		x"0f",	--2159
		x"e7",	--2160
		x"81",	--2161
		x"0a",	--2162
		x"a6",	--2163
		x"6e",	--2164
		x"36",	--2165
		x"5f",	--2166
		x"d1",	--2167
		x"11",	--2168
		x"19",	--2169
		x"20",	--2170
		x"c1",	--2171
		x"19",	--2172
		x"0f",	--2173
		x"3f",	--2174
		x"18",	--2175
		x"c5",	--2176
		x"0d",	--2177
		x"ba",	--2178
		x"0c",	--2179
		x"0d",	--2180
		x"3c",	--2181
		x"80",	--2182
		x"0d",	--2183
		x"0c",	--2184
		x"b3",	--2185
		x"0d",	--2186
		x"b1",	--2187
		x"81",	--2188
		x"20",	--2189
		x"03",	--2190
		x"81",	--2191
		x"22",	--2192
		x"ab",	--2193
		x"3e",	--2194
		x"40",	--2195
		x"0f",	--2196
		x"3e",	--2197
		x"80",	--2198
		x"3f",	--2199
		x"a4",	--2200
		x"4d",	--2201
		x"7b",	--2202
		x"4f",	--2203
		x"de",	--2204
		x"5f",	--2205
		x"d1",	--2206
		x"11",	--2207
		x"19",	--2208
		x"06",	--2209
		x"c1",	--2210
		x"11",	--2211
		x"0f",	--2212
		x"3f",	--2213
		x"10",	--2214
		x"9e",	--2215
		x"4f",	--2216
		x"f8",	--2217
		x"6f",	--2218
		x"f1",	--2219
		x"3f",	--2220
		x"b8",	--2221
		x"97",	--2222
		x"0b",	--2223
		x"0a",	--2224
		x"09",	--2225
		x"08",	--2226
		x"07",	--2227
		x"31",	--2228
		x"e8",	--2229
		x"81",	--2230
		x"04",	--2231
		x"81",	--2232
		x"06",	--2233
		x"81",	--2234
		x"00",	--2235
		x"81",	--2236
		x"02",	--2237
		x"0e",	--2238
		x"3e",	--2239
		x"10",	--2240
		x"0f",	--2241
		x"2f",	--2242
		x"b0",	--2243
		x"c0",	--2244
		x"0e",	--2245
		x"3e",	--2246
		x"0f",	--2247
		x"b0",	--2248
		x"c0",	--2249
		x"5f",	--2250
		x"10",	--2251
		x"6f",	--2252
		x"5d",	--2253
		x"5e",	--2254
		x"08",	--2255
		x"6e",	--2256
		x"82",	--2257
		x"d1",	--2258
		x"09",	--2259
		x"11",	--2260
		x"6f",	--2261
		x"58",	--2262
		x"6f",	--2263
		x"56",	--2264
		x"6e",	--2265
		x"6f",	--2266
		x"6e",	--2267
		x"4c",	--2268
		x"1d",	--2269
		x"12",	--2270
		x"1d",	--2271
		x"0a",	--2272
		x"81",	--2273
		x"12",	--2274
		x"1e",	--2275
		x"14",	--2276
		x"1f",	--2277
		x"16",	--2278
		x"18",	--2279
		x"0c",	--2280
		x"19",	--2281
		x"0e",	--2282
		x"0f",	--2283
		x"1e",	--2284
		x"0e",	--2285
		x"0f",	--2286
		x"3d",	--2287
		x"81",	--2288
		x"12",	--2289
		x"37",	--2290
		x"1f",	--2291
		x"0c",	--2292
		x"3d",	--2293
		x"00",	--2294
		x"0a",	--2295
		x"0b",	--2296
		x"0b",	--2297
		x"0a",	--2298
		x"0b",	--2299
		x"0e",	--2300
		x"0f",	--2301
		x"12",	--2302
		x"0d",	--2303
		x"0c",	--2304
		x"0e",	--2305
		x"0f",	--2306
		x"37",	--2307
		x"0b",	--2308
		x"0f",	--2309
		x"f7",	--2310
		x"f2",	--2311
		x"0e",	--2312
		x"f4",	--2313
		x"ef",	--2314
		x"09",	--2315
		x"e5",	--2316
		x"0e",	--2317
		x"e3",	--2318
		x"dd",	--2319
		x"0c",	--2320
		x"0d",	--2321
		x"3c",	--2322
		x"7f",	--2323
		x"0d",	--2324
		x"3c",	--2325
		x"40",	--2326
		x"1c",	--2327
		x"81",	--2328
		x"14",	--2329
		x"81",	--2330
		x"16",	--2331
		x"0f",	--2332
		x"3f",	--2333
		x"10",	--2334
		x"b0",	--2335
		x"e2",	--2336
		x"31",	--2337
		x"18",	--2338
		x"37",	--2339
		x"38",	--2340
		x"39",	--2341
		x"3a",	--2342
		x"3b",	--2343
		x"30",	--2344
		x"e1",	--2345
		x"10",	--2346
		x"0f",	--2347
		x"3f",	--2348
		x"10",	--2349
		x"f0",	--2350
		x"4f",	--2351
		x"fa",	--2352
		x"3f",	--2353
		x"b8",	--2354
		x"eb",	--2355
		x"0d",	--2356
		x"e2",	--2357
		x"0c",	--2358
		x"0d",	--2359
		x"3c",	--2360
		x"80",	--2361
		x"0d",	--2362
		x"0c",	--2363
		x"db",	--2364
		x"0d",	--2365
		x"d9",	--2366
		x"0e",	--2367
		x"02",	--2368
		x"0f",	--2369
		x"d5",	--2370
		x"3a",	--2371
		x"40",	--2372
		x"0b",	--2373
		x"3a",	--2374
		x"80",	--2375
		x"3b",	--2376
		x"ce",	--2377
		x"81",	--2378
		x"14",	--2379
		x"81",	--2380
		x"16",	--2381
		x"81",	--2382
		x"12",	--2383
		x"0f",	--2384
		x"3f",	--2385
		x"10",	--2386
		x"cb",	--2387
		x"0f",	--2388
		x"3f",	--2389
		x"c8",	--2390
		x"31",	--2391
		x"e8",	--2392
		x"81",	--2393
		x"04",	--2394
		x"81",	--2395
		x"06",	--2396
		x"81",	--2397
		x"00",	--2398
		x"81",	--2399
		x"02",	--2400
		x"0e",	--2401
		x"3e",	--2402
		x"10",	--2403
		x"0f",	--2404
		x"2f",	--2405
		x"b0",	--2406
		x"c0",	--2407
		x"0e",	--2408
		x"3e",	--2409
		x"0f",	--2410
		x"b0",	--2411
		x"c0",	--2412
		x"e1",	--2413
		x"10",	--2414
		x"0d",	--2415
		x"e1",	--2416
		x"08",	--2417
		x"0a",	--2418
		x"0e",	--2419
		x"3e",	--2420
		x"0f",	--2421
		x"3f",	--2422
		x"10",	--2423
		x"b0",	--2424
		x"e4",	--2425
		x"31",	--2426
		x"18",	--2427
		x"30",	--2428
		x"3f",	--2429
		x"fb",	--2430
		x"31",	--2431
		x"f4",	--2432
		x"81",	--2433
		x"00",	--2434
		x"81",	--2435
		x"02",	--2436
		x"0e",	--2437
		x"2e",	--2438
		x"0f",	--2439
		x"b0",	--2440
		x"c0",	--2441
		x"5f",	--2442
		x"04",	--2443
		x"6f",	--2444
		x"28",	--2445
		x"27",	--2446
		x"6f",	--2447
		x"07",	--2448
		x"1d",	--2449
		x"06",	--2450
		x"0d",	--2451
		x"21",	--2452
		x"3d",	--2453
		x"1f",	--2454
		x"09",	--2455
		x"c1",	--2456
		x"05",	--2457
		x"26",	--2458
		x"3e",	--2459
		x"3f",	--2460
		x"ff",	--2461
		x"31",	--2462
		x"0c",	--2463
		x"30",	--2464
		x"1e",	--2465
		x"08",	--2466
		x"1f",	--2467
		x"0a",	--2468
		x"3c",	--2469
		x"1e",	--2470
		x"4c",	--2471
		x"4d",	--2472
		x"7d",	--2473
		x"1f",	--2474
		x"0f",	--2475
		x"c1",	--2476
		x"05",	--2477
		x"ef",	--2478
		x"3e",	--2479
		x"3f",	--2480
		x"1e",	--2481
		x"0f",	--2482
		x"31",	--2483
		x"0c",	--2484
		x"30",	--2485
		x"0e",	--2486
		x"0f",	--2487
		x"31",	--2488
		x"0c",	--2489
		x"30",	--2490
		x"12",	--2491
		x"0f",	--2492
		x"0e",	--2493
		x"7d",	--2494
		x"fb",	--2495
		x"eb",	--2496
		x"0e",	--2497
		x"3f",	--2498
		x"00",	--2499
		x"31",	--2500
		x"0c",	--2501
		x"30",	--2502
		x"0b",	--2503
		x"0a",	--2504
		x"09",	--2505
		x"08",	--2506
		x"31",	--2507
		x"0a",	--2508
		x"0b",	--2509
		x"c1",	--2510
		x"01",	--2511
		x"0e",	--2512
		x"0d",	--2513
		x"0b",	--2514
		x"0b",	--2515
		x"e1",	--2516
		x"00",	--2517
		x"0f",	--2518
		x"b0",	--2519
		x"e2",	--2520
		x"31",	--2521
		x"38",	--2522
		x"39",	--2523
		x"3a",	--2524
		x"3b",	--2525
		x"30",	--2526
		x"f1",	--2527
		x"03",	--2528
		x"00",	--2529
		x"b1",	--2530
		x"1e",	--2531
		x"02",	--2532
		x"81",	--2533
		x"04",	--2534
		x"81",	--2535
		x"06",	--2536
		x"0e",	--2537
		x"0f",	--2538
		x"b0",	--2539
		x"70",	--2540
		x"3f",	--2541
		x"0f",	--2542
		x"18",	--2543
		x"e5",	--2544
		x"81",	--2545
		x"04",	--2546
		x"81",	--2547
		x"06",	--2548
		x"4e",	--2549
		x"7e",	--2550
		x"1f",	--2551
		x"06",	--2552
		x"3e",	--2553
		x"1e",	--2554
		x"0e",	--2555
		x"81",	--2556
		x"02",	--2557
		x"d7",	--2558
		x"91",	--2559
		x"04",	--2560
		x"04",	--2561
		x"91",	--2562
		x"06",	--2563
		x"06",	--2564
		x"7e",	--2565
		x"f8",	--2566
		x"f1",	--2567
		x"0e",	--2568
		x"3e",	--2569
		x"1e",	--2570
		x"1c",	--2571
		x"0d",	--2572
		x"48",	--2573
		x"78",	--2574
		x"1f",	--2575
		x"04",	--2576
		x"0c",	--2577
		x"0d",	--2578
		x"78",	--2579
		x"fc",	--2580
		x"3c",	--2581
		x"3d",	--2582
		x"0c",	--2583
		x"0d",	--2584
		x"18",	--2585
		x"09",	--2586
		x"0c",	--2587
		x"04",	--2588
		x"0d",	--2589
		x"02",	--2590
		x"08",	--2591
		x"09",	--2592
		x"7e",	--2593
		x"1f",	--2594
		x"0e",	--2595
		x"0d",	--2596
		x"0e",	--2597
		x"0d",	--2598
		x"0e",	--2599
		x"81",	--2600
		x"04",	--2601
		x"81",	--2602
		x"06",	--2603
		x"3e",	--2604
		x"1e",	--2605
		x"0e",	--2606
		x"81",	--2607
		x"02",	--2608
		x"a4",	--2609
		x"12",	--2610
		x"0b",	--2611
		x"0a",	--2612
		x"7e",	--2613
		x"fb",	--2614
		x"ec",	--2615
		x"0b",	--2616
		x"0a",	--2617
		x"09",	--2618
		x"1f",	--2619
		x"17",	--2620
		x"3e",	--2621
		x"00",	--2622
		x"2c",	--2623
		x"3a",	--2624
		x"18",	--2625
		x"0b",	--2626
		x"39",	--2627
		x"0c",	--2628
		x"0d",	--2629
		x"4f",	--2630
		x"4f",	--2631
		x"17",	--2632
		x"3c",	--2633
		x"c0",	--2634
		x"6e",	--2635
		x"0f",	--2636
		x"0a",	--2637
		x"0b",	--2638
		x"0f",	--2639
		x"39",	--2640
		x"3a",	--2641
		x"3b",	--2642
		x"30",	--2643
		x"3f",	--2644
		x"00",	--2645
		x"0f",	--2646
		x"3a",	--2647
		x"0b",	--2648
		x"39",	--2649
		x"18",	--2650
		x"0c",	--2651
		x"0d",	--2652
		x"4f",	--2653
		x"4f",	--2654
		x"e9",	--2655
		x"12",	--2656
		x"0d",	--2657
		x"0c",	--2658
		x"7f",	--2659
		x"fb",	--2660
		x"e3",	--2661
		x"3a",	--2662
		x"10",	--2663
		x"0b",	--2664
		x"39",	--2665
		x"10",	--2666
		x"ef",	--2667
		x"3a",	--2668
		x"20",	--2669
		x"0b",	--2670
		x"09",	--2671
		x"ea",	--2672
		x"0b",	--2673
		x"0a",	--2674
		x"09",	--2675
		x"08",	--2676
		x"07",	--2677
		x"0d",	--2678
		x"1e",	--2679
		x"04",	--2680
		x"1f",	--2681
		x"06",	--2682
		x"5a",	--2683
		x"01",	--2684
		x"6c",	--2685
		x"6c",	--2686
		x"70",	--2687
		x"6c",	--2688
		x"6a",	--2689
		x"6c",	--2690
		x"36",	--2691
		x"0e",	--2692
		x"32",	--2693
		x"1b",	--2694
		x"02",	--2695
		x"3b",	--2696
		x"82",	--2697
		x"6d",	--2698
		x"3b",	--2699
		x"80",	--2700
		x"5e",	--2701
		x"0c",	--2702
		x"0d",	--2703
		x"3c",	--2704
		x"7f",	--2705
		x"0d",	--2706
		x"3c",	--2707
		x"40",	--2708
		x"40",	--2709
		x"3e",	--2710
		x"3f",	--2711
		x"0f",	--2712
		x"0f",	--2713
		x"4a",	--2714
		x"0d",	--2715
		x"3d",	--2716
		x"7f",	--2717
		x"12",	--2718
		x"0f",	--2719
		x"0e",	--2720
		x"12",	--2721
		x"0f",	--2722
		x"0e",	--2723
		x"12",	--2724
		x"0f",	--2725
		x"0e",	--2726
		x"12",	--2727
		x"0f",	--2728
		x"0e",	--2729
		x"12",	--2730
		x"0f",	--2731
		x"0e",	--2732
		x"12",	--2733
		x"0f",	--2734
		x"0e",	--2735
		x"12",	--2736
		x"0f",	--2737
		x"0e",	--2738
		x"3e",	--2739
		x"3f",	--2740
		x"7f",	--2741
		x"4d",	--2742
		x"05",	--2743
		x"0f",	--2744
		x"cc",	--2745
		x"4d",	--2746
		x"0e",	--2747
		x"0f",	--2748
		x"4d",	--2749
		x"0d",	--2750
		x"0d",	--2751
		x"0d",	--2752
		x"0d",	--2753
		x"0d",	--2754
		x"0d",	--2755
		x"0d",	--2756
		x"0c",	--2757
		x"3c",	--2758
		x"7f",	--2759
		x"0c",	--2760
		x"4f",	--2761
		x"0f",	--2762
		x"0f",	--2763
		x"0f",	--2764
		x"0d",	--2765
		x"0d",	--2766
		x"0f",	--2767
		x"37",	--2768
		x"38",	--2769
		x"39",	--2770
		x"3a",	--2771
		x"3b",	--2772
		x"30",	--2773
		x"0d",	--2774
		x"be",	--2775
		x"0c",	--2776
		x"0d",	--2777
		x"3c",	--2778
		x"80",	--2779
		x"0d",	--2780
		x"0c",	--2781
		x"02",	--2782
		x"0d",	--2783
		x"b8",	--2784
		x"3e",	--2785
		x"40",	--2786
		x"0f",	--2787
		x"b4",	--2788
		x"12",	--2789
		x"0f",	--2790
		x"0e",	--2791
		x"0d",	--2792
		x"3d",	--2793
		x"80",	--2794
		x"b2",	--2795
		x"7d",	--2796
		x"0e",	--2797
		x"0f",	--2798
		x"cd",	--2799
		x"0e",	--2800
		x"3f",	--2801
		x"10",	--2802
		x"3e",	--2803
		x"3f",	--2804
		x"7f",	--2805
		x"7d",	--2806
		x"c5",	--2807
		x"37",	--2808
		x"82",	--2809
		x"07",	--2810
		x"37",	--2811
		x"1a",	--2812
		x"4f",	--2813
		x"0c",	--2814
		x"0d",	--2815
		x"4b",	--2816
		x"7b",	--2817
		x"1f",	--2818
		x"05",	--2819
		x"12",	--2820
		x"0d",	--2821
		x"0c",	--2822
		x"7b",	--2823
		x"fb",	--2824
		x"18",	--2825
		x"09",	--2826
		x"77",	--2827
		x"1f",	--2828
		x"04",	--2829
		x"08",	--2830
		x"09",	--2831
		x"77",	--2832
		x"fc",	--2833
		x"38",	--2834
		x"39",	--2835
		x"08",	--2836
		x"09",	--2837
		x"1e",	--2838
		x"0f",	--2839
		x"08",	--2840
		x"04",	--2841
		x"09",	--2842
		x"02",	--2843
		x"0e",	--2844
		x"0f",	--2845
		x"08",	--2846
		x"09",	--2847
		x"08",	--2848
		x"09",	--2849
		x"0e",	--2850
		x"0f",	--2851
		x"3e",	--2852
		x"7f",	--2853
		x"0f",	--2854
		x"3e",	--2855
		x"40",	--2856
		x"26",	--2857
		x"38",	--2858
		x"3f",	--2859
		x"09",	--2860
		x"0e",	--2861
		x"0f",	--2862
		x"12",	--2863
		x"0f",	--2864
		x"0e",	--2865
		x"12",	--2866
		x"0f",	--2867
		x"0e",	--2868
		x"12",	--2869
		x"0f",	--2870
		x"0e",	--2871
		x"12",	--2872
		x"0f",	--2873
		x"0e",	--2874
		x"12",	--2875
		x"0f",	--2876
		x"0e",	--2877
		x"12",	--2878
		x"0f",	--2879
		x"0e",	--2880
		x"12",	--2881
		x"0f",	--2882
		x"0e",	--2883
		x"3e",	--2884
		x"3f",	--2885
		x"7f",	--2886
		x"5d",	--2887
		x"39",	--2888
		x"00",	--2889
		x"72",	--2890
		x"4d",	--2891
		x"70",	--2892
		x"08",	--2893
		x"09",	--2894
		x"da",	--2895
		x"0f",	--2896
		x"d8",	--2897
		x"0e",	--2898
		x"0f",	--2899
		x"3e",	--2900
		x"80",	--2901
		x"0f",	--2902
		x"0e",	--2903
		x"04",	--2904
		x"38",	--2905
		x"40",	--2906
		x"09",	--2907
		x"d0",	--2908
		x"0f",	--2909
		x"ce",	--2910
		x"f9",	--2911
		x"0b",	--2912
		x"0a",	--2913
		x"2a",	--2914
		x"5b",	--2915
		x"02",	--2916
		x"3b",	--2917
		x"7f",	--2918
		x"1d",	--2919
		x"02",	--2920
		x"12",	--2921
		x"0d",	--2922
		x"12",	--2923
		x"0d",	--2924
		x"12",	--2925
		x"0d",	--2926
		x"12",	--2927
		x"0d",	--2928
		x"12",	--2929
		x"0d",	--2930
		x"12",	--2931
		x"0d",	--2932
		x"12",	--2933
		x"0d",	--2934
		x"4d",	--2935
		x"5f",	--2936
		x"03",	--2937
		x"3f",	--2938
		x"80",	--2939
		x"0f",	--2940
		x"0f",	--2941
		x"ce",	--2942
		x"01",	--2943
		x"0d",	--2944
		x"2d",	--2945
		x"0a",	--2946
		x"51",	--2947
		x"be",	--2948
		x"82",	--2949
		x"02",	--2950
		x"0c",	--2951
		x"0d",	--2952
		x"0c",	--2953
		x"0d",	--2954
		x"0c",	--2955
		x"0d",	--2956
		x"0c",	--2957
		x"0d",	--2958
		x"0c",	--2959
		x"0d",	--2960
		x"0c",	--2961
		x"0d",	--2962
		x"0c",	--2963
		x"0d",	--2964
		x"0c",	--2965
		x"0d",	--2966
		x"fe",	--2967
		x"03",	--2968
		x"00",	--2969
		x"3d",	--2970
		x"00",	--2971
		x"0b",	--2972
		x"3f",	--2973
		x"81",	--2974
		x"0c",	--2975
		x"0d",	--2976
		x"0a",	--2977
		x"3f",	--2978
		x"3d",	--2979
		x"00",	--2980
		x"f9",	--2981
		x"8e",	--2982
		x"02",	--2983
		x"8e",	--2984
		x"04",	--2985
		x"8e",	--2986
		x"06",	--2987
		x"3a",	--2988
		x"3b",	--2989
		x"30",	--2990
		x"3d",	--2991
		x"ff",	--2992
		x"2a",	--2993
		x"3d",	--2994
		x"81",	--2995
		x"8e",	--2996
		x"02",	--2997
		x"fe",	--2998
		x"03",	--2999
		x"00",	--3000
		x"0c",	--3001
		x"0d",	--3002
		x"0c",	--3003
		x"0d",	--3004
		x"0c",	--3005
		x"0d",	--3006
		x"0c",	--3007
		x"0d",	--3008
		x"0c",	--3009
		x"0d",	--3010
		x"0c",	--3011
		x"0d",	--3012
		x"0c",	--3013
		x"0d",	--3014
		x"0c",	--3015
		x"0d",	--3016
		x"0a",	--3017
		x"0b",	--3018
		x"0a",	--3019
		x"3b",	--3020
		x"00",	--3021
		x"8e",	--3022
		x"04",	--3023
		x"8e",	--3024
		x"06",	--3025
		x"3a",	--3026
		x"3b",	--3027
		x"30",	--3028
		x"0b",	--3029
		x"ad",	--3030
		x"ee",	--3031
		x"00",	--3032
		x"3a",	--3033
		x"3b",	--3034
		x"30",	--3035
		x"0a",	--3036
		x"0c",	--3037
		x"0c",	--3038
		x"0d",	--3039
		x"0c",	--3040
		x"3d",	--3041
		x"10",	--3042
		x"0c",	--3043
		x"02",	--3044
		x"0d",	--3045
		x"08",	--3046
		x"de",	--3047
		x"00",	--3048
		x"e4",	--3049
		x"0b",	--3050
		x"f2",	--3051
		x"ee",	--3052
		x"00",	--3053
		x"e3",	--3054
		x"ce",	--3055
		x"00",	--3056
		x"dc",	--3057
		x"0b",	--3058
		x"6d",	--3059
		x"6d",	--3060
		x"12",	--3061
		x"6c",	--3062
		x"6c",	--3063
		x"0f",	--3064
		x"6d",	--3065
		x"41",	--3066
		x"6c",	--3067
		x"11",	--3068
		x"6d",	--3069
		x"0d",	--3070
		x"6c",	--3071
		x"14",	--3072
		x"5d",	--3073
		x"01",	--3074
		x"5d",	--3075
		x"01",	--3076
		x"14",	--3077
		x"4d",	--3078
		x"09",	--3079
		x"1e",	--3080
		x"0f",	--3081
		x"3b",	--3082
		x"30",	--3083
		x"6c",	--3084
		x"28",	--3085
		x"ce",	--3086
		x"01",	--3087
		x"f7",	--3088
		x"3e",	--3089
		x"0f",	--3090
		x"3b",	--3091
		x"30",	--3092
		x"cf",	--3093
		x"01",	--3094
		x"f0",	--3095
		x"3e",	--3096
		x"f8",	--3097
		x"1b",	--3098
		x"02",	--3099
		x"1c",	--3100
		x"02",	--3101
		x"0c",	--3102
		x"e6",	--3103
		x"0b",	--3104
		x"16",	--3105
		x"1b",	--3106
		x"04",	--3107
		x"1f",	--3108
		x"06",	--3109
		x"1c",	--3110
		x"04",	--3111
		x"1e",	--3112
		x"06",	--3113
		x"0e",	--3114
		x"da",	--3115
		x"0f",	--3116
		x"02",	--3117
		x"0c",	--3118
		x"d6",	--3119
		x"0f",	--3120
		x"06",	--3121
		x"0e",	--3122
		x"02",	--3123
		x"0b",	--3124
		x"02",	--3125
		x"0e",	--3126
		x"d1",	--3127
		x"4d",	--3128
		x"ce",	--3129
		x"3e",	--3130
		x"d6",	--3131
		x"6c",	--3132
		x"d7",	--3133
		x"5e",	--3134
		x"01",	--3135
		x"5f",	--3136
		x"01",	--3137
		x"0e",	--3138
		x"c5",	--3139
		x"0d",	--3140
		x"0f",	--3141
		x"04",	--3142
		x"3d",	--3143
		x"03",	--3144
		x"3f",	--3145
		x"1f",	--3146
		x"0e",	--3147
		x"03",	--3148
		x"5d",	--3149
		x"3e",	--3150
		x"1e",	--3151
		x"0d",	--3152
		x"b0",	--3153
		x"0e",	--3154
		x"3d",	--3155
		x"6d",	--3156
		x"02",	--3157
		x"3e",	--3158
		x"1e",	--3159
		x"5d",	--3160
		x"02",	--3161
		x"3f",	--3162
		x"1f",	--3163
		x"30",	--3164
		x"b0",	--3165
		x"88",	--3166
		x"0f",	--3167
		x"30",	--3168
		x"0b",	--3169
		x"0b",	--3170
		x"0f",	--3171
		x"06",	--3172
		x"3b",	--3173
		x"03",	--3174
		x"3e",	--3175
		x"3f",	--3176
		x"1e",	--3177
		x"0f",	--3178
		x"0d",	--3179
		x"05",	--3180
		x"5b",	--3181
		x"3c",	--3182
		x"3d",	--3183
		x"1c",	--3184
		x"0d",	--3185
		x"b0",	--3186
		x"30",	--3187
		x"6b",	--3188
		x"04",	--3189
		x"3c",	--3190
		x"3d",	--3191
		x"1c",	--3192
		x"0d",	--3193
		x"5b",	--3194
		x"04",	--3195
		x"3e",	--3196
		x"3f",	--3197
		x"1e",	--3198
		x"0f",	--3199
		x"3b",	--3200
		x"30",	--3201
		x"b0",	--3202
		x"c2",	--3203
		x"0e",	--3204
		x"0f",	--3205
		x"30",	--3206
		x"7c",	--3207
		x"10",	--3208
		x"0d",	--3209
		x"0e",	--3210
		x"0f",	--3211
		x"0e",	--3212
		x"0e",	--3213
		x"02",	--3214
		x"0e",	--3215
		x"1f",	--3216
		x"1c",	--3217
		x"f8",	--3218
		x"30",	--3219
		x"b0",	--3220
		x"0e",	--3221
		x"0f",	--3222
		x"30",	--3223
		x"0b",	--3224
		x"0a",	--3225
		x"09",	--3226
		x"79",	--3227
		x"20",	--3228
		x"0a",	--3229
		x"0b",	--3230
		x"0c",	--3231
		x"0d",	--3232
		x"0e",	--3233
		x"0f",	--3234
		x"0c",	--3235
		x"0d",	--3236
		x"0d",	--3237
		x"06",	--3238
		x"02",	--3239
		x"0c",	--3240
		x"03",	--3241
		x"0c",	--3242
		x"0d",	--3243
		x"1e",	--3244
		x"19",	--3245
		x"f2",	--3246
		x"39",	--3247
		x"3a",	--3248
		x"3b",	--3249
		x"30",	--3250
		x"b0",	--3251
		x"30",	--3252
		x"0e",	--3253
		x"0f",	--3254
		x"30",	--3255
		x"00",	--3256
		x"32",	--3257
		x"f0",	--3258
		x"fd",	--3259
		x"57",	--3260
		x"69",	--3261
		x"69",	--3262
		x"67",	--3263
		x"66",	--3264
		x"72",	--3265
		x"61",	--3266
		x"6e",	--3267
		x"77",	--3268
		x"2e",	--3269
		x"69",	--3270
		x"20",	--3271
		x"69",	--3272
		x"65",	--3273
		x"0a",	--3274
		x"57",	--3275
		x"20",	--3276
		x"68",	--3277
		x"75",	--3278
		x"64",	--3279
		x"6e",	--3280
		x"74",	--3281
		x"73",	--3282
		x"65",	--3283
		x"74",	--3284
		x"61",	--3285
		x"0d",	--3286
		x"00",	--3287
		x"6f",	--3288
		x"72",	--3289
		x"63",	--3290
		x"20",	--3291
		x"73",	--3292
		x"67",	--3293
		x"3a",	--3294
		x"0a",	--3295
		x"09",	--3296
		x"63",	--3297
		x"4c",	--3298
		x"46",	--3299
		x"20",	--3300
		x"49",	--3301
		x"48",	--3302
		x"0d",	--3303
		x"00",	--3304
		x"6f",	--3305
		x"65",	--3306
		x"68",	--3307
		x"6e",	--3308
		x"20",	--3309
		x"65",	--3310
		x"74",	--3311
		x"74",	--3312
		x"72",	--3313
		x"69",	--3314
		x"6c",	--3315
		x"20",	--3316
		x"72",	--3317
		x"6e",	--3318
		x"0d",	--3319
		x"00",	--3320
		x"77",	--3321
		x"25",	--3322
		x"20",	--3323
		x"77",	--3324
		x"25",	--3325
		x"0d",	--3326
		x"00",	--3327
		x"e6",	--3328
		x"0e",	--3329
		x"14",	--3330
		x"1c",	--3331
		x"24",	--3332
		x"2c",	--3333
		x"fe",	--3334
		x"06",	--3335
		x"0d",	--3336
		x"3d",	--3337
		x"3d",	--3338
		x"3d",	--3339
		x"20",	--3340
		x"61",	--3341
		x"63",	--3342
		x"6c",	--3343
		x"4d",	--3344
		x"55",	--3345
		x"3d",	--3346
		x"3d",	--3347
		x"3d",	--3348
		x"0d",	--3349
		x"00",	--3350
		x"72",	--3351
		x"74",	--3352
		x"00",	--3353
		x"65",	--3354
		x"64",	--3355
		x"70",	--3356
		x"6d",	--3357
		x"65",	--3358
		x"63",	--3359
		x"64",	--3360
		x"72",	--3361
		x"62",	--3362
		x"6f",	--3363
		x"6c",	--3364
		x"61",	--3365
		x"65",	--3366
		x"00",	--3367
		x"0a",	--3368
		x"08",	--3369
		x"08",	--3370
		x"25",	--3371
		x"00",	--3372
		x"77",	--3373
		x"69",	--3374
		x"65",	--3375
		x"0d",	--3376
		x"63",	--3377
		x"72",	--3378
		x"65",	--3379
		x"74",	--3380
		x"75",	--3381
		x"61",	--3382
		x"65",	--3383
		x"0d",	--3384
		x"00",	--3385
		x"25",	--3386
		x"20",	--3387
		x"45",	--3388
		x"49",	--3389
		x"54",	--3390
		x"52",	--3391
		x"56",	--3392
		x"4c",	--3393
		x"45",	--3394
		x"0a",	--3395
		x"53",	--3396
		x"6d",	--3397
		x"74",	--3398
		x"69",	--3399
		x"67",	--3400
		x"77",	--3401
		x"6e",	--3402
		x"20",	--3403
		x"65",	--3404
		x"72",	--3405
		x"62",	--3406
		x"79",	--3407
		x"77",	--3408
		x"6f",	--3409
		x"67",	--3410
		x"0a",	--3411
		x"72",	--3412
		x"25",	--3413
		x"20",	--3414
		x"3d",	--3415
		x"64",	--3416
		x"0a",	--3417
		x"72",	--3418
		x"61",	--3419
		x"0a",	--3420
		x"00",	--3421
		x"25",	--3422
		x"20",	--3423
		x"45",	--3424
		x"49",	--3425
		x"54",	--3426
		x"52",	--3427
		x"0a",	--3428
		x"25",	--3429
		x"20",	--3430
		x"73",	--3431
		x"6e",	--3432
		x"74",	--3433
		x"61",	--3434
		x"6e",	--3435
		x"6d",	--3436
		x"65",	--3437
		x"0d",	--3438
		x"00",	--3439
		x"63",	--3440
		x"25",	--3441
		x"0d",	--3442
		x"00",	--3443
		x"63",	--3444
		x"20",	--3445
		x"6f",	--3446
		x"73",	--3447
		x"63",	--3448
		x"20",	--3449
		x"6f",	--3450
		x"6d",	--3451
		x"6e",	--3452
		x"0d",	--3453
		x"00",	--3454
		x"18",	--3455
		x"46",	--3456
		x"46",	--3457
		x"46",	--3458
		x"46",	--3459
		x"46",	--3460
		x"46",	--3461
		x"46",	--3462
		x"46",	--3463
		x"46",	--3464
		x"46",	--3465
		x"46",	--3466
		x"46",	--3467
		x"46",	--3468
		x"46",	--3469
		x"46",	--3470
		x"46",	--3471
		x"46",	--3472
		x"46",	--3473
		x"46",	--3474
		x"46",	--3475
		x"46",	--3476
		x"46",	--3477
		x"46",	--3478
		x"46",	--3479
		x"46",	--3480
		x"46",	--3481
		x"46",	--3482
		x"46",	--3483
		x"0a",	--3484
		x"46",	--3485
		x"46",	--3486
		x"46",	--3487
		x"46",	--3488
		x"46",	--3489
		x"46",	--3490
		x"46",	--3491
		x"46",	--3492
		x"46",	--3493
		x"46",	--3494
		x"46",	--3495
		x"46",	--3496
		x"46",	--3497
		x"46",	--3498
		x"46",	--3499
		x"46",	--3500
		x"46",	--3501
		x"46",	--3502
		x"46",	--3503
		x"46",	--3504
		x"46",	--3505
		x"46",	--3506
		x"46",	--3507
		x"46",	--3508
		x"46",	--3509
		x"46",	--3510
		x"46",	--3511
		x"46",	--3512
		x"46",	--3513
		x"46",	--3514
		x"46",	--3515
		x"fc",	--3516
		x"ee",	--3517
		x"e0",	--3518
		x"46",	--3519
		x"46",	--3520
		x"46",	--3521
		x"46",	--3522
		x"46",	--3523
		x"46",	--3524
		x"46",	--3525
		x"c8",	--3526
		x"46",	--3527
		x"b6",	--3528
		x"46",	--3529
		x"46",	--3530
		x"46",	--3531
		x"46",	--3532
		x"9a",	--3533
		x"46",	--3534
		x"46",	--3535
		x"46",	--3536
		x"8c",	--3537
		x"7a",	--3538
		x"30",	--3539
		x"32",	--3540
		x"34",	--3541
		x"36",	--3542
		x"38",	--3543
		x"61",	--3544
		x"63",	--3545
		x"65",	--3546
		x"00",	--3547
		x"00",	--3548
		x"00",	--3549
		x"00",	--3550
		x"00",	--3551
		x"00",	--3552
		x"02",	--3553
		x"03",	--3554
		x"03",	--3555
		x"04",	--3556
		x"04",	--3557
		x"04",	--3558
		x"04",	--3559
		x"05",	--3560
		x"05",	--3561
		x"05",	--3562
		x"05",	--3563
		x"05",	--3564
		x"05",	--3565
		x"05",	--3566
		x"05",	--3567
		x"06",	--3568
		x"06",	--3569
		x"06",	--3570
		x"06",	--3571
		x"06",	--3572
		x"06",	--3573
		x"06",	--3574
		x"06",	--3575
		x"06",	--3576
		x"06",	--3577
		x"06",	--3578
		x"06",	--3579
		x"06",	--3580
		x"06",	--3581
		x"06",	--3582
		x"06",	--3583
		x"07",	--3584
		x"07",	--3585
		x"07",	--3586
		x"07",	--3587
		x"07",	--3588
		x"07",	--3589
		x"07",	--3590
		x"07",	--3591
		x"07",	--3592
		x"07",	--3593
		x"07",	--3594
		x"07",	--3595
		x"07",	--3596
		x"07",	--3597
		x"07",	--3598
		x"07",	--3599
		x"07",	--3600
		x"07",	--3601
		x"07",	--3602
		x"07",	--3603
		x"07",	--3604
		x"07",	--3605
		x"07",	--3606
		x"07",	--3607
		x"07",	--3608
		x"07",	--3609
		x"07",	--3610
		x"07",	--3611
		x"07",	--3612
		x"07",	--3613
		x"07",	--3614
		x"07",	--3615
		x"08",	--3616
		x"08",	--3617
		x"08",	--3618
		x"08",	--3619
		x"08",	--3620
		x"08",	--3621
		x"08",	--3622
		x"08",	--3623
		x"08",	--3624
		x"08",	--3625
		x"08",	--3626
		x"08",	--3627
		x"08",	--3628
		x"08",	--3629
		x"08",	--3630
		x"08",	--3631
		x"08",	--3632
		x"08",	--3633
		x"08",	--3634
		x"08",	--3635
		x"08",	--3636
		x"08",	--3637
		x"08",	--3638
		x"08",	--3639
		x"08",	--3640
		x"08",	--3641
		x"08",	--3642
		x"08",	--3643
		x"08",	--3644
		x"08",	--3645
		x"08",	--3646
		x"08",	--3647
		x"08",	--3648
		x"08",	--3649
		x"08",	--3650
		x"08",	--3651
		x"08",	--3652
		x"08",	--3653
		x"08",	--3654
		x"08",	--3655
		x"08",	--3656
		x"08",	--3657
		x"08",	--3658
		x"08",	--3659
		x"08",	--3660
		x"08",	--3661
		x"08",	--3662
		x"08",	--3663
		x"08",	--3664
		x"08",	--3665
		x"08",	--3666
		x"08",	--3667
		x"08",	--3668
		x"08",	--3669
		x"08",	--3670
		x"08",	--3671
		x"08",	--3672
		x"08",	--3673
		x"08",	--3674
		x"08",	--3675
		x"08",	--3676
		x"08",	--3677
		x"08",	--3678
		x"08",	--3679
		x"68",	--3680
		x"6c",	--3681
		x"00",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"b8",	--4080
		x"b8",	--4081
		x"b8",	--4082
		x"b8",	--4083
		x"b8",	--4084
		x"b8",	--4085
		x"b8",	--4086
		x"22",	--4087
		x"da",	--4088
		x"b8",	--4089
		x"b8",	--4090
		x"b8",	--4091
		x"b8",	--4092
		x"b8",	--4093
		x"b8",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"04",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"04",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fc",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"02",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"04",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"25",	--41
		x"43",	--42
		x"12",	--43
		x"eb",	--44
		x"12",	--45
		x"e6",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"fa",	--50
		x"12",	--51
		x"ea",	--52
		x"53",	--53
		x"40",	--54
		x"fa",	--55
		x"40",	--56
		x"e3",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"e6",	--61
		x"40",	--62
		x"fa",	--63
		x"40",	--64
		x"e3",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"e6",	--69
		x"40",	--70
		x"fa",	--71
		x"40",	--72
		x"e1",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"e6",	--77
		x"40",	--78
		x"fa",	--79
		x"40",	--80
		x"e2",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"e6",	--85
		x"40",	--86
		x"fa",	--87
		x"40",	--88
		x"e1",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"e6",	--93
		x"43",	--94
		x"12",	--95
		x"e6",	--96
		x"43",	--97
		x"40",	--98
		x"4e",	--99
		x"40",	--100
		x"01",	--101
		x"41",	--102
		x"50",	--103
		x"00",	--104
		x"12",	--105
		x"e5",	--106
		x"41",	--107
		x"50",	--108
		x"00",	--109
		x"12",	--110
		x"e5",	--111
		x"43",	--112
		x"40",	--113
		x"4e",	--114
		x"40",	--115
		x"01",	--116
		x"41",	--117
		x"52",	--118
		x"12",	--119
		x"e5",	--120
		x"41",	--121
		x"52",	--122
		x"12",	--123
		x"e5",	--124
		x"41",	--125
		x"52",	--126
		x"41",	--127
		x"50",	--128
		x"00",	--129
		x"12",	--130
		x"e1",	--131
		x"40",	--132
		x"01",	--133
		x"41",	--134
		x"53",	--135
		x"12",	--136
		x"e8",	--137
		x"40",	--138
		x"01",	--139
		x"41",	--140
		x"12",	--141
		x"e8",	--142
		x"41",	--143
		x"41",	--144
		x"53",	--145
		x"12",	--146
		x"e2",	--147
		x"12",	--148
		x"e7",	--149
		x"43",	--150
		x"40",	--151
		x"e2",	--152
		x"43",	--153
		x"12",	--154
		x"e7",	--155
		x"12",	--156
		x"e7",	--157
		x"40",	--158
		x"ff",	--159
		x"00",	--160
		x"d2",	--161
		x"43",	--162
		x"12",	--163
		x"eb",	--164
		x"93",	--165
		x"27",	--166
		x"12",	--167
		x"eb",	--168
		x"92",	--169
		x"24",	--170
		x"90",	--171
		x"00",	--172
		x"20",	--173
		x"12",	--174
		x"fa",	--175
		x"12",	--176
		x"ea",	--177
		x"53",	--178
		x"41",	--179
		x"50",	--180
		x"00",	--181
		x"41",	--182
		x"00",	--183
		x"12",	--184
		x"e7",	--185
		x"43",	--186
		x"3f",	--187
		x"93",	--188
		x"27",	--189
		x"53",	--190
		x"12",	--191
		x"fa",	--192
		x"12",	--193
		x"ea",	--194
		x"53",	--195
		x"3f",	--196
		x"90",	--197
		x"00",	--198
		x"2f",	--199
		x"4f",	--200
		x"11",	--201
		x"12",	--202
		x"12",	--203
		x"fa",	--204
		x"4f",	--205
		x"00",	--206
		x"12",	--207
		x"ea",	--208
		x"52",	--209
		x"40",	--210
		x"00",	--211
		x"51",	--212
		x"5b",	--213
		x"41",	--214
		x"00",	--215
		x"4f",	--216
		x"00",	--217
		x"53",	--218
		x"3f",	--219
		x"40",	--220
		x"f9",	--221
		x"40",	--222
		x"e0",	--223
		x"01",	--224
		x"42",	--225
		x"01",	--226
		x"40",	--227
		x"02",	--228
		x"01",	--229
		x"12",	--230
		x"f9",	--231
		x"12",	--232
		x"ea",	--233
		x"43",	--234
		x"01",	--235
		x"40",	--236
		x"f9",	--237
		x"00",	--238
		x"12",	--239
		x"ea",	--240
		x"53",	--241
		x"43",	--242
		x"41",	--243
		x"4f",	--244
		x"02",	--245
		x"4e",	--246
		x"02",	--247
		x"41",	--248
		x"82",	--249
		x"90",	--250
		x"00",	--251
		x"00",	--252
		x"20",	--253
		x"93",	--254
		x"00",	--255
		x"24",	--256
		x"41",	--257
		x"4f",	--258
		x"53",	--259
		x"41",	--260
		x"52",	--261
		x"12",	--262
		x"e4",	--263
		x"93",	--264
		x"00",	--265
		x"24",	--266
		x"41",	--267
		x"4f",	--268
		x"41",	--269
		x"53",	--270
		x"12",	--271
		x"e4",	--272
		x"93",	--273
		x"00",	--274
		x"24",	--275
		x"41",	--276
		x"00",	--277
		x"43",	--278
		x"12",	--279
		x"f3",	--280
		x"43",	--281
		x"40",	--282
		x"42",	--283
		x"12",	--284
		x"f1",	--285
		x"4e",	--286
		x"4f",	--287
		x"42",	--288
		x"02",	--289
		x"12",	--290
		x"e6",	--291
		x"41",	--292
		x"00",	--293
		x"43",	--294
		x"12",	--295
		x"f3",	--296
		x"43",	--297
		x"40",	--298
		x"42",	--299
		x"12",	--300
		x"f1",	--301
		x"4e",	--302
		x"4f",	--303
		x"42",	--304
		x"02",	--305
		x"12",	--306
		x"e6",	--307
		x"43",	--308
		x"52",	--309
		x"41",	--310
		x"12",	--311
		x"f9",	--312
		x"4f",	--313
		x"00",	--314
		x"12",	--315
		x"ea",	--316
		x"41",	--317
		x"00",	--318
		x"4f",	--319
		x"11",	--320
		x"4f",	--321
		x"00",	--322
		x"12",	--323
		x"f9",	--324
		x"12",	--325
		x"ea",	--326
		x"52",	--327
		x"43",	--328
		x"52",	--329
		x"41",	--330
		x"12",	--331
		x"f9",	--332
		x"12",	--333
		x"ea",	--334
		x"53",	--335
		x"43",	--336
		x"3f",	--337
		x"4f",	--338
		x"02",	--339
		x"4e",	--340
		x"02",	--341
		x"41",	--342
		x"42",	--343
		x"02",	--344
		x"4f",	--345
		x"42",	--346
		x"02",	--347
		x"4f",	--348
		x"12",	--349
		x"12",	--350
		x"00",	--351
		x"12",	--352
		x"12",	--353
		x"00",	--354
		x"12",	--355
		x"f9",	--356
		x"12",	--357
		x"ea",	--358
		x"50",	--359
		x"00",	--360
		x"43",	--361
		x"41",	--362
		x"42",	--363
		x"02",	--364
		x"92",	--365
		x"2c",	--366
		x"4e",	--367
		x"5f",	--368
		x"4f",	--369
		x"fa",	--370
		x"43",	--371
		x"00",	--372
		x"90",	--373
		x"00",	--374
		x"38",	--375
		x"43",	--376
		x"02",	--377
		x"41",	--378
		x"53",	--379
		x"4e",	--380
		x"02",	--381
		x"41",	--382
		x"40",	--383
		x"00",	--384
		x"00",	--385
		x"3f",	--386
		x"40",	--387
		x"00",	--388
		x"00",	--389
		x"3f",	--390
		x"42",	--391
		x"00",	--392
		x"3f",	--393
		x"40",	--394
		x"00",	--395
		x"00",	--396
		x"3f",	--397
		x"40",	--398
		x"00",	--399
		x"00",	--400
		x"3f",	--401
		x"40",	--402
		x"00",	--403
		x"00",	--404
		x"3f",	--405
		x"40",	--406
		x"00",	--407
		x"00",	--408
		x"3f",	--409
		x"42",	--410
		x"00",	--411
		x"4e",	--412
		x"be",	--413
		x"20",	--414
		x"df",	--415
		x"00",	--416
		x"41",	--417
		x"cf",	--418
		x"00",	--419
		x"41",	--420
		x"12",	--421
		x"50",	--422
		x"ff",	--423
		x"4f",	--424
		x"12",	--425
		x"fa",	--426
		x"12",	--427
		x"ea",	--428
		x"53",	--429
		x"90",	--430
		x"00",	--431
		x"00",	--432
		x"20",	--433
		x"93",	--434
		x"00",	--435
		x"24",	--436
		x"41",	--437
		x"4b",	--438
		x"53",	--439
		x"41",	--440
		x"52",	--441
		x"12",	--442
		x"e4",	--443
		x"93",	--444
		x"00",	--445
		x"24",	--446
		x"41",	--447
		x"4f",	--448
		x"41",	--449
		x"53",	--450
		x"12",	--451
		x"e4",	--452
		x"93",	--453
		x"00",	--454
		x"24",	--455
		x"12",	--456
		x"00",	--457
		x"12",	--458
		x"00",	--459
		x"12",	--460
		x"fa",	--461
		x"12",	--462
		x"ea",	--463
		x"50",	--464
		x"00",	--465
		x"41",	--466
		x"00",	--467
		x"41",	--468
		x"00",	--469
		x"00",	--470
		x"43",	--471
		x"50",	--472
		x"00",	--473
		x"41",	--474
		x"41",	--475
		x"12",	--476
		x"fa",	--477
		x"12",	--478
		x"ea",	--479
		x"4b",	--480
		x"11",	--481
		x"4f",	--482
		x"00",	--483
		x"12",	--484
		x"fa",	--485
		x"12",	--486
		x"ea",	--487
		x"52",	--488
		x"43",	--489
		x"50",	--490
		x"00",	--491
		x"41",	--492
		x"41",	--493
		x"12",	--494
		x"fa",	--495
		x"12",	--496
		x"ea",	--497
		x"53",	--498
		x"43",	--499
		x"3f",	--500
		x"12",	--501
		x"82",	--502
		x"4f",	--503
		x"12",	--504
		x"fa",	--505
		x"12",	--506
		x"ea",	--507
		x"53",	--508
		x"90",	--509
		x"00",	--510
		x"00",	--511
		x"20",	--512
		x"93",	--513
		x"00",	--514
		x"24",	--515
		x"41",	--516
		x"4b",	--517
		x"53",	--518
		x"41",	--519
		x"53",	--520
		x"12",	--521
		x"e4",	--522
		x"93",	--523
		x"00",	--524
		x"24",	--525
		x"41",	--526
		x"00",	--527
		x"12",	--528
		x"12",	--529
		x"12",	--530
		x"fa",	--531
		x"12",	--532
		x"ea",	--533
		x"50",	--534
		x"00",	--535
		x"43",	--536
		x"52",	--537
		x"41",	--538
		x"41",	--539
		x"12",	--540
		x"fa",	--541
		x"12",	--542
		x"ea",	--543
		x"4b",	--544
		x"11",	--545
		x"4f",	--546
		x"00",	--547
		x"12",	--548
		x"fa",	--549
		x"12",	--550
		x"ea",	--551
		x"52",	--552
		x"43",	--553
		x"52",	--554
		x"41",	--555
		x"41",	--556
		x"12",	--557
		x"fa",	--558
		x"12",	--559
		x"ea",	--560
		x"53",	--561
		x"43",	--562
		x"3f",	--563
		x"12",	--564
		x"12",	--565
		x"12",	--566
		x"12",	--567
		x"12",	--568
		x"43",	--569
		x"00",	--570
		x"43",	--571
		x"00",	--572
		x"4e",	--573
		x"93",	--574
		x"24",	--575
		x"4e",	--576
		x"53",	--577
		x"4e",	--578
		x"43",	--579
		x"43",	--580
		x"43",	--581
		x"3c",	--582
		x"90",	--583
		x"00",	--584
		x"2c",	--585
		x"4f",	--586
		x"5c",	--587
		x"5c",	--588
		x"5c",	--589
		x"5c",	--590
		x"4c",	--591
		x"00",	--592
		x"50",	--593
		x"ff",	--594
		x"48",	--595
		x"11",	--596
		x"5a",	--597
		x"4c",	--598
		x"00",	--599
		x"43",	--600
		x"53",	--601
		x"49",	--602
		x"4b",	--603
		x"4b",	--604
		x"93",	--605
		x"24",	--606
		x"90",	--607
		x"00",	--608
		x"24",	--609
		x"90",	--610
		x"00",	--611
		x"24",	--612
		x"4c",	--613
		x"50",	--614
		x"ff",	--615
		x"93",	--616
		x"23",	--617
		x"90",	--618
		x"00",	--619
		x"2c",	--620
		x"4f",	--621
		x"5a",	--622
		x"4a",	--623
		x"5c",	--624
		x"5c",	--625
		x"5a",	--626
		x"4c",	--627
		x"00",	--628
		x"50",	--629
		x"ff",	--630
		x"48",	--631
		x"11",	--632
		x"58",	--633
		x"4c",	--634
		x"00",	--635
		x"3f",	--636
		x"43",	--637
		x"3f",	--638
		x"4c",	--639
		x"50",	--640
		x"ff",	--641
		x"90",	--642
		x"00",	--643
		x"2c",	--644
		x"4f",	--645
		x"5c",	--646
		x"5c",	--647
		x"5c",	--648
		x"5c",	--649
		x"4c",	--650
		x"00",	--651
		x"50",	--652
		x"ff",	--653
		x"3f",	--654
		x"4c",	--655
		x"50",	--656
		x"ff",	--657
		x"90",	--658
		x"00",	--659
		x"2c",	--660
		x"4f",	--661
		x"5c",	--662
		x"5c",	--663
		x"5c",	--664
		x"5c",	--665
		x"4c",	--666
		x"00",	--667
		x"50",	--668
		x"ff",	--669
		x"3f",	--670
		x"43",	--671
		x"00",	--672
		x"43",	--673
		x"41",	--674
		x"41",	--675
		x"41",	--676
		x"41",	--677
		x"41",	--678
		x"41",	--679
		x"43",	--680
		x"00",	--681
		x"4a",	--682
		x"53",	--683
		x"5e",	--684
		x"41",	--685
		x"41",	--686
		x"41",	--687
		x"41",	--688
		x"41",	--689
		x"41",	--690
		x"11",	--691
		x"12",	--692
		x"12",	--693
		x"fa",	--694
		x"12",	--695
		x"ea",	--696
		x"52",	--697
		x"43",	--698
		x"41",	--699
		x"41",	--700
		x"41",	--701
		x"41",	--702
		x"41",	--703
		x"41",	--704
		x"12",	--705
		x"12",	--706
		x"4e",	--707
		x"4c",	--708
		x"4e",	--709
		x"00",	--710
		x"4d",	--711
		x"00",	--712
		x"4c",	--713
		x"00",	--714
		x"4d",	--715
		x"43",	--716
		x"40",	--717
		x"36",	--718
		x"40",	--719
		x"01",	--720
		x"12",	--721
		x"f8",	--722
		x"4e",	--723
		x"00",	--724
		x"12",	--725
		x"c2",	--726
		x"43",	--727
		x"4a",	--728
		x"01",	--729
		x"40",	--730
		x"00",	--731
		x"01",	--732
		x"42",	--733
		x"01",	--734
		x"00",	--735
		x"41",	--736
		x"43",	--737
		x"41",	--738
		x"41",	--739
		x"41",	--740
		x"12",	--741
		x"12",	--742
		x"12",	--743
		x"43",	--744
		x"00",	--745
		x"40",	--746
		x"3f",	--747
		x"00",	--748
		x"4f",	--749
		x"4b",	--750
		x"00",	--751
		x"43",	--752
		x"12",	--753
		x"f3",	--754
		x"43",	--755
		x"40",	--756
		x"3f",	--757
		x"12",	--758
		x"ef",	--759
		x"4e",	--760
		x"4f",	--761
		x"4b",	--762
		x"00",	--763
		x"43",	--764
		x"12",	--765
		x"f3",	--766
		x"4e",	--767
		x"4f",	--768
		x"48",	--769
		x"49",	--770
		x"12",	--771
		x"ee",	--772
		x"12",	--773
		x"eb",	--774
		x"4e",	--775
		x"00",	--776
		x"43",	--777
		x"00",	--778
		x"41",	--779
		x"41",	--780
		x"41",	--781
		x"41",	--782
		x"12",	--783
		x"12",	--784
		x"12",	--785
		x"4d",	--786
		x"4e",	--787
		x"4d",	--788
		x"00",	--789
		x"4e",	--790
		x"00",	--791
		x"4f",	--792
		x"49",	--793
		x"00",	--794
		x"43",	--795
		x"12",	--796
		x"f3",	--797
		x"4e",	--798
		x"4f",	--799
		x"4a",	--800
		x"4b",	--801
		x"12",	--802
		x"ef",	--803
		x"4e",	--804
		x"4f",	--805
		x"49",	--806
		x"00",	--807
		x"43",	--808
		x"12",	--809
		x"f3",	--810
		x"4e",	--811
		x"4f",	--812
		x"4a",	--813
		x"4b",	--814
		x"12",	--815
		x"ee",	--816
		x"12",	--817
		x"eb",	--818
		x"4e",	--819
		x"00",	--820
		x"41",	--821
		x"41",	--822
		x"41",	--823
		x"41",	--824
		x"12",	--825
		x"12",	--826
		x"93",	--827
		x"02",	--828
		x"38",	--829
		x"40",	--830
		x"02",	--831
		x"43",	--832
		x"12",	--833
		x"4b",	--834
		x"ff",	--835
		x"11",	--836
		x"12",	--837
		x"12",	--838
		x"fa",	--839
		x"12",	--840
		x"ea",	--841
		x"50",	--842
		x"00",	--843
		x"53",	--844
		x"50",	--845
		x"00",	--846
		x"92",	--847
		x"02",	--848
		x"3b",	--849
		x"43",	--850
		x"41",	--851
		x"41",	--852
		x"41",	--853
		x"42",	--854
		x"02",	--855
		x"90",	--856
		x"00",	--857
		x"34",	--858
		x"4e",	--859
		x"5f",	--860
		x"5e",	--861
		x"5f",	--862
		x"50",	--863
		x"02",	--864
		x"40",	--865
		x"00",	--866
		x"00",	--867
		x"40",	--868
		x"e6",	--869
		x"00",	--870
		x"40",	--871
		x"02",	--872
		x"00",	--873
		x"53",	--874
		x"4e",	--875
		x"02",	--876
		x"41",	--877
		x"12",	--878
		x"42",	--879
		x"02",	--880
		x"90",	--881
		x"00",	--882
		x"34",	--883
		x"4b",	--884
		x"5c",	--885
		x"5b",	--886
		x"5c",	--887
		x"50",	--888
		x"02",	--889
		x"4f",	--890
		x"00",	--891
		x"4e",	--892
		x"00",	--893
		x"4d",	--894
		x"00",	--895
		x"53",	--896
		x"4b",	--897
		x"02",	--898
		x"43",	--899
		x"41",	--900
		x"41",	--901
		x"43",	--902
		x"3f",	--903
		x"12",	--904
		x"42",	--905
		x"02",	--906
		x"93",	--907
		x"38",	--908
		x"92",	--909
		x"02",	--910
		x"24",	--911
		x"40",	--912
		x"02",	--913
		x"43",	--914
		x"3c",	--915
		x"50",	--916
		x"00",	--917
		x"9f",	--918
		x"ff",	--919
		x"24",	--920
		x"53",	--921
		x"9b",	--922
		x"23",	--923
		x"12",	--924
		x"fa",	--925
		x"12",	--926
		x"ea",	--927
		x"53",	--928
		x"43",	--929
		x"41",	--930
		x"41",	--931
		x"43",	--932
		x"4c",	--933
		x"5d",	--934
		x"5d",	--935
		x"5c",	--936
		x"50",	--937
		x"02",	--938
		x"4e",	--939
		x"12",	--940
		x"00",	--941
		x"41",	--942
		x"41",	--943
		x"d0",	--944
		x"02",	--945
		x"01",	--946
		x"40",	--947
		x"0b",	--948
		x"01",	--949
		x"43",	--950
		x"41",	--951
		x"12",	--952
		x"12",	--953
		x"4f",	--954
		x"42",	--955
		x"02",	--956
		x"90",	--957
		x"00",	--958
		x"34",	--959
		x"4f",	--960
		x"5b",	--961
		x"4b",	--962
		x"5c",	--963
		x"5c",	--964
		x"5b",	--965
		x"50",	--966
		x"02",	--967
		x"43",	--968
		x"00",	--969
		x"43",	--970
		x"00",	--971
		x"4a",	--972
		x"00",	--973
		x"4e",	--974
		x"00",	--975
		x"4d",	--976
		x"00",	--977
		x"4f",	--978
		x"53",	--979
		x"4e",	--980
		x"02",	--981
		x"41",	--982
		x"41",	--983
		x"41",	--984
		x"43",	--985
		x"3f",	--986
		x"5f",	--987
		x"4f",	--988
		x"5e",	--989
		x"5e",	--990
		x"5f",	--991
		x"43",	--992
		x"02",	--993
		x"43",	--994
		x"41",	--995
		x"5f",	--996
		x"4f",	--997
		x"5e",	--998
		x"5e",	--999
		x"5f",	--1000
		x"43",	--1001
		x"02",	--1002
		x"43",	--1003
		x"41",	--1004
		x"12",	--1005
		x"12",	--1006
		x"12",	--1007
		x"12",	--1008
		x"12",	--1009
		x"12",	--1010
		x"93",	--1011
		x"02",	--1012
		x"38",	--1013
		x"40",	--1014
		x"02",	--1015
		x"43",	--1016
		x"3c",	--1017
		x"53",	--1018
		x"4f",	--1019
		x"00",	--1020
		x"53",	--1021
		x"50",	--1022
		x"00",	--1023
		x"92",	--1024
		x"02",	--1025
		x"34",	--1026
		x"93",	--1027
		x"ff",	--1028
		x"27",	--1029
		x"4b",	--1030
		x"9b",	--1031
		x"00",	--1032
		x"2b",	--1033
		x"43",	--1034
		x"00",	--1035
		x"4b",	--1036
		x"00",	--1037
		x"12",	--1038
		x"00",	--1039
		x"53",	--1040
		x"50",	--1041
		x"00",	--1042
		x"92",	--1043
		x"02",	--1044
		x"3b",	--1045
		x"f0",	--1046
		x"ff",	--1047
		x"01",	--1048
		x"41",	--1049
		x"41",	--1050
		x"41",	--1051
		x"41",	--1052
		x"41",	--1053
		x"41",	--1054
		x"13",	--1055
		x"4e",	--1056
		x"00",	--1057
		x"43",	--1058
		x"41",	--1059
		x"4f",	--1060
		x"4f",	--1061
		x"41",	--1062
		x"42",	--1063
		x"00",	--1064
		x"f2",	--1065
		x"23",	--1066
		x"4f",	--1067
		x"00",	--1068
		x"43",	--1069
		x"41",	--1070
		x"f0",	--1071
		x"00",	--1072
		x"4f",	--1073
		x"fb",	--1074
		x"11",	--1075
		x"12",	--1076
		x"e8",	--1077
		x"41",	--1078
		x"12",	--1079
		x"4f",	--1080
		x"4f",	--1081
		x"11",	--1082
		x"11",	--1083
		x"11",	--1084
		x"11",	--1085
		x"4e",	--1086
		x"12",	--1087
		x"e8",	--1088
		x"4b",	--1089
		x"12",	--1090
		x"e8",	--1091
		x"41",	--1092
		x"41",	--1093
		x"12",	--1094
		x"12",	--1095
		x"4f",	--1096
		x"40",	--1097
		x"00",	--1098
		x"4a",	--1099
		x"4b",	--1100
		x"f0",	--1101
		x"00",	--1102
		x"24",	--1103
		x"11",	--1104
		x"53",	--1105
		x"23",	--1106
		x"f3",	--1107
		x"24",	--1108
		x"40",	--1109
		x"00",	--1110
		x"12",	--1111
		x"e8",	--1112
		x"53",	--1113
		x"93",	--1114
		x"23",	--1115
		x"41",	--1116
		x"41",	--1117
		x"41",	--1118
		x"40",	--1119
		x"00",	--1120
		x"3f",	--1121
		x"12",	--1122
		x"4f",	--1123
		x"4f",	--1124
		x"10",	--1125
		x"11",	--1126
		x"4e",	--1127
		x"12",	--1128
		x"e8",	--1129
		x"4b",	--1130
		x"12",	--1131
		x"e8",	--1132
		x"41",	--1133
		x"41",	--1134
		x"12",	--1135
		x"12",	--1136
		x"4e",	--1137
		x"4f",	--1138
		x"4f",	--1139
		x"10",	--1140
		x"11",	--1141
		x"4d",	--1142
		x"12",	--1143
		x"e8",	--1144
		x"4b",	--1145
		x"12",	--1146
		x"e8",	--1147
		x"4b",	--1148
		x"4a",	--1149
		x"10",	--1150
		x"10",	--1151
		x"ec",	--1152
		x"ec",	--1153
		x"4d",	--1154
		x"12",	--1155
		x"e8",	--1156
		x"4a",	--1157
		x"12",	--1158
		x"e8",	--1159
		x"41",	--1160
		x"41",	--1161
		x"41",	--1162
		x"12",	--1163
		x"12",	--1164
		x"12",	--1165
		x"4f",	--1166
		x"93",	--1167
		x"24",	--1168
		x"4e",	--1169
		x"53",	--1170
		x"43",	--1171
		x"4a",	--1172
		x"5b",	--1173
		x"4d",	--1174
		x"11",	--1175
		x"12",	--1176
		x"e8",	--1177
		x"99",	--1178
		x"24",	--1179
		x"53",	--1180
		x"b0",	--1181
		x"00",	--1182
		x"20",	--1183
		x"40",	--1184
		x"00",	--1185
		x"12",	--1186
		x"e8",	--1187
		x"3f",	--1188
		x"40",	--1189
		x"00",	--1190
		x"12",	--1191
		x"e8",	--1192
		x"3f",	--1193
		x"41",	--1194
		x"41",	--1195
		x"41",	--1196
		x"41",	--1197
		x"12",	--1198
		x"12",	--1199
		x"12",	--1200
		x"4f",	--1201
		x"93",	--1202
		x"24",	--1203
		x"4e",	--1204
		x"53",	--1205
		x"43",	--1206
		x"4a",	--1207
		x"11",	--1208
		x"12",	--1209
		x"e8",	--1210
		x"99",	--1211
		x"24",	--1212
		x"53",	--1213
		x"b0",	--1214
		x"00",	--1215
		x"23",	--1216
		x"40",	--1217
		x"00",	--1218
		x"12",	--1219
		x"e8",	--1220
		x"4a",	--1221
		x"11",	--1222
		x"12",	--1223
		x"e8",	--1224
		x"99",	--1225
		x"23",	--1226
		x"41",	--1227
		x"41",	--1228
		x"41",	--1229
		x"41",	--1230
		x"12",	--1231
		x"12",	--1232
		x"12",	--1233
		x"50",	--1234
		x"ff",	--1235
		x"4f",	--1236
		x"93",	--1237
		x"38",	--1238
		x"90",	--1239
		x"00",	--1240
		x"38",	--1241
		x"43",	--1242
		x"41",	--1243
		x"59",	--1244
		x"40",	--1245
		x"00",	--1246
		x"4b",	--1247
		x"12",	--1248
		x"f8",	--1249
		x"50",	--1250
		x"00",	--1251
		x"4f",	--1252
		x"00",	--1253
		x"53",	--1254
		x"40",	--1255
		x"00",	--1256
		x"4b",	--1257
		x"12",	--1258
		x"f8",	--1259
		x"4f",	--1260
		x"90",	--1261
		x"00",	--1262
		x"37",	--1263
		x"49",	--1264
		x"53",	--1265
		x"51",	--1266
		x"40",	--1267
		x"00",	--1268
		x"4b",	--1269
		x"12",	--1270
		x"f8",	--1271
		x"50",	--1272
		x"00",	--1273
		x"4f",	--1274
		x"00",	--1275
		x"53",	--1276
		x"41",	--1277
		x"5a",	--1278
		x"4f",	--1279
		x"11",	--1280
		x"12",	--1281
		x"e8",	--1282
		x"93",	--1283
		x"23",	--1284
		x"50",	--1285
		x"00",	--1286
		x"41",	--1287
		x"41",	--1288
		x"41",	--1289
		x"41",	--1290
		x"40",	--1291
		x"00",	--1292
		x"12",	--1293
		x"e8",	--1294
		x"e3",	--1295
		x"53",	--1296
		x"3f",	--1297
		x"43",	--1298
		x"43",	--1299
		x"3f",	--1300
		x"12",	--1301
		x"12",	--1302
		x"12",	--1303
		x"41",	--1304
		x"52",	--1305
		x"4b",	--1306
		x"49",	--1307
		x"93",	--1308
		x"20",	--1309
		x"3c",	--1310
		x"11",	--1311
		x"12",	--1312
		x"e8",	--1313
		x"49",	--1314
		x"4a",	--1315
		x"53",	--1316
		x"4a",	--1317
		x"00",	--1318
		x"93",	--1319
		x"24",	--1320
		x"90",	--1321
		x"00",	--1322
		x"23",	--1323
		x"49",	--1324
		x"53",	--1325
		x"49",	--1326
		x"00",	--1327
		x"50",	--1328
		x"ff",	--1329
		x"90",	--1330
		x"00",	--1331
		x"2f",	--1332
		x"4f",	--1333
		x"5f",	--1334
		x"4f",	--1335
		x"fa",	--1336
		x"41",	--1337
		x"41",	--1338
		x"41",	--1339
		x"41",	--1340
		x"4b",	--1341
		x"52",	--1342
		x"4b",	--1343
		x"00",	--1344
		x"4b",	--1345
		x"12",	--1346
		x"e9",	--1347
		x"49",	--1348
		x"3f",	--1349
		x"4b",	--1350
		x"53",	--1351
		x"4b",	--1352
		x"12",	--1353
		x"e8",	--1354
		x"49",	--1355
		x"3f",	--1356
		x"4b",	--1357
		x"53",	--1358
		x"4f",	--1359
		x"49",	--1360
		x"93",	--1361
		x"27",	--1362
		x"53",	--1363
		x"11",	--1364
		x"12",	--1365
		x"e8",	--1366
		x"49",	--1367
		x"93",	--1368
		x"23",	--1369
		x"3f",	--1370
		x"4b",	--1371
		x"52",	--1372
		x"4b",	--1373
		x"00",	--1374
		x"4b",	--1375
		x"12",	--1376
		x"e9",	--1377
		x"49",	--1378
		x"3f",	--1379
		x"4b",	--1380
		x"53",	--1381
		x"4b",	--1382
		x"4e",	--1383
		x"10",	--1384
		x"11",	--1385
		x"10",	--1386
		x"11",	--1387
		x"12",	--1388
		x"e8",	--1389
		x"49",	--1390
		x"3f",	--1391
		x"4b",	--1392
		x"53",	--1393
		x"4b",	--1394
		x"12",	--1395
		x"e9",	--1396
		x"49",	--1397
		x"3f",	--1398
		x"4b",	--1399
		x"53",	--1400
		x"4b",	--1401
		x"12",	--1402
		x"e8",	--1403
		x"49",	--1404
		x"3f",	--1405
		x"4b",	--1406
		x"53",	--1407
		x"4b",	--1408
		x"12",	--1409
		x"e8",	--1410
		x"49",	--1411
		x"3f",	--1412
		x"4b",	--1413
		x"53",	--1414
		x"4b",	--1415
		x"12",	--1416
		x"e8",	--1417
		x"49",	--1418
		x"3f",	--1419
		x"40",	--1420
		x"00",	--1421
		x"12",	--1422
		x"e8",	--1423
		x"3f",	--1424
		x"12",	--1425
		x"12",	--1426
		x"42",	--1427
		x"02",	--1428
		x"42",	--1429
		x"00",	--1430
		x"04",	--1431
		x"42",	--1432
		x"02",	--1433
		x"90",	--1434
		x"00",	--1435
		x"34",	--1436
		x"53",	--1437
		x"02",	--1438
		x"42",	--1439
		x"02",	--1440
		x"42",	--1441
		x"02",	--1442
		x"9f",	--1443
		x"20",	--1444
		x"53",	--1445
		x"02",	--1446
		x"40",	--1447
		x"00",	--1448
		x"00",	--1449
		x"41",	--1450
		x"41",	--1451
		x"c0",	--1452
		x"00",	--1453
		x"00",	--1454
		x"13",	--1455
		x"43",	--1456
		x"02",	--1457
		x"3f",	--1458
		x"40",	--1459
		x"09",	--1460
		x"00",	--1461
		x"40",	--1462
		x"00",	--1463
		x"00",	--1464
		x"41",	--1465
		x"42",	--1466
		x"02",	--1467
		x"42",	--1468
		x"02",	--1469
		x"9f",	--1470
		x"38",	--1471
		x"42",	--1472
		x"02",	--1473
		x"82",	--1474
		x"02",	--1475
		x"41",	--1476
		x"42",	--1477
		x"02",	--1478
		x"42",	--1479
		x"02",	--1480
		x"40",	--1481
		x"00",	--1482
		x"8d",	--1483
		x"8e",	--1484
		x"41",	--1485
		x"42",	--1486
		x"02",	--1487
		x"4f",	--1488
		x"04",	--1489
		x"42",	--1490
		x"02",	--1491
		x"42",	--1492
		x"02",	--1493
		x"9e",	--1494
		x"24",	--1495
		x"42",	--1496
		x"02",	--1497
		x"90",	--1498
		x"00",	--1499
		x"38",	--1500
		x"43",	--1501
		x"02",	--1502
		x"41",	--1503
		x"53",	--1504
		x"02",	--1505
		x"41",	--1506
		x"43",	--1507
		x"41",	--1508
		x"12",	--1509
		x"12",	--1510
		x"4e",	--1511
		x"4f",	--1512
		x"43",	--1513
		x"40",	--1514
		x"4f",	--1515
		x"12",	--1516
		x"f2",	--1517
		x"93",	--1518
		x"34",	--1519
		x"4a",	--1520
		x"4b",	--1521
		x"12",	--1522
		x"f2",	--1523
		x"41",	--1524
		x"41",	--1525
		x"41",	--1526
		x"43",	--1527
		x"40",	--1528
		x"4f",	--1529
		x"4a",	--1530
		x"4b",	--1531
		x"12",	--1532
		x"ee",	--1533
		x"12",	--1534
		x"f2",	--1535
		x"53",	--1536
		x"60",	--1537
		x"80",	--1538
		x"41",	--1539
		x"41",	--1540
		x"41",	--1541
		x"12",	--1542
		x"12",	--1543
		x"12",	--1544
		x"12",	--1545
		x"12",	--1546
		x"12",	--1547
		x"12",	--1548
		x"12",	--1549
		x"50",	--1550
		x"ff",	--1551
		x"4d",	--1552
		x"4f",	--1553
		x"93",	--1554
		x"28",	--1555
		x"4e",	--1556
		x"93",	--1557
		x"28",	--1558
		x"92",	--1559
		x"20",	--1560
		x"40",	--1561
		x"ee",	--1562
		x"92",	--1563
		x"24",	--1564
		x"93",	--1565
		x"24",	--1566
		x"93",	--1567
		x"24",	--1568
		x"4f",	--1569
		x"00",	--1570
		x"00",	--1571
		x"4e",	--1572
		x"00",	--1573
		x"4f",	--1574
		x"00",	--1575
		x"4f",	--1576
		x"00",	--1577
		x"4e",	--1578
		x"00",	--1579
		x"4e",	--1580
		x"00",	--1581
		x"41",	--1582
		x"8b",	--1583
		x"4c",	--1584
		x"93",	--1585
		x"38",	--1586
		x"90",	--1587
		x"00",	--1588
		x"34",	--1589
		x"93",	--1590
		x"38",	--1591
		x"46",	--1592
		x"00",	--1593
		x"47",	--1594
		x"00",	--1595
		x"49",	--1596
		x"f0",	--1597
		x"00",	--1598
		x"24",	--1599
		x"46",	--1600
		x"47",	--1601
		x"c3",	--1602
		x"10",	--1603
		x"10",	--1604
		x"53",	--1605
		x"23",	--1606
		x"4a",	--1607
		x"00",	--1608
		x"4b",	--1609
		x"00",	--1610
		x"43",	--1611
		x"43",	--1612
		x"f0",	--1613
		x"00",	--1614
		x"24",	--1615
		x"5c",	--1616
		x"6d",	--1617
		x"53",	--1618
		x"23",	--1619
		x"53",	--1620
		x"63",	--1621
		x"f6",	--1622
		x"f7",	--1623
		x"43",	--1624
		x"43",	--1625
		x"93",	--1626
		x"20",	--1627
		x"93",	--1628
		x"24",	--1629
		x"41",	--1630
		x"00",	--1631
		x"41",	--1632
		x"00",	--1633
		x"da",	--1634
		x"db",	--1635
		x"4f",	--1636
		x"00",	--1637
		x"9e",	--1638
		x"00",	--1639
		x"20",	--1640
		x"4f",	--1641
		x"00",	--1642
		x"41",	--1643
		x"00",	--1644
		x"46",	--1645
		x"47",	--1646
		x"54",	--1647
		x"65",	--1648
		x"4e",	--1649
		x"00",	--1650
		x"4f",	--1651
		x"00",	--1652
		x"40",	--1653
		x"00",	--1654
		x"00",	--1655
		x"93",	--1656
		x"38",	--1657
		x"48",	--1658
		x"50",	--1659
		x"00",	--1660
		x"41",	--1661
		x"41",	--1662
		x"41",	--1663
		x"41",	--1664
		x"41",	--1665
		x"41",	--1666
		x"41",	--1667
		x"41",	--1668
		x"41",	--1669
		x"91",	--1670
		x"38",	--1671
		x"4b",	--1672
		x"00",	--1673
		x"43",	--1674
		x"43",	--1675
		x"4f",	--1676
		x"00",	--1677
		x"9e",	--1678
		x"00",	--1679
		x"27",	--1680
		x"93",	--1681
		x"24",	--1682
		x"46",	--1683
		x"47",	--1684
		x"84",	--1685
		x"75",	--1686
		x"93",	--1687
		x"38",	--1688
		x"43",	--1689
		x"00",	--1690
		x"41",	--1691
		x"00",	--1692
		x"4e",	--1693
		x"00",	--1694
		x"4f",	--1695
		x"00",	--1696
		x"4e",	--1697
		x"4f",	--1698
		x"53",	--1699
		x"63",	--1700
		x"90",	--1701
		x"3f",	--1702
		x"28",	--1703
		x"90",	--1704
		x"40",	--1705
		x"2c",	--1706
		x"93",	--1707
		x"2c",	--1708
		x"48",	--1709
		x"00",	--1710
		x"53",	--1711
		x"5e",	--1712
		x"6f",	--1713
		x"4b",	--1714
		x"53",	--1715
		x"4e",	--1716
		x"4f",	--1717
		x"53",	--1718
		x"63",	--1719
		x"90",	--1720
		x"3f",	--1721
		x"2b",	--1722
		x"24",	--1723
		x"4e",	--1724
		x"00",	--1725
		x"4f",	--1726
		x"00",	--1727
		x"4a",	--1728
		x"00",	--1729
		x"40",	--1730
		x"00",	--1731
		x"00",	--1732
		x"93",	--1733
		x"37",	--1734
		x"4e",	--1735
		x"4f",	--1736
		x"f3",	--1737
		x"f3",	--1738
		x"c3",	--1739
		x"10",	--1740
		x"10",	--1741
		x"4c",	--1742
		x"4d",	--1743
		x"de",	--1744
		x"df",	--1745
		x"4a",	--1746
		x"00",	--1747
		x"4b",	--1748
		x"00",	--1749
		x"53",	--1750
		x"00",	--1751
		x"48",	--1752
		x"3f",	--1753
		x"93",	--1754
		x"23",	--1755
		x"4f",	--1756
		x"00",	--1757
		x"4f",	--1758
		x"00",	--1759
		x"00",	--1760
		x"4f",	--1761
		x"00",	--1762
		x"00",	--1763
		x"4f",	--1764
		x"00",	--1765
		x"00",	--1766
		x"4e",	--1767
		x"00",	--1768
		x"ff",	--1769
		x"00",	--1770
		x"4e",	--1771
		x"00",	--1772
		x"4d",	--1773
		x"3f",	--1774
		x"43",	--1775
		x"43",	--1776
		x"3f",	--1777
		x"e3",	--1778
		x"53",	--1779
		x"90",	--1780
		x"00",	--1781
		x"37",	--1782
		x"3f",	--1783
		x"93",	--1784
		x"2b",	--1785
		x"3f",	--1786
		x"44",	--1787
		x"45",	--1788
		x"86",	--1789
		x"77",	--1790
		x"3f",	--1791
		x"4e",	--1792
		x"3f",	--1793
		x"43",	--1794
		x"00",	--1795
		x"41",	--1796
		x"00",	--1797
		x"e3",	--1798
		x"e3",	--1799
		x"53",	--1800
		x"63",	--1801
		x"4e",	--1802
		x"00",	--1803
		x"4f",	--1804
		x"00",	--1805
		x"3f",	--1806
		x"93",	--1807
		x"27",	--1808
		x"59",	--1809
		x"00",	--1810
		x"44",	--1811
		x"00",	--1812
		x"45",	--1813
		x"00",	--1814
		x"49",	--1815
		x"f0",	--1816
		x"00",	--1817
		x"24",	--1818
		x"4d",	--1819
		x"44",	--1820
		x"45",	--1821
		x"c3",	--1822
		x"10",	--1823
		x"10",	--1824
		x"53",	--1825
		x"23",	--1826
		x"4c",	--1827
		x"00",	--1828
		x"4d",	--1829
		x"00",	--1830
		x"43",	--1831
		x"43",	--1832
		x"f0",	--1833
		x"00",	--1834
		x"24",	--1835
		x"5c",	--1836
		x"6d",	--1837
		x"53",	--1838
		x"23",	--1839
		x"53",	--1840
		x"63",	--1841
		x"f4",	--1842
		x"f5",	--1843
		x"43",	--1844
		x"43",	--1845
		x"93",	--1846
		x"20",	--1847
		x"93",	--1848
		x"20",	--1849
		x"43",	--1850
		x"43",	--1851
		x"41",	--1852
		x"00",	--1853
		x"41",	--1854
		x"00",	--1855
		x"da",	--1856
		x"db",	--1857
		x"3f",	--1858
		x"43",	--1859
		x"43",	--1860
		x"3f",	--1861
		x"92",	--1862
		x"23",	--1863
		x"9e",	--1864
		x"00",	--1865
		x"00",	--1866
		x"27",	--1867
		x"40",	--1868
		x"fb",	--1869
		x"3f",	--1870
		x"50",	--1871
		x"ff",	--1872
		x"4e",	--1873
		x"00",	--1874
		x"4f",	--1875
		x"00",	--1876
		x"4c",	--1877
		x"00",	--1878
		x"4d",	--1879
		x"00",	--1880
		x"41",	--1881
		x"50",	--1882
		x"00",	--1883
		x"41",	--1884
		x"52",	--1885
		x"12",	--1886
		x"f6",	--1887
		x"41",	--1888
		x"50",	--1889
		x"00",	--1890
		x"41",	--1891
		x"12",	--1892
		x"f6",	--1893
		x"41",	--1894
		x"52",	--1895
		x"41",	--1896
		x"50",	--1897
		x"00",	--1898
		x"41",	--1899
		x"50",	--1900
		x"00",	--1901
		x"12",	--1902
		x"ec",	--1903
		x"12",	--1904
		x"f4",	--1905
		x"50",	--1906
		x"00",	--1907
		x"41",	--1908
		x"50",	--1909
		x"ff",	--1910
		x"4e",	--1911
		x"00",	--1912
		x"4f",	--1913
		x"00",	--1914
		x"4c",	--1915
		x"00",	--1916
		x"4d",	--1917
		x"00",	--1918
		x"41",	--1919
		x"50",	--1920
		x"00",	--1921
		x"41",	--1922
		x"52",	--1923
		x"12",	--1924
		x"f6",	--1925
		x"41",	--1926
		x"50",	--1927
		x"00",	--1928
		x"41",	--1929
		x"12",	--1930
		x"f6",	--1931
		x"e3",	--1932
		x"00",	--1933
		x"41",	--1934
		x"52",	--1935
		x"41",	--1936
		x"50",	--1937
		x"00",	--1938
		x"41",	--1939
		x"50",	--1940
		x"00",	--1941
		x"12",	--1942
		x"ec",	--1943
		x"12",	--1944
		x"f4",	--1945
		x"50",	--1946
		x"00",	--1947
		x"41",	--1948
		x"12",	--1949
		x"12",	--1950
		x"12",	--1951
		x"12",	--1952
		x"12",	--1953
		x"12",	--1954
		x"12",	--1955
		x"12",	--1956
		x"50",	--1957
		x"ff",	--1958
		x"4e",	--1959
		x"00",	--1960
		x"4f",	--1961
		x"00",	--1962
		x"4c",	--1963
		x"00",	--1964
		x"4d",	--1965
		x"00",	--1966
		x"41",	--1967
		x"50",	--1968
		x"00",	--1969
		x"41",	--1970
		x"52",	--1971
		x"12",	--1972
		x"f6",	--1973
		x"41",	--1974
		x"50",	--1975
		x"00",	--1976
		x"41",	--1977
		x"12",	--1978
		x"f6",	--1979
		x"41",	--1980
		x"00",	--1981
		x"93",	--1982
		x"28",	--1983
		x"41",	--1984
		x"00",	--1985
		x"93",	--1986
		x"28",	--1987
		x"92",	--1988
		x"24",	--1989
		x"92",	--1990
		x"24",	--1991
		x"93",	--1992
		x"24",	--1993
		x"93",	--1994
		x"24",	--1995
		x"41",	--1996
		x"00",	--1997
		x"41",	--1998
		x"00",	--1999
		x"41",	--2000
		x"00",	--2001
		x"41",	--2002
		x"00",	--2003
		x"40",	--2004
		x"00",	--2005
		x"43",	--2006
		x"43",	--2007
		x"43",	--2008
		x"43",	--2009
		x"43",	--2010
		x"00",	--2011
		x"43",	--2012
		x"00",	--2013
		x"43",	--2014
		x"43",	--2015
		x"4c",	--2016
		x"00",	--2017
		x"3c",	--2018
		x"58",	--2019
		x"69",	--2020
		x"c3",	--2021
		x"10",	--2022
		x"10",	--2023
		x"53",	--2024
		x"00",	--2025
		x"24",	--2026
		x"b3",	--2027
		x"24",	--2028
		x"58",	--2029
		x"69",	--2030
		x"56",	--2031
		x"67",	--2032
		x"43",	--2033
		x"43",	--2034
		x"99",	--2035
		x"28",	--2036
		x"24",	--2037
		x"43",	--2038
		x"43",	--2039
		x"5c",	--2040
		x"6d",	--2041
		x"56",	--2042
		x"67",	--2043
		x"93",	--2044
		x"37",	--2045
		x"d3",	--2046
		x"d3",	--2047
		x"3f",	--2048
		x"98",	--2049
		x"2b",	--2050
		x"3f",	--2051
		x"4a",	--2052
		x"00",	--2053
		x"4b",	--2054
		x"00",	--2055
		x"4f",	--2056
		x"41",	--2057
		x"00",	--2058
		x"51",	--2059
		x"00",	--2060
		x"4a",	--2061
		x"53",	--2062
		x"46",	--2063
		x"00",	--2064
		x"43",	--2065
		x"91",	--2066
		x"00",	--2067
		x"00",	--2068
		x"24",	--2069
		x"4d",	--2070
		x"00",	--2071
		x"93",	--2072
		x"38",	--2073
		x"90",	--2074
		x"40",	--2075
		x"2c",	--2076
		x"41",	--2077
		x"00",	--2078
		x"53",	--2079
		x"41",	--2080
		x"00",	--2081
		x"41",	--2082
		x"00",	--2083
		x"4d",	--2084
		x"5e",	--2085
		x"6f",	--2086
		x"93",	--2087
		x"38",	--2088
		x"5a",	--2089
		x"6b",	--2090
		x"53",	--2091
		x"90",	--2092
		x"40",	--2093
		x"2b",	--2094
		x"4a",	--2095
		x"00",	--2096
		x"4b",	--2097
		x"00",	--2098
		x"4c",	--2099
		x"00",	--2100
		x"4e",	--2101
		x"4f",	--2102
		x"f0",	--2103
		x"00",	--2104
		x"f3",	--2105
		x"90",	--2106
		x"00",	--2107
		x"24",	--2108
		x"4e",	--2109
		x"00",	--2110
		x"4f",	--2111
		x"00",	--2112
		x"40",	--2113
		x"00",	--2114
		x"00",	--2115
		x"41",	--2116
		x"52",	--2117
		x"12",	--2118
		x"f4",	--2119
		x"50",	--2120
		x"00",	--2121
		x"41",	--2122
		x"41",	--2123
		x"41",	--2124
		x"41",	--2125
		x"41",	--2126
		x"41",	--2127
		x"41",	--2128
		x"41",	--2129
		x"41",	--2130
		x"d3",	--2131
		x"d3",	--2132
		x"3f",	--2133
		x"50",	--2134
		x"00",	--2135
		x"4a",	--2136
		x"b3",	--2137
		x"24",	--2138
		x"41",	--2139
		x"00",	--2140
		x"41",	--2141
		x"00",	--2142
		x"c3",	--2143
		x"10",	--2144
		x"10",	--2145
		x"4c",	--2146
		x"4d",	--2147
		x"d3",	--2148
		x"d0",	--2149
		x"80",	--2150
		x"46",	--2151
		x"00",	--2152
		x"47",	--2153
		x"00",	--2154
		x"c3",	--2155
		x"10",	--2156
		x"10",	--2157
		x"53",	--2158
		x"93",	--2159
		x"3b",	--2160
		x"48",	--2161
		x"00",	--2162
		x"3f",	--2163
		x"93",	--2164
		x"24",	--2165
		x"43",	--2166
		x"91",	--2167
		x"00",	--2168
		x"00",	--2169
		x"24",	--2170
		x"4f",	--2171
		x"00",	--2172
		x"41",	--2173
		x"50",	--2174
		x"00",	--2175
		x"3f",	--2176
		x"93",	--2177
		x"23",	--2178
		x"4e",	--2179
		x"4f",	--2180
		x"f0",	--2181
		x"00",	--2182
		x"f3",	--2183
		x"93",	--2184
		x"23",	--2185
		x"93",	--2186
		x"23",	--2187
		x"93",	--2188
		x"00",	--2189
		x"20",	--2190
		x"93",	--2191
		x"00",	--2192
		x"27",	--2193
		x"50",	--2194
		x"00",	--2195
		x"63",	--2196
		x"f0",	--2197
		x"ff",	--2198
		x"f3",	--2199
		x"3f",	--2200
		x"43",	--2201
		x"3f",	--2202
		x"43",	--2203
		x"3f",	--2204
		x"43",	--2205
		x"91",	--2206
		x"00",	--2207
		x"00",	--2208
		x"24",	--2209
		x"4f",	--2210
		x"00",	--2211
		x"41",	--2212
		x"50",	--2213
		x"00",	--2214
		x"3f",	--2215
		x"43",	--2216
		x"3f",	--2217
		x"93",	--2218
		x"23",	--2219
		x"40",	--2220
		x"fb",	--2221
		x"3f",	--2222
		x"12",	--2223
		x"12",	--2224
		x"12",	--2225
		x"12",	--2226
		x"12",	--2227
		x"50",	--2228
		x"ff",	--2229
		x"4e",	--2230
		x"00",	--2231
		x"4f",	--2232
		x"00",	--2233
		x"4c",	--2234
		x"00",	--2235
		x"4d",	--2236
		x"00",	--2237
		x"41",	--2238
		x"50",	--2239
		x"00",	--2240
		x"41",	--2241
		x"52",	--2242
		x"12",	--2243
		x"f6",	--2244
		x"41",	--2245
		x"52",	--2246
		x"41",	--2247
		x"12",	--2248
		x"f6",	--2249
		x"41",	--2250
		x"00",	--2251
		x"93",	--2252
		x"28",	--2253
		x"41",	--2254
		x"00",	--2255
		x"93",	--2256
		x"28",	--2257
		x"e1",	--2258
		x"00",	--2259
		x"00",	--2260
		x"92",	--2261
		x"24",	--2262
		x"93",	--2263
		x"24",	--2264
		x"92",	--2265
		x"24",	--2266
		x"93",	--2267
		x"24",	--2268
		x"41",	--2269
		x"00",	--2270
		x"81",	--2271
		x"00",	--2272
		x"4d",	--2273
		x"00",	--2274
		x"41",	--2275
		x"00",	--2276
		x"41",	--2277
		x"00",	--2278
		x"41",	--2279
		x"00",	--2280
		x"41",	--2281
		x"00",	--2282
		x"99",	--2283
		x"2c",	--2284
		x"5e",	--2285
		x"6f",	--2286
		x"53",	--2287
		x"4d",	--2288
		x"00",	--2289
		x"40",	--2290
		x"00",	--2291
		x"43",	--2292
		x"40",	--2293
		x"40",	--2294
		x"43",	--2295
		x"43",	--2296
		x"3c",	--2297
		x"dc",	--2298
		x"dd",	--2299
		x"88",	--2300
		x"79",	--2301
		x"c3",	--2302
		x"10",	--2303
		x"10",	--2304
		x"5e",	--2305
		x"6f",	--2306
		x"53",	--2307
		x"24",	--2308
		x"99",	--2309
		x"2b",	--2310
		x"23",	--2311
		x"98",	--2312
		x"2b",	--2313
		x"3f",	--2314
		x"9f",	--2315
		x"2b",	--2316
		x"98",	--2317
		x"2f",	--2318
		x"3f",	--2319
		x"4a",	--2320
		x"4b",	--2321
		x"f0",	--2322
		x"00",	--2323
		x"f3",	--2324
		x"90",	--2325
		x"00",	--2326
		x"24",	--2327
		x"4a",	--2328
		x"00",	--2329
		x"4b",	--2330
		x"00",	--2331
		x"41",	--2332
		x"50",	--2333
		x"00",	--2334
		x"12",	--2335
		x"f4",	--2336
		x"50",	--2337
		x"00",	--2338
		x"41",	--2339
		x"41",	--2340
		x"41",	--2341
		x"41",	--2342
		x"41",	--2343
		x"41",	--2344
		x"42",	--2345
		x"00",	--2346
		x"41",	--2347
		x"50",	--2348
		x"00",	--2349
		x"3f",	--2350
		x"9e",	--2351
		x"23",	--2352
		x"40",	--2353
		x"fb",	--2354
		x"3f",	--2355
		x"93",	--2356
		x"23",	--2357
		x"4a",	--2358
		x"4b",	--2359
		x"f0",	--2360
		x"00",	--2361
		x"f3",	--2362
		x"93",	--2363
		x"23",	--2364
		x"93",	--2365
		x"23",	--2366
		x"93",	--2367
		x"20",	--2368
		x"93",	--2369
		x"27",	--2370
		x"50",	--2371
		x"00",	--2372
		x"63",	--2373
		x"f0",	--2374
		x"ff",	--2375
		x"f3",	--2376
		x"3f",	--2377
		x"43",	--2378
		x"00",	--2379
		x"43",	--2380
		x"00",	--2381
		x"43",	--2382
		x"00",	--2383
		x"41",	--2384
		x"50",	--2385
		x"00",	--2386
		x"3f",	--2387
		x"41",	--2388
		x"52",	--2389
		x"3f",	--2390
		x"50",	--2391
		x"ff",	--2392
		x"4e",	--2393
		x"00",	--2394
		x"4f",	--2395
		x"00",	--2396
		x"4c",	--2397
		x"00",	--2398
		x"4d",	--2399
		x"00",	--2400
		x"41",	--2401
		x"50",	--2402
		x"00",	--2403
		x"41",	--2404
		x"52",	--2405
		x"12",	--2406
		x"f6",	--2407
		x"41",	--2408
		x"52",	--2409
		x"41",	--2410
		x"12",	--2411
		x"f6",	--2412
		x"93",	--2413
		x"00",	--2414
		x"28",	--2415
		x"93",	--2416
		x"00",	--2417
		x"28",	--2418
		x"41",	--2419
		x"52",	--2420
		x"41",	--2421
		x"50",	--2422
		x"00",	--2423
		x"12",	--2424
		x"f7",	--2425
		x"50",	--2426
		x"00",	--2427
		x"41",	--2428
		x"43",	--2429
		x"3f",	--2430
		x"50",	--2431
		x"ff",	--2432
		x"4e",	--2433
		x"00",	--2434
		x"4f",	--2435
		x"00",	--2436
		x"41",	--2437
		x"52",	--2438
		x"41",	--2439
		x"12",	--2440
		x"f6",	--2441
		x"41",	--2442
		x"00",	--2443
		x"93",	--2444
		x"24",	--2445
		x"28",	--2446
		x"92",	--2447
		x"24",	--2448
		x"41",	--2449
		x"00",	--2450
		x"93",	--2451
		x"38",	--2452
		x"90",	--2453
		x"00",	--2454
		x"38",	--2455
		x"93",	--2456
		x"00",	--2457
		x"20",	--2458
		x"43",	--2459
		x"40",	--2460
		x"7f",	--2461
		x"50",	--2462
		x"00",	--2463
		x"41",	--2464
		x"41",	--2465
		x"00",	--2466
		x"41",	--2467
		x"00",	--2468
		x"40",	--2469
		x"00",	--2470
		x"8d",	--2471
		x"4c",	--2472
		x"f0",	--2473
		x"00",	--2474
		x"20",	--2475
		x"93",	--2476
		x"00",	--2477
		x"27",	--2478
		x"e3",	--2479
		x"e3",	--2480
		x"53",	--2481
		x"63",	--2482
		x"50",	--2483
		x"00",	--2484
		x"41",	--2485
		x"43",	--2486
		x"43",	--2487
		x"50",	--2488
		x"00",	--2489
		x"41",	--2490
		x"c3",	--2491
		x"10",	--2492
		x"10",	--2493
		x"53",	--2494
		x"23",	--2495
		x"3f",	--2496
		x"43",	--2497
		x"40",	--2498
		x"80",	--2499
		x"50",	--2500
		x"00",	--2501
		x"41",	--2502
		x"12",	--2503
		x"12",	--2504
		x"12",	--2505
		x"12",	--2506
		x"82",	--2507
		x"4e",	--2508
		x"4f",	--2509
		x"43",	--2510
		x"00",	--2511
		x"93",	--2512
		x"20",	--2513
		x"93",	--2514
		x"20",	--2515
		x"43",	--2516
		x"00",	--2517
		x"41",	--2518
		x"12",	--2519
		x"f4",	--2520
		x"52",	--2521
		x"41",	--2522
		x"41",	--2523
		x"41",	--2524
		x"41",	--2525
		x"41",	--2526
		x"40",	--2527
		x"00",	--2528
		x"00",	--2529
		x"40",	--2530
		x"00",	--2531
		x"00",	--2532
		x"4a",	--2533
		x"00",	--2534
		x"4b",	--2535
		x"00",	--2536
		x"4a",	--2537
		x"4b",	--2538
		x"12",	--2539
		x"f4",	--2540
		x"53",	--2541
		x"93",	--2542
		x"38",	--2543
		x"27",	--2544
		x"4a",	--2545
		x"00",	--2546
		x"4b",	--2547
		x"00",	--2548
		x"4f",	--2549
		x"f0",	--2550
		x"00",	--2551
		x"20",	--2552
		x"40",	--2553
		x"00",	--2554
		x"8f",	--2555
		x"4e",	--2556
		x"00",	--2557
		x"3f",	--2558
		x"51",	--2559
		x"00",	--2560
		x"00",	--2561
		x"61",	--2562
		x"00",	--2563
		x"00",	--2564
		x"53",	--2565
		x"23",	--2566
		x"3f",	--2567
		x"4f",	--2568
		x"e3",	--2569
		x"53",	--2570
		x"43",	--2571
		x"43",	--2572
		x"4e",	--2573
		x"f0",	--2574
		x"00",	--2575
		x"24",	--2576
		x"5c",	--2577
		x"6d",	--2578
		x"53",	--2579
		x"23",	--2580
		x"53",	--2581
		x"63",	--2582
		x"fa",	--2583
		x"fb",	--2584
		x"43",	--2585
		x"43",	--2586
		x"93",	--2587
		x"20",	--2588
		x"93",	--2589
		x"20",	--2590
		x"43",	--2591
		x"43",	--2592
		x"f0",	--2593
		x"00",	--2594
		x"20",	--2595
		x"48",	--2596
		x"49",	--2597
		x"da",	--2598
		x"db",	--2599
		x"4d",	--2600
		x"00",	--2601
		x"4e",	--2602
		x"00",	--2603
		x"40",	--2604
		x"00",	--2605
		x"8f",	--2606
		x"4e",	--2607
		x"00",	--2608
		x"3f",	--2609
		x"c3",	--2610
		x"10",	--2611
		x"10",	--2612
		x"53",	--2613
		x"23",	--2614
		x"3f",	--2615
		x"12",	--2616
		x"12",	--2617
		x"12",	--2618
		x"93",	--2619
		x"2c",	--2620
		x"90",	--2621
		x"01",	--2622
		x"28",	--2623
		x"40",	--2624
		x"00",	--2625
		x"43",	--2626
		x"42",	--2627
		x"4e",	--2628
		x"4f",	--2629
		x"49",	--2630
		x"93",	--2631
		x"20",	--2632
		x"50",	--2633
		x"fb",	--2634
		x"4c",	--2635
		x"43",	--2636
		x"8e",	--2637
		x"7f",	--2638
		x"4a",	--2639
		x"41",	--2640
		x"41",	--2641
		x"41",	--2642
		x"41",	--2643
		x"90",	--2644
		x"01",	--2645
		x"28",	--2646
		x"42",	--2647
		x"43",	--2648
		x"40",	--2649
		x"00",	--2650
		x"4e",	--2651
		x"4f",	--2652
		x"49",	--2653
		x"93",	--2654
		x"27",	--2655
		x"c3",	--2656
		x"10",	--2657
		x"10",	--2658
		x"53",	--2659
		x"23",	--2660
		x"3f",	--2661
		x"40",	--2662
		x"00",	--2663
		x"43",	--2664
		x"40",	--2665
		x"00",	--2666
		x"3f",	--2667
		x"40",	--2668
		x"00",	--2669
		x"43",	--2670
		x"43",	--2671
		x"3f",	--2672
		x"12",	--2673
		x"12",	--2674
		x"12",	--2675
		x"12",	--2676
		x"12",	--2677
		x"4f",	--2678
		x"4f",	--2679
		x"00",	--2680
		x"4f",	--2681
		x"00",	--2682
		x"4d",	--2683
		x"00",	--2684
		x"4d",	--2685
		x"93",	--2686
		x"28",	--2687
		x"92",	--2688
		x"24",	--2689
		x"93",	--2690
		x"24",	--2691
		x"93",	--2692
		x"24",	--2693
		x"4d",	--2694
		x"00",	--2695
		x"90",	--2696
		x"ff",	--2697
		x"38",	--2698
		x"90",	--2699
		x"00",	--2700
		x"34",	--2701
		x"4e",	--2702
		x"4f",	--2703
		x"f0",	--2704
		x"00",	--2705
		x"f3",	--2706
		x"90",	--2707
		x"00",	--2708
		x"24",	--2709
		x"50",	--2710
		x"00",	--2711
		x"63",	--2712
		x"93",	--2713
		x"38",	--2714
		x"4b",	--2715
		x"50",	--2716
		x"00",	--2717
		x"c3",	--2718
		x"10",	--2719
		x"10",	--2720
		x"c3",	--2721
		x"10",	--2722
		x"10",	--2723
		x"c3",	--2724
		x"10",	--2725
		x"10",	--2726
		x"c3",	--2727
		x"10",	--2728
		x"10",	--2729
		x"c3",	--2730
		x"10",	--2731
		x"10",	--2732
		x"c3",	--2733
		x"10",	--2734
		x"10",	--2735
		x"c3",	--2736
		x"10",	--2737
		x"10",	--2738
		x"f3",	--2739
		x"f0",	--2740
		x"00",	--2741
		x"4d",	--2742
		x"3c",	--2743
		x"93",	--2744
		x"23",	--2745
		x"43",	--2746
		x"43",	--2747
		x"43",	--2748
		x"4d",	--2749
		x"5d",	--2750
		x"5d",	--2751
		x"5d",	--2752
		x"5d",	--2753
		x"5d",	--2754
		x"5d",	--2755
		x"5d",	--2756
		x"4f",	--2757
		x"f0",	--2758
		x"00",	--2759
		x"dd",	--2760
		x"4a",	--2761
		x"11",	--2762
		x"43",	--2763
		x"10",	--2764
		x"4c",	--2765
		x"df",	--2766
		x"4d",	--2767
		x"41",	--2768
		x"41",	--2769
		x"41",	--2770
		x"41",	--2771
		x"41",	--2772
		x"41",	--2773
		x"93",	--2774
		x"23",	--2775
		x"4e",	--2776
		x"4f",	--2777
		x"f0",	--2778
		x"00",	--2779
		x"f3",	--2780
		x"93",	--2781
		x"20",	--2782
		x"93",	--2783
		x"27",	--2784
		x"50",	--2785
		x"00",	--2786
		x"63",	--2787
		x"3f",	--2788
		x"c3",	--2789
		x"10",	--2790
		x"10",	--2791
		x"4b",	--2792
		x"50",	--2793
		x"00",	--2794
		x"3f",	--2795
		x"43",	--2796
		x"43",	--2797
		x"43",	--2798
		x"3f",	--2799
		x"d3",	--2800
		x"d0",	--2801
		x"00",	--2802
		x"f3",	--2803
		x"f0",	--2804
		x"00",	--2805
		x"43",	--2806
		x"3f",	--2807
		x"40",	--2808
		x"ff",	--2809
		x"8b",	--2810
		x"90",	--2811
		x"00",	--2812
		x"34",	--2813
		x"4e",	--2814
		x"4f",	--2815
		x"47",	--2816
		x"f0",	--2817
		x"00",	--2818
		x"24",	--2819
		x"c3",	--2820
		x"10",	--2821
		x"10",	--2822
		x"53",	--2823
		x"23",	--2824
		x"43",	--2825
		x"43",	--2826
		x"f0",	--2827
		x"00",	--2828
		x"24",	--2829
		x"58",	--2830
		x"69",	--2831
		x"53",	--2832
		x"23",	--2833
		x"53",	--2834
		x"63",	--2835
		x"fe",	--2836
		x"ff",	--2837
		x"43",	--2838
		x"43",	--2839
		x"93",	--2840
		x"20",	--2841
		x"93",	--2842
		x"20",	--2843
		x"43",	--2844
		x"43",	--2845
		x"4e",	--2846
		x"4f",	--2847
		x"dc",	--2848
		x"dd",	--2849
		x"48",	--2850
		x"49",	--2851
		x"f0",	--2852
		x"00",	--2853
		x"f3",	--2854
		x"90",	--2855
		x"00",	--2856
		x"24",	--2857
		x"50",	--2858
		x"00",	--2859
		x"63",	--2860
		x"48",	--2861
		x"49",	--2862
		x"c3",	--2863
		x"10",	--2864
		x"10",	--2865
		x"c3",	--2866
		x"10",	--2867
		x"10",	--2868
		x"c3",	--2869
		x"10",	--2870
		x"10",	--2871
		x"c3",	--2872
		x"10",	--2873
		x"10",	--2874
		x"c3",	--2875
		x"10",	--2876
		x"10",	--2877
		x"c3",	--2878
		x"10",	--2879
		x"10",	--2880
		x"c3",	--2881
		x"10",	--2882
		x"10",	--2883
		x"f3",	--2884
		x"f0",	--2885
		x"00",	--2886
		x"43",	--2887
		x"90",	--2888
		x"40",	--2889
		x"2f",	--2890
		x"43",	--2891
		x"3f",	--2892
		x"43",	--2893
		x"43",	--2894
		x"3f",	--2895
		x"93",	--2896
		x"23",	--2897
		x"48",	--2898
		x"49",	--2899
		x"f0",	--2900
		x"00",	--2901
		x"f3",	--2902
		x"93",	--2903
		x"24",	--2904
		x"50",	--2905
		x"00",	--2906
		x"63",	--2907
		x"3f",	--2908
		x"93",	--2909
		x"27",	--2910
		x"3f",	--2911
		x"12",	--2912
		x"12",	--2913
		x"4f",	--2914
		x"4f",	--2915
		x"00",	--2916
		x"f0",	--2917
		x"00",	--2918
		x"4f",	--2919
		x"00",	--2920
		x"c3",	--2921
		x"10",	--2922
		x"c3",	--2923
		x"10",	--2924
		x"c3",	--2925
		x"10",	--2926
		x"c3",	--2927
		x"10",	--2928
		x"c3",	--2929
		x"10",	--2930
		x"c3",	--2931
		x"10",	--2932
		x"c3",	--2933
		x"10",	--2934
		x"4d",	--2935
		x"4f",	--2936
		x"00",	--2937
		x"b0",	--2938
		x"00",	--2939
		x"43",	--2940
		x"6f",	--2941
		x"4f",	--2942
		x"00",	--2943
		x"93",	--2944
		x"20",	--2945
		x"93",	--2946
		x"24",	--2947
		x"40",	--2948
		x"ff",	--2949
		x"00",	--2950
		x"4a",	--2951
		x"4b",	--2952
		x"5c",	--2953
		x"6d",	--2954
		x"5c",	--2955
		x"6d",	--2956
		x"5c",	--2957
		x"6d",	--2958
		x"5c",	--2959
		x"6d",	--2960
		x"5c",	--2961
		x"6d",	--2962
		x"5c",	--2963
		x"6d",	--2964
		x"5c",	--2965
		x"6d",	--2966
		x"40",	--2967
		x"00",	--2968
		x"00",	--2969
		x"90",	--2970
		x"40",	--2971
		x"2c",	--2972
		x"40",	--2973
		x"ff",	--2974
		x"5c",	--2975
		x"6d",	--2976
		x"4f",	--2977
		x"53",	--2978
		x"90",	--2979
		x"40",	--2980
		x"2b",	--2981
		x"4a",	--2982
		x"00",	--2983
		x"4c",	--2984
		x"00",	--2985
		x"4d",	--2986
		x"00",	--2987
		x"41",	--2988
		x"41",	--2989
		x"41",	--2990
		x"90",	--2991
		x"00",	--2992
		x"24",	--2993
		x"50",	--2994
		x"ff",	--2995
		x"4d",	--2996
		x"00",	--2997
		x"40",	--2998
		x"00",	--2999
		x"00",	--3000
		x"4a",	--3001
		x"4b",	--3002
		x"5c",	--3003
		x"6d",	--3004
		x"5c",	--3005
		x"6d",	--3006
		x"5c",	--3007
		x"6d",	--3008
		x"5c",	--3009
		x"6d",	--3010
		x"5c",	--3011
		x"6d",	--3012
		x"5c",	--3013
		x"6d",	--3014
		x"5c",	--3015
		x"6d",	--3016
		x"4c",	--3017
		x"4d",	--3018
		x"d3",	--3019
		x"d0",	--3020
		x"40",	--3021
		x"4a",	--3022
		x"00",	--3023
		x"4b",	--3024
		x"00",	--3025
		x"41",	--3026
		x"41",	--3027
		x"41",	--3028
		x"93",	--3029
		x"23",	--3030
		x"43",	--3031
		x"00",	--3032
		x"41",	--3033
		x"41",	--3034
		x"41",	--3035
		x"93",	--3036
		x"24",	--3037
		x"4a",	--3038
		x"4b",	--3039
		x"f3",	--3040
		x"f0",	--3041
		x"00",	--3042
		x"93",	--3043
		x"20",	--3044
		x"93",	--3045
		x"24",	--3046
		x"43",	--3047
		x"00",	--3048
		x"3f",	--3049
		x"93",	--3050
		x"23",	--3051
		x"42",	--3052
		x"00",	--3053
		x"3f",	--3054
		x"43",	--3055
		x"00",	--3056
		x"3f",	--3057
		x"12",	--3058
		x"4f",	--3059
		x"93",	--3060
		x"28",	--3061
		x"4e",	--3062
		x"93",	--3063
		x"28",	--3064
		x"92",	--3065
		x"24",	--3066
		x"92",	--3067
		x"24",	--3068
		x"93",	--3069
		x"24",	--3070
		x"93",	--3071
		x"24",	--3072
		x"4f",	--3073
		x"00",	--3074
		x"9e",	--3075
		x"00",	--3076
		x"24",	--3077
		x"93",	--3078
		x"20",	--3079
		x"43",	--3080
		x"4e",	--3081
		x"41",	--3082
		x"41",	--3083
		x"93",	--3084
		x"24",	--3085
		x"93",	--3086
		x"00",	--3087
		x"23",	--3088
		x"43",	--3089
		x"4e",	--3090
		x"41",	--3091
		x"41",	--3092
		x"93",	--3093
		x"00",	--3094
		x"27",	--3095
		x"43",	--3096
		x"3f",	--3097
		x"4f",	--3098
		x"00",	--3099
		x"4e",	--3100
		x"00",	--3101
		x"9b",	--3102
		x"3b",	--3103
		x"9c",	--3104
		x"38",	--3105
		x"4f",	--3106
		x"00",	--3107
		x"4f",	--3108
		x"00",	--3109
		x"4e",	--3110
		x"00",	--3111
		x"4e",	--3112
		x"00",	--3113
		x"9f",	--3114
		x"2b",	--3115
		x"9e",	--3116
		x"28",	--3117
		x"9b",	--3118
		x"2b",	--3119
		x"9e",	--3120
		x"28",	--3121
		x"9f",	--3122
		x"28",	--3123
		x"9c",	--3124
		x"28",	--3125
		x"43",	--3126
		x"3f",	--3127
		x"93",	--3128
		x"23",	--3129
		x"43",	--3130
		x"3f",	--3131
		x"92",	--3132
		x"23",	--3133
		x"4e",	--3134
		x"00",	--3135
		x"4f",	--3136
		x"00",	--3137
		x"8f",	--3138
		x"3f",	--3139
		x"43",	--3140
		x"93",	--3141
		x"34",	--3142
		x"40",	--3143
		x"00",	--3144
		x"e3",	--3145
		x"53",	--3146
		x"93",	--3147
		x"34",	--3148
		x"e3",	--3149
		x"e3",	--3150
		x"53",	--3151
		x"12",	--3152
		x"12",	--3153
		x"f9",	--3154
		x"41",	--3155
		x"b3",	--3156
		x"24",	--3157
		x"e3",	--3158
		x"53",	--3159
		x"b3",	--3160
		x"24",	--3161
		x"e3",	--3162
		x"53",	--3163
		x"41",	--3164
		x"12",	--3165
		x"f8",	--3166
		x"4e",	--3167
		x"41",	--3168
		x"12",	--3169
		x"43",	--3170
		x"93",	--3171
		x"34",	--3172
		x"40",	--3173
		x"00",	--3174
		x"e3",	--3175
		x"e3",	--3176
		x"53",	--3177
		x"63",	--3178
		x"93",	--3179
		x"34",	--3180
		x"e3",	--3181
		x"e3",	--3182
		x"e3",	--3183
		x"53",	--3184
		x"63",	--3185
		x"12",	--3186
		x"f9",	--3187
		x"b3",	--3188
		x"24",	--3189
		x"e3",	--3190
		x"e3",	--3191
		x"53",	--3192
		x"63",	--3193
		x"b3",	--3194
		x"24",	--3195
		x"e3",	--3196
		x"e3",	--3197
		x"53",	--3198
		x"63",	--3199
		x"41",	--3200
		x"41",	--3201
		x"12",	--3202
		x"f8",	--3203
		x"4c",	--3204
		x"4d",	--3205
		x"41",	--3206
		x"40",	--3207
		x"00",	--3208
		x"4e",	--3209
		x"43",	--3210
		x"5f",	--3211
		x"6e",	--3212
		x"9d",	--3213
		x"28",	--3214
		x"8d",	--3215
		x"d3",	--3216
		x"83",	--3217
		x"23",	--3218
		x"41",	--3219
		x"12",	--3220
		x"f9",	--3221
		x"4e",	--3222
		x"41",	--3223
		x"12",	--3224
		x"12",	--3225
		x"12",	--3226
		x"40",	--3227
		x"00",	--3228
		x"4c",	--3229
		x"4d",	--3230
		x"43",	--3231
		x"43",	--3232
		x"5e",	--3233
		x"6f",	--3234
		x"6c",	--3235
		x"6d",	--3236
		x"9b",	--3237
		x"28",	--3238
		x"20",	--3239
		x"9a",	--3240
		x"28",	--3241
		x"8a",	--3242
		x"7b",	--3243
		x"d3",	--3244
		x"83",	--3245
		x"23",	--3246
		x"41",	--3247
		x"41",	--3248
		x"41",	--3249
		x"41",	--3250
		x"12",	--3251
		x"f9",	--3252
		x"4c",	--3253
		x"4d",	--3254
		x"41",	--3255
		x"13",	--3256
		x"d0",	--3257
		x"00",	--3258
		x"3f",	--3259
		x"61",	--3260
		x"74",	--3261
		x"6e",	--3262
		x"20",	--3263
		x"6f",	--3264
		x"20",	--3265
		x"20",	--3266
		x"65",	--3267
		x"20",	--3268
		x"62",	--3269
		x"6e",	--3270
		x"66",	--3271
		x"6c",	--3272
		x"0d",	--3273
		x"00",	--3274
		x"65",	--3275
		x"73",	--3276
		x"6f",	--3277
		x"6c",	--3278
		x"20",	--3279
		x"6f",	--3280
		x"20",	--3281
		x"65",	--3282
		x"20",	--3283
		x"68",	--3284
		x"74",	--3285
		x"0a",	--3286
		x"63",	--3287
		x"72",	--3288
		x"65",	--3289
		x"74",	--3290
		x"75",	--3291
		x"61",	--3292
		x"65",	--3293
		x"0d",	--3294
		x"00",	--3295
		x"25",	--3296
		x"20",	--3297
		x"45",	--3298
		x"54",	--3299
		x"52",	--3300
		x"47",	--3301
		x"54",	--3302
		x"0a",	--3303
		x"53",	--3304
		x"6d",	--3305
		x"74",	--3306
		x"69",	--3307
		x"67",	--3308
		x"77",	--3309
		x"6e",	--3310
		x"20",	--3311
		x"65",	--3312
		x"72",	--3313
		x"62",	--3314
		x"79",	--3315
		x"77",	--3316
		x"6f",	--3317
		x"67",	--3318
		x"0a",	--3319
		x"25",	--3320
		x"20",	--3321
		x"77",	--3322
		x"25",	--3323
		x"20",	--3324
		x"77",	--3325
		x"0a",	--3326
		x"00",	--3327
		x"e2",	--3328
		x"e3",	--3329
		x"e3",	--3330
		x"e3",	--3331
		x"e3",	--3332
		x"e3",	--3333
		x"e2",	--3334
		x"e3",	--3335
		x"0a",	--3336
		x"3d",	--3337
		x"3d",	--3338
		x"3d",	--3339
		x"4d",	--3340
		x"72",	--3341
		x"65",	--3342
		x"20",	--3343
		x"43",	--3344
		x"20",	--3345
		x"3d",	--3346
		x"3d",	--3347
		x"3d",	--3348
		x"0a",	--3349
		x"77",	--3350
		x"69",	--3351
		x"65",	--3352
		x"72",	--3353
		x"61",	--3354
		x"00",	--3355
		x"77",	--3356
		x"00",	--3357
		x"6e",	--3358
		x"6f",	--3359
		x"65",	--3360
		x"00",	--3361
		x"6f",	--3362
		x"74",	--3363
		x"6f",	--3364
		x"64",	--3365
		x"72",	--3366
		x"0d",	--3367
		x"00",	--3368
		x"20",	--3369
		x"00",	--3370
		x"63",	--3371
		x"00",	--3372
		x"72",	--3373
		x"74",	--3374
		x"0a",	--3375
		x"00",	--3376
		x"6f",	--3377
		x"72",	--3378
		x"63",	--3379
		x"20",	--3380
		x"73",	--3381
		x"67",	--3382
		x"3a",	--3383
		x"0a",	--3384
		x"09",	--3385
		x"63",	--3386
		x"52",	--3387
		x"47",	--3388
		x"53",	--3389
		x"45",	--3390
		x"20",	--3391
		x"41",	--3392
		x"55",	--3393
		x"0d",	--3394
		x"00",	--3395
		x"6f",	--3396
		x"65",	--3397
		x"68",	--3398
		x"6e",	--3399
		x"20",	--3400
		x"65",	--3401
		x"74",	--3402
		x"74",	--3403
		x"72",	--3404
		x"69",	--3405
		x"6c",	--3406
		x"20",	--3407
		x"72",	--3408
		x"6e",	--3409
		x"0d",	--3410
		x"00",	--3411
		x"3d",	--3412
		x"64",	--3413
		x"76",	--3414
		x"25",	--3415
		x"0d",	--3416
		x"00",	--3417
		x"65",	--3418
		x"64",	--3419
		x"0d",	--3420
		x"09",	--3421
		x"63",	--3422
		x"52",	--3423
		x"47",	--3424
		x"53",	--3425
		x"45",	--3426
		x"0d",	--3427
		x"00",	--3428
		x"63",	--3429
		x"69",	--3430
		x"20",	--3431
		x"6f",	--3432
		x"20",	--3433
		x"20",	--3434
		x"75",	--3435
		x"62",	--3436
		x"72",	--3437
		x"0a",	--3438
		x"25",	--3439
		x"20",	--3440
		x"73",	--3441
		x"0a",	--3442
		x"25",	--3443
		x"3a",	--3444
		x"6e",	--3445
		x"20",	--3446
		x"75",	--3447
		x"68",	--3448
		x"63",	--3449
		x"6d",	--3450
		x"61",	--3451
		x"64",	--3452
		x"0a",	--3453
		x"00",	--3454
		x"eb",	--3455
		x"ea",	--3456
		x"ea",	--3457
		x"ea",	--3458
		x"ea",	--3459
		x"ea",	--3460
		x"ea",	--3461
		x"ea",	--3462
		x"ea",	--3463
		x"ea",	--3464
		x"ea",	--3465
		x"ea",	--3466
		x"ea",	--3467
		x"ea",	--3468
		x"ea",	--3469
		x"ea",	--3470
		x"ea",	--3471
		x"ea",	--3472
		x"ea",	--3473
		x"ea",	--3474
		x"ea",	--3475
		x"ea",	--3476
		x"ea",	--3477
		x"ea",	--3478
		x"ea",	--3479
		x"ea",	--3480
		x"ea",	--3481
		x"ea",	--3482
		x"ea",	--3483
		x"eb",	--3484
		x"ea",	--3485
		x"ea",	--3486
		x"ea",	--3487
		x"ea",	--3488
		x"ea",	--3489
		x"ea",	--3490
		x"ea",	--3491
		x"ea",	--3492
		x"ea",	--3493
		x"ea",	--3494
		x"ea",	--3495
		x"ea",	--3496
		x"ea",	--3497
		x"ea",	--3498
		x"ea",	--3499
		x"ea",	--3500
		x"ea",	--3501
		x"ea",	--3502
		x"ea",	--3503
		x"ea",	--3504
		x"ea",	--3505
		x"ea",	--3506
		x"ea",	--3507
		x"ea",	--3508
		x"ea",	--3509
		x"ea",	--3510
		x"ea",	--3511
		x"ea",	--3512
		x"ea",	--3513
		x"ea",	--3514
		x"ea",	--3515
		x"ea",	--3516
		x"ea",	--3517
		x"ea",	--3518
		x"ea",	--3519
		x"ea",	--3520
		x"ea",	--3521
		x"ea",	--3522
		x"ea",	--3523
		x"ea",	--3524
		x"ea",	--3525
		x"ea",	--3526
		x"ea",	--3527
		x"ea",	--3528
		x"ea",	--3529
		x"ea",	--3530
		x"ea",	--3531
		x"ea",	--3532
		x"ea",	--3533
		x"ea",	--3534
		x"ea",	--3535
		x"ea",	--3536
		x"ea",	--3537
		x"ea",	--3538
		x"31",	--3539
		x"33",	--3540
		x"35",	--3541
		x"37",	--3542
		x"39",	--3543
		x"62",	--3544
		x"64",	--3545
		x"66",	--3546
		x"00",	--3547
		x"00",	--3548
		x"00",	--3549
		x"00",	--3550
		x"00",	--3551
		x"01",	--3552
		x"02",	--3553
		x"03",	--3554
		x"03",	--3555
		x"04",	--3556
		x"04",	--3557
		x"04",	--3558
		x"04",	--3559
		x"05",	--3560
		x"05",	--3561
		x"05",	--3562
		x"05",	--3563
		x"05",	--3564
		x"05",	--3565
		x"05",	--3566
		x"05",	--3567
		x"06",	--3568
		x"06",	--3569
		x"06",	--3570
		x"06",	--3571
		x"06",	--3572
		x"06",	--3573
		x"06",	--3574
		x"06",	--3575
		x"06",	--3576
		x"06",	--3577
		x"06",	--3578
		x"06",	--3579
		x"06",	--3580
		x"06",	--3581
		x"06",	--3582
		x"06",	--3583
		x"07",	--3584
		x"07",	--3585
		x"07",	--3586
		x"07",	--3587
		x"07",	--3588
		x"07",	--3589
		x"07",	--3590
		x"07",	--3591
		x"07",	--3592
		x"07",	--3593
		x"07",	--3594
		x"07",	--3595
		x"07",	--3596
		x"07",	--3597
		x"07",	--3598
		x"07",	--3599
		x"07",	--3600
		x"07",	--3601
		x"07",	--3602
		x"07",	--3603
		x"07",	--3604
		x"07",	--3605
		x"07",	--3606
		x"07",	--3607
		x"07",	--3608
		x"07",	--3609
		x"07",	--3610
		x"07",	--3611
		x"07",	--3612
		x"07",	--3613
		x"07",	--3614
		x"07",	--3615
		x"08",	--3616
		x"08",	--3617
		x"08",	--3618
		x"08",	--3619
		x"08",	--3620
		x"08",	--3621
		x"08",	--3622
		x"08",	--3623
		x"08",	--3624
		x"08",	--3625
		x"08",	--3626
		x"08",	--3627
		x"08",	--3628
		x"08",	--3629
		x"08",	--3630
		x"08",	--3631
		x"08",	--3632
		x"08",	--3633
		x"08",	--3634
		x"08",	--3635
		x"08",	--3636
		x"08",	--3637
		x"08",	--3638
		x"08",	--3639
		x"08",	--3640
		x"08",	--3641
		x"08",	--3642
		x"08",	--3643
		x"08",	--3644
		x"08",	--3645
		x"08",	--3646
		x"08",	--3647
		x"08",	--3648
		x"08",	--3649
		x"08",	--3650
		x"08",	--3651
		x"08",	--3652
		x"08",	--3653
		x"08",	--3654
		x"08",	--3655
		x"08",	--3656
		x"08",	--3657
		x"08",	--3658
		x"08",	--3659
		x"08",	--3660
		x"08",	--3661
		x"08",	--3662
		x"08",	--3663
		x"08",	--3664
		x"08",	--3665
		x"08",	--3666
		x"08",	--3667
		x"08",	--3668
		x"08",	--3669
		x"08",	--3670
		x"08",	--3671
		x"08",	--3672
		x"08",	--3673
		x"08",	--3674
		x"08",	--3675
		x"08",	--3676
		x"08",	--3677
		x"08",	--3678
		x"08",	--3679
		x"65",	--3680
		x"70",	--3681
		x"00",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"eb",	--4087
		x"e7",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
