library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"2e",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"0e",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"2e",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"d2",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"20",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"2e",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"0e",	--29
		x"f9",	--30
		x"31",	--31
		x"74",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"7c",	--44
		x"b0",	--45
		x"fe",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"c8",	--50
		x"b0",	--51
		x"40",	--52
		x"21",	--53
		x"3d",	--54
		x"e5",	--55
		x"3e",	--56
		x"0e",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"2e",	--61
		x"3d",	--62
		x"f6",	--63
		x"3e",	--64
		x"ae",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"2e",	--69
		x"3d",	--70
		x"fc",	--71
		x"3e",	--72
		x"22",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"2e",	--77
		x"3d",	--78
		x"01",	--79
		x"3e",	--80
		x"46",	--81
		x"7f",	--82
		x"61",	--83
		x"b0",	--84
		x"2e",	--85
		x"3d",	--86
		x"08",	--87
		x"3e",	--88
		x"c4",	--89
		x"7f",	--90
		x"70",	--91
		x"b0",	--92
		x"2e",	--93
		x"3d",	--94
		x"0c",	--95
		x"3e",	--96
		x"04",	--97
		x"7f",	--98
		x"65",	--99
		x"b0",	--100
		x"2e",	--101
		x"3d",	--102
		x"14",	--103
		x"3e",	--104
		x"ec",	--105
		x"7f",	--106
		x"73",	--107
		x"b0",	--108
		x"2e",	--109
		x"3d",	--110
		x"25",	--111
		x"3e",	--112
		x"14",	--113
		x"7f",	--114
		x"63",	--115
		x"b0",	--116
		x"2e",	--117
		x"3d",	--118
		x"39",	--119
		x"3e",	--120
		x"22",	--121
		x"7f",	--122
		x"62",	--123
		x"b0",	--124
		x"2e",	--125
		x"0e",	--126
		x"0f",	--127
		x"b0",	--128
		x"c4",	--129
		x"2c",	--130
		x"3d",	--131
		x"20",	--132
		x"3e",	--133
		x"80",	--134
		x"0f",	--135
		x"3f",	--136
		x"10",	--137
		x"b0",	--138
		x"cc",	--139
		x"0f",	--140
		x"3f",	--141
		x"10",	--142
		x"b0",	--143
		x"14",	--144
		x"2c",	--145
		x"3d",	--146
		x"20",	--147
		x"3e",	--148
		x"88",	--149
		x"0f",	--150
		x"3f",	--151
		x"06",	--152
		x"b0",	--153
		x"cc",	--154
		x"0f",	--155
		x"3f",	--156
		x"06",	--157
		x"b0",	--158
		x"14",	--159
		x"0e",	--160
		x"3e",	--161
		x"06",	--162
		x"0f",	--163
		x"3f",	--164
		x"10",	--165
		x"b0",	--166
		x"ba",	--167
		x"3e",	--168
		x"98",	--169
		x"0f",	--170
		x"2f",	--171
		x"b0",	--172
		x"22",	--173
		x"3e",	--174
		x"9c",	--175
		x"0f",	--176
		x"2f",	--177
		x"b0",	--178
		x"22",	--179
		x"0e",	--180
		x"2e",	--181
		x"0f",	--182
		x"2f",	--183
		x"b0",	--184
		x"f0",	--185
		x"0e",	--186
		x"3e",	--187
		x"06",	--188
		x"0f",	--189
		x"3f",	--190
		x"10",	--191
		x"b0",	--192
		x"fa",	--193
		x"b0",	--194
		x"fa",	--195
		x"3e",	--196
		x"a0",	--197
		x"0f",	--198
		x"b0",	--199
		x"3a",	--200
		x"0f",	--201
		x"b0",	--202
		x"40",	--203
		x"3d",	--204
		x"64",	--205
		x"3e",	--206
		x"2a",	--207
		x"0f",	--208
		x"b0",	--209
		x"4e",	--210
		x"03",	--211
		x"03",	--212
		x"30",	--213
		x"d1",	--214
		x"30",	--215
		x"17",	--216
		x"30",	--217
		x"1d",	--218
		x"30",	--219
		x"52",	--220
		x"3c",	--221
		x"32",	--222
		x"0d",	--223
		x"3d",	--224
		x"10",	--225
		x"0e",	--226
		x"3e",	--227
		x"1c",	--228
		x"0f",	--229
		x"3f",	--230
		x"4a",	--231
		x"b0",	--232
		x"dc",	--233
		x"31",	--234
		x"0c",	--235
		x"03",	--236
		x"03",	--237
		x"30",	--238
		x"d1",	--239
		x"30",	--240
		x"17",	--241
		x"30",	--242
		x"1d",	--243
		x"30",	--244
		x"52",	--245
		x"3c",	--246
		x"32",	--247
		x"0d",	--248
		x"3d",	--249
		x"0e",	--250
		x"0e",	--251
		x"3e",	--252
		x"12",	--253
		x"0f",	--254
		x"3f",	--255
		x"26",	--256
		x"b0",	--257
		x"dc",	--258
		x"31",	--259
		x"0c",	--260
		x"0e",	--261
		x"3e",	--262
		x"1a",	--263
		x"0f",	--264
		x"3f",	--265
		x"3e",	--266
		x"b0",	--267
		x"e2",	--268
		x"b0",	--269
		x"ba",	--270
		x"f2",	--271
		x"80",	--272
		x"19",	--273
		x"32",	--274
		x"0b",	--275
		x"0a",	--276
		x"05",	--277
		x"1b",	--278
		x"03",	--279
		x"2b",	--280
		x"01",	--281
		x"0b",	--282
		x"b0",	--283
		x"9a",	--284
		x"0f",	--285
		x"fc",	--286
		x"b0",	--287
		x"c2",	--288
		x"0b",	--289
		x"3e",	--290
		x"7f",	--291
		x"0d",	--292
		x"06",	--293
		x"7f",	--294
		x"1b",	--295
		x"ed",	--296
		x"7f",	--297
		x"1c",	--298
		x"12",	--299
		x"30",	--300
		x"44",	--301
		x"b0",	--302
		x"40",	--303
		x"21",	--304
		x"3f",	--305
		x"62",	--306
		x"0f",	--307
		x"0a",	--308
		x"ca",	--309
		x"00",	--310
		x"0e",	--311
		x"5f",	--312
		x"62",	--313
		x"b0",	--314
		x"62",	--315
		x"0a",	--316
		x"dd",	--317
		x"0a",	--318
		x"db",	--319
		x"3a",	--320
		x"30",	--321
		x"47",	--322
		x"b0",	--323
		x"40",	--324
		x"21",	--325
		x"d4",	--326
		x"3a",	--327
		x"28",	--328
		x"d1",	--329
		x"82",	--330
		x"10",	--331
		x"0c",	--332
		x"4e",	--333
		x"8e",	--334
		x"0e",	--335
		x"30",	--336
		x"4b",	--337
		x"81",	--338
		x"8e",	--339
		x"b0",	--340
		x"40",	--341
		x"21",	--342
		x"1f",	--343
		x"8a",	--344
		x"3e",	--345
		x"62",	--346
		x"0e",	--347
		x"0e",	--348
		x"ce",	--349
		x"00",	--350
		x"1a",	--351
		x"ba",	--352
		x"1b",	--353
		x"04",	--354
		x"7f",	--355
		x"5b",	--356
		x"b5",	--357
		x"b1",	--358
		x"2b",	--359
		x"b2",	--360
		x"7f",	--361
		x"42",	--362
		x"17",	--363
		x"7f",	--364
		x"43",	--365
		x"04",	--366
		x"7f",	--367
		x"41",	--368
		x"a8",	--369
		x"07",	--370
		x"7f",	--371
		x"43",	--372
		x"16",	--373
		x"7f",	--374
		x"44",	--375
		x"a1",	--376
		x"1b",	--377
		x"30",	--378
		x"4e",	--379
		x"b0",	--380
		x"40",	--381
		x"21",	--382
		x"b0",	--383
		x"74",	--384
		x"0b",	--385
		x"98",	--386
		x"30",	--387
		x"53",	--388
		x"b0",	--389
		x"40",	--390
		x"21",	--391
		x"b0",	--392
		x"9c",	--393
		x"0b",	--394
		x"8f",	--395
		x"30",	--396
		x"5a",	--397
		x"b0",	--398
		x"40",	--399
		x"21",	--400
		x"b0",	--401
		x"c4",	--402
		x"0b",	--403
		x"86",	--404
		x"30",	--405
		x"62",	--406
		x"b0",	--407
		x"40",	--408
		x"21",	--409
		x"b0",	--410
		x"ec",	--411
		x"0b",	--412
		x"7d",	--413
		x"30",	--414
		x"be",	--415
		x"82",	--416
		x"20",	--417
		x"30",	--418
		x"0b",	--419
		x"0a",	--420
		x"21",	--421
		x"0a",	--422
		x"0b",	--423
		x"2f",	--424
		x"1b",	--425
		x"0e",	--426
		x"1f",	--427
		x"02",	--428
		x"b0",	--429
		x"7e",	--430
		x"0d",	--431
		x"2a",	--432
		x"18",	--433
		x"0e",	--434
		x"1f",	--435
		x"04",	--436
		x"81",	--437
		x"02",	--438
		x"b0",	--439
		x"7e",	--440
		x"0e",	--441
		x"1d",	--442
		x"02",	--443
		x"1f",	--444
		x"20",	--445
		x"b0",	--446
		x"4e",	--447
		x"0f",	--448
		x"21",	--449
		x"3a",	--450
		x"3b",	--451
		x"30",	--452
		x"3d",	--453
		x"64",	--454
		x"3e",	--455
		x"2a",	--456
		x"f2",	--457
		x"3e",	--458
		x"2a",	--459
		x"ef",	--460
		x"0e",	--461
		x"1f",	--462
		x"24",	--463
		x"b0",	--464
		x"66",	--465
		x"0e",	--466
		x"1f",	--467
		x"22",	--468
		x"b0",	--469
		x"66",	--470
		x"30",	--471
		x"c6",	--472
		x"b0",	--473
		x"40",	--474
		x"21",	--475
		x"30",	--476
		x"b2",	--477
		x"00",	--478
		x"09",	--479
		x"1f",	--480
		x"24",	--481
		x"b0",	--482
		x"22",	--483
		x"1f",	--484
		x"22",	--485
		x"b0",	--486
		x"22",	--487
		x"30",	--488
		x"0e",	--489
		x"3f",	--490
		x"9a",	--491
		x"b0",	--492
		x"0a",	--493
		x"82",	--494
		x"00",	--495
		x"ef",	--496
		x"82",	--497
		x"24",	--498
		x"82",	--499
		x"22",	--500
		x"30",	--501
		x"0b",	--502
		x"0a",	--503
		x"21",	--504
		x"0b",	--505
		x"3f",	--506
		x"03",	--507
		x"30",	--508
		x"23",	--509
		x"0e",	--510
		x"1f",	--511
		x"02",	--512
		x"b0",	--513
		x"4c",	--514
		x"0a",	--515
		x"0e",	--516
		x"1f",	--517
		x"04",	--518
		x"b0",	--519
		x"4c",	--520
		x"0b",	--521
		x"0f",	--522
		x"0a",	--523
		x"30",	--524
		x"f9",	--525
		x"b0",	--526
		x"40",	--527
		x"31",	--528
		x"06",	--529
		x"0e",	--530
		x"1f",	--531
		x"24",	--532
		x"b0",	--533
		x"66",	--534
		x"0e",	--535
		x"1f",	--536
		x"22",	--537
		x"b0",	--538
		x"66",	--539
		x"0f",	--540
		x"21",	--541
		x"3a",	--542
		x"3b",	--543
		x"30",	--544
		x"0e",	--545
		x"1f",	--546
		x"06",	--547
		x"b0",	--548
		x"7e",	--549
		x"1d",	--550
		x"0e",	--551
		x"1f",	--552
		x"00",	--553
		x"b0",	--554
		x"4e",	--555
		x"d1",	--556
		x"30",	--557
		x"cd",	--558
		x"b0",	--559
		x"40",	--560
		x"a1",	--561
		x"00",	--562
		x"30",	--563
		x"de",	--564
		x"b0",	--565
		x"40",	--566
		x"21",	--567
		x"3f",	--568
		x"e3",	--569
		x"3e",	--570
		x"9c",	--571
		x"1f",	--572
		x"24",	--573
		x"b0",	--574
		x"66",	--575
		x"3e",	--576
		x"64",	--577
		x"1f",	--578
		x"22",	--579
		x"b0",	--580
		x"66",	--581
		x"1d",	--582
		x"3e",	--583
		x"c8",	--584
		x"1f",	--585
		x"00",	--586
		x"b0",	--587
		x"4e",	--588
		x"30",	--589
		x"3e",	--590
		x"64",	--591
		x"1f",	--592
		x"24",	--593
		x"b0",	--594
		x"66",	--595
		x"3e",	--596
		x"9c",	--597
		x"1f",	--598
		x"22",	--599
		x"b0",	--600
		x"66",	--601
		x"1d",	--602
		x"3e",	--603
		x"c8",	--604
		x"1f",	--605
		x"00",	--606
		x"b0",	--607
		x"4e",	--608
		x"30",	--609
		x"3e",	--610
		x"c4",	--611
		x"1f",	--612
		x"24",	--613
		x"b0",	--614
		x"66",	--615
		x"3e",	--616
		x"c4",	--617
		x"1f",	--618
		x"22",	--619
		x"b0",	--620
		x"66",	--621
		x"1d",	--622
		x"3e",	--623
		x"c8",	--624
		x"1f",	--625
		x"00",	--626
		x"b0",	--627
		x"4e",	--628
		x"30",	--629
		x"3e",	--630
		x"3c",	--631
		x"1f",	--632
		x"24",	--633
		x"b0",	--634
		x"66",	--635
		x"3e",	--636
		x"3c",	--637
		x"1f",	--638
		x"22",	--639
		x"b0",	--640
		x"66",	--641
		x"1d",	--642
		x"3e",	--643
		x"c8",	--644
		x"1f",	--645
		x"00",	--646
		x"b0",	--647
		x"4e",	--648
		x"30",	--649
		x"30",	--650
		x"01",	--651
		x"b0",	--652
		x"40",	--653
		x"21",	--654
		x"0f",	--655
		x"30",	--656
		x"b2",	--657
		x"00",	--658
		x"92",	--659
		x"b2",	--660
		x"30",	--661
		x"94",	--662
		x"b2",	--663
		x"41",	--664
		x"96",	--665
		x"30",	--666
		x"17",	--667
		x"b0",	--668
		x"40",	--669
		x"92",	--670
		x"90",	--671
		x"b1",	--672
		x"35",	--673
		x"00",	--674
		x"b0",	--675
		x"40",	--676
		x"21",	--677
		x"0f",	--678
		x"30",	--679
		x"0b",	--680
		x"0a",	--681
		x"09",	--682
		x"09",	--683
		x"1f",	--684
		x"1a",	--685
		x"b0",	--686
		x"2a",	--687
		x"0a",	--688
		x"0b",	--689
		x"1e",	--690
		x"1c",	--691
		x"1f",	--692
		x"1e",	--693
		x"b0",	--694
		x"c4",	--695
		x"89",	--696
		x"1c",	--697
		x"89",	--698
		x"1e",	--699
		x"0d",	--700
		x"0e",	--701
		x"0f",	--702
		x"b0",	--703
		x"10",	--704
		x"0c",	--705
		x"3d",	--706
		x"00",	--707
		x"b0",	--708
		x"c4",	--709
		x"0a",	--710
		x"0b",	--711
		x"3c",	--712
		x"66",	--713
		x"3d",	--714
		x"66",	--715
		x"b0",	--716
		x"d4",	--717
		x"0f",	--718
		x"01",	--719
		x"18",	--720
		x"3c",	--721
		x"cd",	--722
		x"3d",	--723
		x"cc",	--724
		x"0e",	--725
		x"0f",	--726
		x"b0",	--727
		x"74",	--728
		x"0f",	--729
		x"04",	--730
		x"3a",	--731
		x"cd",	--732
		x"3b",	--733
		x"cc",	--734
		x"0d",	--735
		x"0e",	--736
		x"1f",	--737
		x"18",	--738
		x"b0",	--739
		x"68",	--740
		x"39",	--741
		x"3a",	--742
		x"3b",	--743
		x"30",	--744
		x"3a",	--745
		x"66",	--746
		x"3b",	--747
		x"66",	--748
		x"f1",	--749
		x"0b",	--750
		x"0a",	--751
		x"0b",	--752
		x"0a",	--753
		x"8f",	--754
		x"18",	--755
		x"8f",	--756
		x"1a",	--757
		x"11",	--758
		x"12",	--759
		x"11",	--760
		x"12",	--761
		x"11",	--762
		x"12",	--763
		x"11",	--764
		x"12",	--765
		x"1d",	--766
		x"0e",	--767
		x"1e",	--768
		x"10",	--769
		x"b0",	--770
		x"94",	--771
		x"31",	--772
		x"8b",	--773
		x"20",	--774
		x"0e",	--775
		x"3f",	--776
		x"50",	--777
		x"b0",	--778
		x"0a",	--779
		x"8b",	--780
		x"22",	--781
		x"3a",	--782
		x"3b",	--783
		x"30",	--784
		x"0b",	--785
		x"0b",	--786
		x"1f",	--787
		x"1a",	--788
		x"b0",	--789
		x"2a",	--790
		x"8b",	--791
		x"1c",	--792
		x"8b",	--793
		x"1e",	--794
		x"0d",	--795
		x"1e",	--796
		x"20",	--797
		x"1f",	--798
		x"22",	--799
		x"b0",	--800
		x"4e",	--801
		x"3b",	--802
		x"30",	--803
		x"0b",	--804
		x"0b",	--805
		x"0d",	--806
		x"3e",	--807
		x"00",	--808
		x"1f",	--809
		x"18",	--810
		x"b0",	--811
		x"68",	--812
		x"1f",	--813
		x"22",	--814
		x"b0",	--815
		x"76",	--816
		x"3b",	--817
		x"30",	--818
		x"0b",	--819
		x"0b",	--820
		x"0d",	--821
		x"8d",	--822
		x"8d",	--823
		x"8d",	--824
		x"8d",	--825
		x"0f",	--826
		x"b0",	--827
		x"c4",	--828
		x"0d",	--829
		x"0e",	--830
		x"0f",	--831
		x"b0",	--832
		x"06",	--833
		x"3b",	--834
		x"30",	--835
		x"0b",	--836
		x"0a",	--837
		x"0a",	--838
		x"3b",	--839
		x"00",	--840
		x"0d",	--841
		x"0e",	--842
		x"1f",	--843
		x"68",	--844
		x"b0",	--845
		x"68",	--846
		x"0d",	--847
		x"0e",	--848
		x"1f",	--849
		x"66",	--850
		x"b0",	--851
		x"68",	--852
		x"30",	--853
		x"4e",	--854
		x"b0",	--855
		x"40",	--856
		x"21",	--857
		x"3a",	--858
		x"3b",	--859
		x"30",	--860
		x"82",	--861
		x"68",	--862
		x"82",	--863
		x"66",	--864
		x"30",	--865
		x"0b",	--866
		x"0a",	--867
		x"21",	--868
		x"0a",	--869
		x"0b",	--870
		x"b2",	--871
		x"02",	--872
		x"4e",	--873
		x"3a",	--874
		x"03",	--875
		x"53",	--876
		x"3e",	--877
		x"0e",	--878
		x"1f",	--879
		x"02",	--880
		x"b0",	--881
		x"7e",	--882
		x"0a",	--883
		x"0e",	--884
		x"1f",	--885
		x"04",	--886
		x"b0",	--887
		x"7e",	--888
		x"0b",	--889
		x"0f",	--890
		x"0a",	--891
		x"30",	--892
		x"9b",	--893
		x"b0",	--894
		x"40",	--895
		x"31",	--896
		x"06",	--897
		x"0e",	--898
		x"0f",	--899
		x"b0",	--900
		x"fa",	--901
		x"0c",	--902
		x"3d",	--903
		x"c8",	--904
		x"b0",	--905
		x"84",	--906
		x"0c",	--907
		x"0d",	--908
		x"0e",	--909
		x"3f",	--910
		x"80",	--911
		x"b0",	--912
		x"10",	--913
		x"0d",	--914
		x"0e",	--915
		x"1f",	--916
		x"68",	--917
		x"b0",	--918
		x"68",	--919
		x"0e",	--920
		x"0f",	--921
		x"b0",	--922
		x"fa",	--923
		x"0c",	--924
		x"3d",	--925
		x"c8",	--926
		x"b0",	--927
		x"84",	--928
		x"0d",	--929
		x"0e",	--930
		x"1f",	--931
		x"66",	--932
		x"b0",	--933
		x"68",	--934
		x"0f",	--935
		x"21",	--936
		x"3a",	--937
		x"3b",	--938
		x"30",	--939
		x"0e",	--940
		x"1f",	--941
		x"06",	--942
		x"b0",	--943
		x"7e",	--944
		x"1d",	--945
		x"0e",	--946
		x"1f",	--947
		x"02",	--948
		x"b0",	--949
		x"4e",	--950
		x"b6",	--951
		x"0e",	--952
		x"3f",	--953
		x"88",	--954
		x"b0",	--955
		x"0a",	--956
		x"82",	--957
		x"02",	--958
		x"aa",	--959
		x"30",	--960
		x"55",	--961
		x"b0",	--962
		x"40",	--963
		x"b1",	--964
		x"6f",	--965
		x"00",	--966
		x"b0",	--967
		x"40",	--968
		x"a1",	--969
		x"00",	--970
		x"30",	--971
		x"80",	--972
		x"b0",	--973
		x"40",	--974
		x"21",	--975
		x"3f",	--976
		x"d6",	--977
		x"0b",	--978
		x"0a",	--979
		x"1f",	--980
		x"6c",	--981
		x"b0",	--982
		x"2a",	--983
		x"0a",	--984
		x"0b",	--985
		x"1f",	--986
		x"6a",	--987
		x"b0",	--988
		x"2a",	--989
		x"0b",	--990
		x"0a",	--991
		x"3e",	--992
		x"3f",	--993
		x"1e",	--994
		x"0f",	--995
		x"0f",	--996
		x"0e",	--997
		x"30",	--998
		x"a3",	--999
		x"30",	--1000
		x"26",	--1001
		x"b0",	--1002
		x"52",	--1003
		x"31",	--1004
		x"0c",	--1005
		x"30",	--1006
		x"26",	--1007
		x"30",	--1008
		x"ab",	--1009
		x"b0",	--1010
		x"40",	--1011
		x"21",	--1012
		x"3a",	--1013
		x"3b",	--1014
		x"30",	--1015
		x"82",	--1016
		x"6a",	--1017
		x"82",	--1018
		x"6c",	--1019
		x"30",	--1020
		x"82",	--1021
		x"68",	--1022
		x"82",	--1023
		x"66",	--1024
		x"30",	--1025
		x"0b",	--1026
		x"0a",	--1027
		x"09",	--1028
		x"08",	--1029
		x"21",	--1030
		x"0a",	--1031
		x"0b",	--1032
		x"81",	--1033
		x"00",	--1034
		x"1f",	--1035
		x"1c",	--1036
		x"b2",	--1037
		x"04",	--1038
		x"6f",	--1039
		x"92",	--1040
		x"0e",	--1041
		x"0e",	--1042
		x"1f",	--1043
		x"02",	--1044
		x"b0",	--1045
		x"7e",	--1046
		x"08",	--1047
		x"3a",	--1048
		x"03",	--1049
		x"1e",	--1050
		x"09",	--1051
		x"0d",	--1052
		x"0e",	--1053
		x"1f",	--1054
		x"04",	--1055
		x"b0",	--1056
		x"4e",	--1057
		x"0f",	--1058
		x"21",	--1059
		x"38",	--1060
		x"39",	--1061
		x"3a",	--1062
		x"3b",	--1063
		x"30",	--1064
		x"82",	--1065
		x"0e",	--1066
		x"49",	--1067
		x"82",	--1068
		x"0e",	--1069
		x"1f",	--1070
		x"04",	--1071
		x"b0",	--1072
		x"76",	--1073
		x"0f",	--1074
		x"21",	--1075
		x"38",	--1076
		x"39",	--1077
		x"3a",	--1078
		x"3b",	--1079
		x"30",	--1080
		x"0e",	--1081
		x"1f",	--1082
		x"04",	--1083
		x"b0",	--1084
		x"7e",	--1085
		x"09",	--1086
		x"3a",	--1087
		x"05",	--1088
		x"da",	--1089
		x"0e",	--1090
		x"1f",	--1091
		x"06",	--1092
		x"b0",	--1093
		x"7e",	--1094
		x"0a",	--1095
		x"0e",	--1096
		x"1f",	--1097
		x"08",	--1098
		x"b0",	--1099
		x"7e",	--1100
		x"0b",	--1101
		x"0f",	--1102
		x"0a",	--1103
		x"30",	--1104
		x"b0",	--1105
		x"b0",	--1106
		x"40",	--1107
		x"31",	--1108
		x"06",	--1109
		x"0e",	--1110
		x"0f",	--1111
		x"b0",	--1112
		x"fa",	--1113
		x"0c",	--1114
		x"3d",	--1115
		x"c8",	--1116
		x"b0",	--1117
		x"84",	--1118
		x"0d",	--1119
		x"0e",	--1120
		x"1f",	--1121
		x"68",	--1122
		x"b0",	--1123
		x"68",	--1124
		x"0e",	--1125
		x"0f",	--1126
		x"b0",	--1127
		x"fa",	--1128
		x"0c",	--1129
		x"3d",	--1130
		x"c8",	--1131
		x"b0",	--1132
		x"84",	--1133
		x"0d",	--1134
		x"0e",	--1135
		x"1f",	--1136
		x"66",	--1137
		x"b0",	--1138
		x"68",	--1139
		x"a7",	--1140
		x"0f",	--1141
		x"b0",	--1142
		x"a4",	--1143
		x"0f",	--1144
		x"21",	--1145
		x"38",	--1146
		x"39",	--1147
		x"3a",	--1148
		x"3b",	--1149
		x"30",	--1150
		x"0e",	--1151
		x"3f",	--1152
		x"a4",	--1153
		x"b0",	--1154
		x"0a",	--1155
		x"82",	--1156
		x"04",	--1157
		x"89",	--1158
		x"1f",	--1159
		x"82",	--1160
		x"10",	--1161
		x"01",	--1162
		x"0f",	--1163
		x"82",	--1164
		x"10",	--1165
		x"0f",	--1166
		x"30",	--1167
		x"5e",	--1168
		x"19",	--1169
		x"4e",	--1170
		x"0f",	--1171
		x"03",	--1172
		x"c2",	--1173
		x"19",	--1174
		x"30",	--1175
		x"c2",	--1176
		x"19",	--1177
		x"30",	--1178
		x"1e",	--1179
		x"12",	--1180
		x"3e",	--1181
		x"06",	--1182
		x"0f",	--1183
		x"0f",	--1184
		x"10",	--1185
		x"b8",	--1186
		x"c2",	--1187
		x"19",	--1188
		x"3e",	--1189
		x"07",	--1190
		x"03",	--1191
		x"82",	--1192
		x"12",	--1193
		x"30",	--1194
		x"1e",	--1195
		x"82",	--1196
		x"12",	--1197
		x"30",	--1198
		x"f2",	--1199
		x"0e",	--1200
		x"19",	--1201
		x"f2",	--1202
		x"f2",	--1203
		x"0a",	--1204
		x"19",	--1205
		x"ee",	--1206
		x"e2",	--1207
		x"19",	--1208
		x"eb",	--1209
		x"f2",	--1210
		x"0d",	--1211
		x"19",	--1212
		x"e7",	--1213
		x"f2",	--1214
		x"09",	--1215
		x"19",	--1216
		x"e3",	--1217
		x"f2",	--1218
		x"03",	--1219
		x"19",	--1220
		x"df",	--1221
		x"f2",	--1222
		x"07",	--1223
		x"19",	--1224
		x"db",	--1225
		x"8f",	--1226
		x"00",	--1227
		x"8f",	--1228
		x"02",	--1229
		x"9f",	--1230
		x"02",	--1231
		x"04",	--1232
		x"9f",	--1233
		x"04",	--1234
		x"06",	--1235
		x"9f",	--1236
		x"06",	--1237
		x"08",	--1238
		x"9f",	--1239
		x"08",	--1240
		x"0a",	--1241
		x"8f",	--1242
		x"0c",	--1243
		x"8f",	--1244
		x"0e",	--1245
		x"8f",	--1246
		x"10",	--1247
		x"8f",	--1248
		x"12",	--1249
		x"8f",	--1250
		x"14",	--1251
		x"8f",	--1252
		x"16",	--1253
		x"30",	--1254
		x"8f",	--1255
		x"0c",	--1256
		x"8f",	--1257
		x"0e",	--1258
		x"8f",	--1259
		x"10",	--1260
		x"8f",	--1261
		x"12",	--1262
		x"8f",	--1263
		x"14",	--1264
		x"8f",	--1265
		x"16",	--1266
		x"30",	--1267
		x"8f",	--1268
		x"00",	--1269
		x"8f",	--1270
		x"02",	--1271
		x"30",	--1272
		x"8f",	--1273
		x"04",	--1274
		x"8f",	--1275
		x"06",	--1276
		x"30",	--1277
		x"8f",	--1278
		x"08",	--1279
		x"8f",	--1280
		x"0a",	--1281
		x"30",	--1282
		x"8f",	--1283
		x"0c",	--1284
		x"8f",	--1285
		x"0e",	--1286
		x"30",	--1287
		x"0b",	--1288
		x"09",	--1289
		x"08",	--1290
		x"07",	--1291
		x"06",	--1292
		x"05",	--1293
		x"04",	--1294
		x"0b",	--1295
		x"0c",	--1296
		x"0d",	--1297
		x"1e",	--1298
		x"0c",	--1299
		x"1f",	--1300
		x"0e",	--1301
		x"b0",	--1302
		x"10",	--1303
		x"08",	--1304
		x"09",	--1305
		x"1c",	--1306
		x"10",	--1307
		x"1d",	--1308
		x"12",	--1309
		x"b0",	--1310
		x"c4",	--1311
		x"06",	--1312
		x"07",	--1313
		x"8b",	--1314
		x"10",	--1315
		x"8b",	--1316
		x"12",	--1317
		x"2c",	--1318
		x"1d",	--1319
		x"02",	--1320
		x"0e",	--1321
		x"0f",	--1322
		x"b0",	--1323
		x"60",	--1324
		x"04",	--1325
		x"05",	--1326
		x"1c",	--1327
		x"04",	--1328
		x"1d",	--1329
		x"06",	--1330
		x"0e",	--1331
		x"0f",	--1332
		x"b0",	--1333
		x"60",	--1334
		x"0c",	--1335
		x"0d",	--1336
		x"b0",	--1337
		x"c4",	--1338
		x"06",	--1339
		x"07",	--1340
		x"1c",	--1341
		x"14",	--1342
		x"1d",	--1343
		x"16",	--1344
		x"0e",	--1345
		x"0f",	--1346
		x"b0",	--1347
		x"10",	--1348
		x"1c",	--1349
		x"08",	--1350
		x"1d",	--1351
		x"0a",	--1352
		x"b0",	--1353
		x"60",	--1354
		x"0c",	--1355
		x"0d",	--1356
		x"b0",	--1357
		x"c4",	--1358
		x"34",	--1359
		x"35",	--1360
		x"36",	--1361
		x"37",	--1362
		x"38",	--1363
		x"39",	--1364
		x"3b",	--1365
		x"30",	--1366
		x"0b",	--1367
		x"0a",	--1368
		x"21",	--1369
		x"0a",	--1370
		x"0b",	--1371
		x"30",	--1372
		x"6a",	--1373
		x"b0",	--1374
		x"40",	--1375
		x"21",	--1376
		x"3a",	--1377
		x"03",	--1378
		x"1b",	--1379
		x"0e",	--1380
		x"1f",	--1381
		x"02",	--1382
		x"b0",	--1383
		x"7e",	--1384
		x"0a",	--1385
		x"0e",	--1386
		x"1f",	--1387
		x"04",	--1388
		x"b0",	--1389
		x"7e",	--1390
		x"0b",	--1391
		x"0f",	--1392
		x"0a",	--1393
		x"30",	--1394
		x"b2",	--1395
		x"b0",	--1396
		x"40",	--1397
		x"31",	--1398
		x"06",	--1399
		x"8a",	--1400
		x"00",	--1401
		x"0f",	--1402
		x"21",	--1403
		x"3a",	--1404
		x"3b",	--1405
		x"30",	--1406
		x"30",	--1407
		x"72",	--1408
		x"b0",	--1409
		x"40",	--1410
		x"b1",	--1411
		x"8c",	--1412
		x"00",	--1413
		x"b0",	--1414
		x"40",	--1415
		x"a1",	--1416
		x"00",	--1417
		x"30",	--1418
		x"9d",	--1419
		x"b0",	--1420
		x"40",	--1421
		x"21",	--1422
		x"3f",	--1423
		x"ea",	--1424
		x"0b",	--1425
		x"21",	--1426
		x"0b",	--1427
		x"1f",	--1428
		x"17",	--1429
		x"16",	--1430
		x"30",	--1431
		x"cd",	--1432
		x"b0",	--1433
		x"40",	--1434
		x"21",	--1435
		x"0e",	--1436
		x"1f",	--1437
		x"02",	--1438
		x"b0",	--1439
		x"7e",	--1440
		x"2f",	--1441
		x"0f",	--1442
		x"30",	--1443
		x"b2",	--1444
		x"b0",	--1445
		x"40",	--1446
		x"31",	--1447
		x"06",	--1448
		x"0f",	--1449
		x"21",	--1450
		x"3b",	--1451
		x"30",	--1452
		x"30",	--1453
		x"72",	--1454
		x"b0",	--1455
		x"40",	--1456
		x"b1",	--1457
		x"8c",	--1458
		x"00",	--1459
		x"b0",	--1460
		x"40",	--1461
		x"a1",	--1462
		x"00",	--1463
		x"30",	--1464
		x"be",	--1465
		x"b0",	--1466
		x"40",	--1467
		x"21",	--1468
		x"3f",	--1469
		x"eb",	--1470
		x"0b",	--1471
		x"0a",	--1472
		x"8e",	--1473
		x"00",	--1474
		x"6d",	--1475
		x"4d",	--1476
		x"5e",	--1477
		x"1f",	--1478
		x"0a",	--1479
		x"0c",	--1480
		x"0f",	--1481
		x"7b",	--1482
		x"0a",	--1483
		x"2b",	--1484
		x"0c",	--1485
		x"0c",	--1486
		x"0c",	--1487
		x"0c",	--1488
		x"8d",	--1489
		x"0c",	--1490
		x"3c",	--1491
		x"d0",	--1492
		x"1a",	--1493
		x"7d",	--1494
		x"4d",	--1495
		x"17",	--1496
		x"7d",	--1497
		x"78",	--1498
		x"1a",	--1499
		x"4b",	--1500
		x"7b",	--1501
		x"d0",	--1502
		x"0a",	--1503
		x"e9",	--1504
		x"7b",	--1505
		x"0a",	--1506
		x"34",	--1507
		x"0c",	--1508
		x"0b",	--1509
		x"0b",	--1510
		x"0b",	--1511
		x"0c",	--1512
		x"8d",	--1513
		x"0c",	--1514
		x"3c",	--1515
		x"d0",	--1516
		x"7d",	--1517
		x"4d",	--1518
		x"e9",	--1519
		x"9e",	--1520
		x"00",	--1521
		x"0f",	--1522
		x"3a",	--1523
		x"3b",	--1524
		x"30",	--1525
		x"1a",	--1526
		x"de",	--1527
		x"4b",	--1528
		x"7b",	--1529
		x"9f",	--1530
		x"7b",	--1531
		x"06",	--1532
		x"0a",	--1533
		x"0c",	--1534
		x"0c",	--1535
		x"0c",	--1536
		x"0c",	--1537
		x"8d",	--1538
		x"0c",	--1539
		x"3c",	--1540
		x"a9",	--1541
		x"1a",	--1542
		x"ce",	--1543
		x"4b",	--1544
		x"7b",	--1545
		x"bf",	--1546
		x"7b",	--1547
		x"06",	--1548
		x"0a",	--1549
		x"0c",	--1550
		x"0c",	--1551
		x"0c",	--1552
		x"0c",	--1553
		x"8d",	--1554
		x"0c",	--1555
		x"3c",	--1556
		x"c9",	--1557
		x"1a",	--1558
		x"be",	--1559
		x"8d",	--1560
		x"0d",	--1561
		x"30",	--1562
		x"d4",	--1563
		x"b0",	--1564
		x"40",	--1565
		x"21",	--1566
		x"0c",	--1567
		x"0f",	--1568
		x"3a",	--1569
		x"3b",	--1570
		x"30",	--1571
		x"0c",	--1572
		x"ca",	--1573
		x"0b",	--1574
		x"0a",	--1575
		x"8e",	--1576
		x"00",	--1577
		x"6b",	--1578
		x"4b",	--1579
		x"37",	--1580
		x"1f",	--1581
		x"1a",	--1582
		x"0c",	--1583
		x"12",	--1584
		x"4d",	--1585
		x"7d",	--1586
		x"d0",	--1587
		x"7d",	--1588
		x"0a",	--1589
		x"22",	--1590
		x"0c",	--1591
		x"0d",	--1592
		x"0d",	--1593
		x"0d",	--1594
		x"0c",	--1595
		x"8b",	--1596
		x"0c",	--1597
		x"3c",	--1598
		x"d0",	--1599
		x"7b",	--1600
		x"4b",	--1601
		x"07",	--1602
		x"7b",	--1603
		x"2d",	--1604
		x"eb",	--1605
		x"3a",	--1606
		x"7b",	--1607
		x"4b",	--1608
		x"f9",	--1609
		x"02",	--1610
		x"32",	--1611
		x"03",	--1612
		x"82",	--1613
		x"32",	--1614
		x"82",	--1615
		x"38",	--1616
		x"1f",	--1617
		x"3a",	--1618
		x"32",	--1619
		x"9e",	--1620
		x"00",	--1621
		x"3a",	--1622
		x"3b",	--1623
		x"30",	--1624
		x"8b",	--1625
		x"0b",	--1626
		x"30",	--1627
		x"d4",	--1628
		x"b0",	--1629
		x"40",	--1630
		x"21",	--1631
		x"0f",	--1632
		x"3a",	--1633
		x"3b",	--1634
		x"30",	--1635
		x"0f",	--1636
		x"ee",	--1637
		x"0b",	--1638
		x"0a",	--1639
		x"0b",	--1640
		x"0a",	--1641
		x"8f",	--1642
		x"00",	--1643
		x"8f",	--1644
		x"02",	--1645
		x"8f",	--1646
		x"04",	--1647
		x"0c",	--1648
		x"0d",	--1649
		x"3e",	--1650
		x"00",	--1651
		x"3f",	--1652
		x"6e",	--1653
		x"b0",	--1654
		x"60",	--1655
		x"8b",	--1656
		x"02",	--1657
		x"02",	--1658
		x"32",	--1659
		x"03",	--1660
		x"82",	--1661
		x"32",	--1662
		x"b2",	--1663
		x"18",	--1664
		x"38",	--1665
		x"9b",	--1666
		x"3a",	--1667
		x"06",	--1668
		x"32",	--1669
		x"0f",	--1670
		x"3a",	--1671
		x"3b",	--1672
		x"30",	--1673
		x"0b",	--1674
		x"09",	--1675
		x"08",	--1676
		x"8f",	--1677
		x"06",	--1678
		x"bf",	--1679
		x"00",	--1680
		x"08",	--1681
		x"2b",	--1682
		x"1e",	--1683
		x"02",	--1684
		x"0f",	--1685
		x"b0",	--1686
		x"fa",	--1687
		x"0c",	--1688
		x"3d",	--1689
		x"00",	--1690
		x"b0",	--1691
		x"60",	--1692
		x"08",	--1693
		x"09",	--1694
		x"1e",	--1695
		x"06",	--1696
		x"0f",	--1697
		x"b0",	--1698
		x"fa",	--1699
		x"0c",	--1700
		x"0d",	--1701
		x"0e",	--1702
		x"0f",	--1703
		x"b0",	--1704
		x"10",	--1705
		x"b0",	--1706
		x"f0",	--1707
		x"8b",	--1708
		x"04",	--1709
		x"9b",	--1710
		x"00",	--1711
		x"38",	--1712
		x"39",	--1713
		x"3b",	--1714
		x"30",	--1715
		x"0b",	--1716
		x"0a",	--1717
		x"09",	--1718
		x"0a",	--1719
		x"0b",	--1720
		x"8f",	--1721
		x"06",	--1722
		x"8f",	--1723
		x"08",	--1724
		x"29",	--1725
		x"1e",	--1726
		x"02",	--1727
		x"0f",	--1728
		x"b0",	--1729
		x"fa",	--1730
		x"0c",	--1731
		x"0d",	--1732
		x"0e",	--1733
		x"0f",	--1734
		x"b0",	--1735
		x"60",	--1736
		x"0a",	--1737
		x"0b",	--1738
		x"1e",	--1739
		x"06",	--1740
		x"0f",	--1741
		x"b0",	--1742
		x"fa",	--1743
		x"0c",	--1744
		x"0d",	--1745
		x"0e",	--1746
		x"0f",	--1747
		x"b0",	--1748
		x"10",	--1749
		x"b0",	--1750
		x"f0",	--1751
		x"89",	--1752
		x"04",	--1753
		x"39",	--1754
		x"3a",	--1755
		x"3b",	--1756
		x"30",	--1757
		x"2f",	--1758
		x"8f",	--1759
		x"04",	--1760
		x"30",	--1761
		x"0b",	--1762
		x"0a",	--1763
		x"92",	--1764
		x"14",	--1765
		x"14",	--1766
		x"3b",	--1767
		x"72",	--1768
		x"0a",	--1769
		x"2b",	--1770
		x"5f",	--1771
		x"fc",	--1772
		x"8f",	--1773
		x"0f",	--1774
		x"30",	--1775
		x"e9",	--1776
		x"b0",	--1777
		x"40",	--1778
		x"31",	--1779
		x"06",	--1780
		x"1a",	--1781
		x"3b",	--1782
		x"06",	--1783
		x"1a",	--1784
		x"14",	--1785
		x"ef",	--1786
		x"0f",	--1787
		x"3a",	--1788
		x"3b",	--1789
		x"30",	--1790
		x"1e",	--1791
		x"14",	--1792
		x"3e",	--1793
		x"20",	--1794
		x"12",	--1795
		x"0f",	--1796
		x"0f",	--1797
		x"0f",	--1798
		x"0f",	--1799
		x"3f",	--1800
		x"6e",	--1801
		x"ff",	--1802
		x"68",	--1803
		x"00",	--1804
		x"bf",	--1805
		x"c4",	--1806
		x"02",	--1807
		x"bf",	--1808
		x"06",	--1809
		x"04",	--1810
		x"1e",	--1811
		x"82",	--1812
		x"14",	--1813
		x"30",	--1814
		x"0b",	--1815
		x"1b",	--1816
		x"14",	--1817
		x"3b",	--1818
		x"20",	--1819
		x"12",	--1820
		x"0c",	--1821
		x"0c",	--1822
		x"0c",	--1823
		x"0c",	--1824
		x"3c",	--1825
		x"6e",	--1826
		x"cc",	--1827
		x"00",	--1828
		x"8c",	--1829
		x"02",	--1830
		x"8c",	--1831
		x"04",	--1832
		x"1b",	--1833
		x"82",	--1834
		x"14",	--1835
		x"0f",	--1836
		x"3b",	--1837
		x"30",	--1838
		x"3f",	--1839
		x"fc",	--1840
		x"0b",	--1841
		x"31",	--1842
		x"f0",	--1843
		x"1b",	--1844
		x"14",	--1845
		x"1b",	--1846
		x"0f",	--1847
		x"5f",	--1848
		x"6e",	--1849
		x"16",	--1850
		x"3d",	--1851
		x"74",	--1852
		x"0c",	--1853
		x"05",	--1854
		x"3d",	--1855
		x"06",	--1856
		x"cd",	--1857
		x"fa",	--1858
		x"0e",	--1859
		x"1c",	--1860
		x"0c",	--1861
		x"f8",	--1862
		x"30",	--1863
		x"f1",	--1864
		x"b0",	--1865
		x"40",	--1866
		x"21",	--1867
		x"3f",	--1868
		x"31",	--1869
		x"10",	--1870
		x"3b",	--1871
		x"30",	--1872
		x"0c",	--1873
		x"81",	--1874
		x"00",	--1875
		x"6d",	--1876
		x"4d",	--1877
		x"24",	--1878
		x"1e",	--1879
		x"1f",	--1880
		x"06",	--1881
		x"6d",	--1882
		x"4d",	--1883
		x"11",	--1884
		x"1e",	--1885
		x"3f",	--1886
		x"0e",	--1887
		x"7d",	--1888
		x"20",	--1889
		x"f7",	--1890
		x"ce",	--1891
		x"ff",	--1892
		x"0d",	--1893
		x"0d",	--1894
		x"0d",	--1895
		x"8d",	--1896
		x"00",	--1897
		x"1f",	--1898
		x"6d",	--1899
		x"4d",	--1900
		x"ef",	--1901
		x"0e",	--1902
		x"0e",	--1903
		x"0c",	--1904
		x"0c",	--1905
		x"3c",	--1906
		x"6e",	--1907
		x"0e",	--1908
		x"9c",	--1909
		x"02",	--1910
		x"31",	--1911
		x"10",	--1912
		x"3b",	--1913
		x"30",	--1914
		x"1f",	--1915
		x"f1",	--1916
		x"b2",	--1917
		x"d2",	--1918
		x"60",	--1919
		x"b2",	--1920
		x"b8",	--1921
		x"72",	--1922
		x"0f",	--1923
		x"30",	--1924
		x"0b",	--1925
		x"0b",	--1926
		x"1f",	--1927
		x"16",	--1928
		x"3f",	--1929
		x"20",	--1930
		x"19",	--1931
		x"0c",	--1932
		x"0c",	--1933
		x"0d",	--1934
		x"0d",	--1935
		x"0d",	--1936
		x"0d",	--1937
		x"0d",	--1938
		x"3d",	--1939
		x"2e",	--1940
		x"8d",	--1941
		x"00",	--1942
		x"8d",	--1943
		x"02",	--1944
		x"8d",	--1945
		x"08",	--1946
		x"8d",	--1947
		x"0a",	--1948
		x"8d",	--1949
		x"0c",	--1950
		x"0e",	--1951
		x"1e",	--1952
		x"82",	--1953
		x"16",	--1954
		x"3b",	--1955
		x"30",	--1956
		x"3f",	--1957
		x"fc",	--1958
		x"0f",	--1959
		x"0c",	--1960
		x"0c",	--1961
		x"0c",	--1962
		x"0c",	--1963
		x"0c",	--1964
		x"3c",	--1965
		x"2e",	--1966
		x"8c",	--1967
		x"02",	--1968
		x"8c",	--1969
		x"04",	--1970
		x"8c",	--1971
		x"06",	--1972
		x"8c",	--1973
		x"08",	--1974
		x"9c",	--1975
		x"00",	--1976
		x"0f",	--1977
		x"30",	--1978
		x"0f",	--1979
		x"0e",	--1980
		x"0e",	--1981
		x"0e",	--1982
		x"0e",	--1983
		x"0e",	--1984
		x"8e",	--1985
		x"2e",	--1986
		x"0f",	--1987
		x"30",	--1988
		x"0f",	--1989
		x"0e",	--1990
		x"0d",	--1991
		x"0c",	--1992
		x"0b",	--1993
		x"0a",	--1994
		x"09",	--1995
		x"08",	--1996
		x"07",	--1997
		x"92",	--1998
		x"16",	--1999
		x"33",	--2000
		x"3a",	--2001
		x"2e",	--2002
		x"0b",	--2003
		x"2b",	--2004
		x"08",	--2005
		x"38",	--2006
		x"07",	--2007
		x"37",	--2008
		x"06",	--2009
		x"09",	--2010
		x"0f",	--2011
		x"1f",	--2012
		x"8b",	--2013
		x"00",	--2014
		x"19",	--2015
		x"3a",	--2016
		x"0e",	--2017
		x"3b",	--2018
		x"0e",	--2019
		x"38",	--2020
		x"0e",	--2021
		x"37",	--2022
		x"0e",	--2023
		x"19",	--2024
		x"16",	--2025
		x"19",	--2026
		x"8a",	--2027
		x"00",	--2028
		x"f1",	--2029
		x"2f",	--2030
		x"1f",	--2031
		x"02",	--2032
		x"ea",	--2033
		x"8b",	--2034
		x"00",	--2035
		x"1f",	--2036
		x"0a",	--2037
		x"9b",	--2038
		x"08",	--2039
		x"88",	--2040
		x"00",	--2041
		x"e4",	--2042
		x"2f",	--2043
		x"1f",	--2044
		x"87",	--2045
		x"00",	--2046
		x"2f",	--2047
		x"de",	--2048
		x"8a",	--2049
		x"00",	--2050
		x"db",	--2051
		x"b2",	--2052
		x"fe",	--2053
		x"60",	--2054
		x"37",	--2055
		x"38",	--2056
		x"39",	--2057
		x"3a",	--2058
		x"3b",	--2059
		x"3c",	--2060
		x"3d",	--2061
		x"3e",	--2062
		x"3f",	--2063
		x"00",	--2064
		x"8f",	--2065
		x"00",	--2066
		x"0f",	--2067
		x"30",	--2068
		x"2f",	--2069
		x"2e",	--2070
		x"1f",	--2071
		x"02",	--2072
		x"30",	--2073
		x"8f",	--2074
		x"00",	--2075
		x"30",	--2076
		x"8f",	--2077
		x"00",	--2078
		x"3f",	--2079
		x"34",	--2080
		x"b0",	--2081
		x"0a",	--2082
		x"82",	--2083
		x"0c",	--2084
		x"0f",	--2085
		x"30",	--2086
		x"0c",	--2087
		x"2f",	--2088
		x"8f",	--2089
		x"00",	--2090
		x"1d",	--2091
		x"0e",	--2092
		x"1f",	--2093
		x"0c",	--2094
		x"b0",	--2095
		x"4e",	--2096
		x"30",	--2097
		x"5e",	--2098
		x"81",	--2099
		x"3e",	--2100
		x"fc",	--2101
		x"c2",	--2102
		x"84",	--2103
		x"0f",	--2104
		x"30",	--2105
		x"3f",	--2106
		x"0f",	--2107
		x"5f",	--2108
		x"b0",	--2109
		x"8f",	--2110
		x"b0",	--2111
		x"64",	--2112
		x"30",	--2113
		x"0b",	--2114
		x"0b",	--2115
		x"0e",	--2116
		x"0e",	--2117
		x"0e",	--2118
		x"0e",	--2119
		x"0e",	--2120
		x"0f",	--2121
		x"b0",	--2122
		x"74",	--2123
		x"0f",	--2124
		x"b0",	--2125
		x"74",	--2126
		x"3b",	--2127
		x"30",	--2128
		x"0b",	--2129
		x"0a",	--2130
		x"0a",	--2131
		x"3b",	--2132
		x"07",	--2133
		x"0e",	--2134
		x"4d",	--2135
		x"7d",	--2136
		x"0f",	--2137
		x"03",	--2138
		x"0e",	--2139
		x"7d",	--2140
		x"fd",	--2141
		x"1e",	--2142
		x"0a",	--2143
		x"3f",	--2144
		x"31",	--2145
		x"b0",	--2146
		x"64",	--2147
		x"3b",	--2148
		x"3b",	--2149
		x"ef",	--2150
		x"3a",	--2151
		x"3b",	--2152
		x"30",	--2153
		x"3f",	--2154
		x"30",	--2155
		x"f5",	--2156
		x"0b",	--2157
		x"0b",	--2158
		x"0e",	--2159
		x"8e",	--2160
		x"8e",	--2161
		x"0f",	--2162
		x"b0",	--2163
		x"84",	--2164
		x"0f",	--2165
		x"b0",	--2166
		x"84",	--2167
		x"3b",	--2168
		x"30",	--2169
		x"0b",	--2170
		x"0a",	--2171
		x"0a",	--2172
		x"0b",	--2173
		x"0d",	--2174
		x"8d",	--2175
		x"8d",	--2176
		x"0f",	--2177
		x"b0",	--2178
		x"84",	--2179
		x"0f",	--2180
		x"b0",	--2181
		x"84",	--2182
		x"0c",	--2183
		x"0d",	--2184
		x"8d",	--2185
		x"8c",	--2186
		x"4d",	--2187
		x"0d",	--2188
		x"0f",	--2189
		x"b0",	--2190
		x"84",	--2191
		x"0f",	--2192
		x"b0",	--2193
		x"84",	--2194
		x"3a",	--2195
		x"3b",	--2196
		x"30",	--2197
		x"0b",	--2198
		x"0a",	--2199
		x"09",	--2200
		x"0a",	--2201
		x"0e",	--2202
		x"19",	--2203
		x"09",	--2204
		x"39",	--2205
		x"0b",	--2206
		x"0d",	--2207
		x"0d",	--2208
		x"6f",	--2209
		x"8f",	--2210
		x"b0",	--2211
		x"84",	--2212
		x"0b",	--2213
		x"0e",	--2214
		x"1b",	--2215
		x"3b",	--2216
		x"07",	--2217
		x"05",	--2218
		x"3f",	--2219
		x"20",	--2220
		x"b0",	--2221
		x"64",	--2222
		x"ef",	--2223
		x"3f",	--2224
		x"3a",	--2225
		x"b0",	--2226
		x"64",	--2227
		x"ea",	--2228
		x"39",	--2229
		x"3a",	--2230
		x"3b",	--2231
		x"30",	--2232
		x"0b",	--2233
		x"0a",	--2234
		x"09",	--2235
		x"0a",	--2236
		x"0e",	--2237
		x"17",	--2238
		x"09",	--2239
		x"39",	--2240
		x"0b",	--2241
		x"6f",	--2242
		x"8f",	--2243
		x"b0",	--2244
		x"74",	--2245
		x"0b",	--2246
		x"0e",	--2247
		x"1b",	--2248
		x"3b",	--2249
		x"07",	--2250
		x"f6",	--2251
		x"3f",	--2252
		x"20",	--2253
		x"b0",	--2254
		x"64",	--2255
		x"6f",	--2256
		x"8f",	--2257
		x"b0",	--2258
		x"74",	--2259
		x"0b",	--2260
		x"f2",	--2261
		x"39",	--2262
		x"3a",	--2263
		x"3b",	--2264
		x"30",	--2265
		x"0b",	--2266
		x"0a",	--2267
		x"09",	--2268
		x"31",	--2269
		x"ec",	--2270
		x"0b",	--2271
		x"0f",	--2272
		x"34",	--2273
		x"3b",	--2274
		x"0a",	--2275
		x"38",	--2276
		x"09",	--2277
		x"0a",	--2278
		x"0a",	--2279
		x"3e",	--2280
		x"0a",	--2281
		x"0f",	--2282
		x"b0",	--2283
		x"18",	--2284
		x"7f",	--2285
		x"30",	--2286
		x"ca",	--2287
		x"00",	--2288
		x"19",	--2289
		x"3e",	--2290
		x"0a",	--2291
		x"0f",	--2292
		x"b0",	--2293
		x"e6",	--2294
		x"0b",	--2295
		x"3f",	--2296
		x"0a",	--2297
		x"eb",	--2298
		x"0a",	--2299
		x"1a",	--2300
		x"09",	--2301
		x"3e",	--2302
		x"0a",	--2303
		x"0f",	--2304
		x"b0",	--2305
		x"18",	--2306
		x"7f",	--2307
		x"30",	--2308
		x"c9",	--2309
		x"00",	--2310
		x"3a",	--2311
		x"0f",	--2312
		x"0f",	--2313
		x"6f",	--2314
		x"8f",	--2315
		x"b0",	--2316
		x"64",	--2317
		x"0a",	--2318
		x"f7",	--2319
		x"31",	--2320
		x"14",	--2321
		x"39",	--2322
		x"3a",	--2323
		x"3b",	--2324
		x"30",	--2325
		x"3f",	--2326
		x"2d",	--2327
		x"b0",	--2328
		x"64",	--2329
		x"3b",	--2330
		x"1b",	--2331
		x"c5",	--2332
		x"1a",	--2333
		x"09",	--2334
		x"dd",	--2335
		x"0b",	--2336
		x"0a",	--2337
		x"09",	--2338
		x"0b",	--2339
		x"3b",	--2340
		x"39",	--2341
		x"6f",	--2342
		x"4f",	--2343
		x"0b",	--2344
		x"1a",	--2345
		x"8f",	--2346
		x"b0",	--2347
		x"64",	--2348
		x"0a",	--2349
		x"09",	--2350
		x"19",	--2351
		x"5f",	--2352
		x"01",	--2353
		x"4f",	--2354
		x"10",	--2355
		x"7f",	--2356
		x"25",	--2357
		x"f3",	--2358
		x"0a",	--2359
		x"1a",	--2360
		x"5f",	--2361
		x"01",	--2362
		x"7f",	--2363
		x"db",	--2364
		x"7f",	--2365
		x"54",	--2366
		x"ee",	--2367
		x"4f",	--2368
		x"0f",	--2369
		x"10",	--2370
		x"08",	--2371
		x"39",	--2372
		x"3a",	--2373
		x"3b",	--2374
		x"30",	--2375
		x"09",	--2376
		x"29",	--2377
		x"1e",	--2378
		x"02",	--2379
		x"2f",	--2380
		x"b0",	--2381
		x"2c",	--2382
		x"0b",	--2383
		x"dd",	--2384
		x"09",	--2385
		x"29",	--2386
		x"2f",	--2387
		x"b0",	--2388
		x"da",	--2389
		x"0b",	--2390
		x"d6",	--2391
		x"0f",	--2392
		x"2b",	--2393
		x"29",	--2394
		x"6f",	--2395
		x"4f",	--2396
		x"d0",	--2397
		x"19",	--2398
		x"8f",	--2399
		x"b0",	--2400
		x"64",	--2401
		x"7f",	--2402
		x"4f",	--2403
		x"fa",	--2404
		x"c8",	--2405
		x"09",	--2406
		x"29",	--2407
		x"1e",	--2408
		x"02",	--2409
		x"2f",	--2410
		x"b0",	--2411
		x"72",	--2412
		x"0b",	--2413
		x"bf",	--2414
		x"09",	--2415
		x"29",	--2416
		x"2e",	--2417
		x"0f",	--2418
		x"8f",	--2419
		x"8f",	--2420
		x"8f",	--2421
		x"8f",	--2422
		x"b0",	--2423
		x"f4",	--2424
		x"0b",	--2425
		x"b3",	--2426
		x"09",	--2427
		x"29",	--2428
		x"2f",	--2429
		x"b0",	--2430
		x"b4",	--2431
		x"0b",	--2432
		x"ac",	--2433
		x"09",	--2434
		x"29",	--2435
		x"2f",	--2436
		x"b0",	--2437
		x"64",	--2438
		x"0b",	--2439
		x"a5",	--2440
		x"09",	--2441
		x"29",	--2442
		x"2f",	--2443
		x"b0",	--2444
		x"84",	--2445
		x"0b",	--2446
		x"9e",	--2447
		x"09",	--2448
		x"29",	--2449
		x"2f",	--2450
		x"b0",	--2451
		x"a2",	--2452
		x"0b",	--2453
		x"97",	--2454
		x"3f",	--2455
		x"25",	--2456
		x"b0",	--2457
		x"64",	--2458
		x"92",	--2459
		x"0f",	--2460
		x"0e",	--2461
		x"1f",	--2462
		x"18",	--2463
		x"df",	--2464
		x"85",	--2465
		x"ee",	--2466
		x"1f",	--2467
		x"18",	--2468
		x"3f",	--2469
		x"3f",	--2470
		x"13",	--2471
		x"92",	--2472
		x"18",	--2473
		x"1e",	--2474
		x"18",	--2475
		x"1f",	--2476
		x"1a",	--2477
		x"0e",	--2478
		x"02",	--2479
		x"92",	--2480
		x"1a",	--2481
		x"f2",	--2482
		x"10",	--2483
		x"81",	--2484
		x"3e",	--2485
		x"3f",	--2486
		x"b1",	--2487
		x"f0",	--2488
		x"00",	--2489
		x"00",	--2490
		x"82",	--2491
		x"18",	--2492
		x"ec",	--2493
		x"0c",	--2494
		x"0d",	--2495
		x"3e",	--2496
		x"00",	--2497
		x"3f",	--2498
		x"6e",	--2499
		x"b0",	--2500
		x"20",	--2501
		x"3e",	--2502
		x"82",	--2503
		x"82",	--2504
		x"f2",	--2505
		x"11",	--2506
		x"80",	--2507
		x"30",	--2508
		x"1e",	--2509
		x"18",	--2510
		x"1f",	--2511
		x"1a",	--2512
		x"0e",	--2513
		x"05",	--2514
		x"1f",	--2515
		x"18",	--2516
		x"1f",	--2517
		x"1a",	--2518
		x"30",	--2519
		x"1d",	--2520
		x"18",	--2521
		x"1e",	--2522
		x"1a",	--2523
		x"3f",	--2524
		x"40",	--2525
		x"0f",	--2526
		x"0f",	--2527
		x"30",	--2528
		x"1f",	--2529
		x"1a",	--2530
		x"5f",	--2531
		x"ee",	--2532
		x"1d",	--2533
		x"1a",	--2534
		x"1e",	--2535
		x"18",	--2536
		x"0d",	--2537
		x"0b",	--2538
		x"1e",	--2539
		x"1a",	--2540
		x"3e",	--2541
		x"3f",	--2542
		x"03",	--2543
		x"82",	--2544
		x"1a",	--2545
		x"30",	--2546
		x"92",	--2547
		x"1a",	--2548
		x"30",	--2549
		x"4f",	--2550
		x"30",	--2551
		x"0b",	--2552
		x"0a",	--2553
		x"0a",	--2554
		x"0b",	--2555
		x"0c",	--2556
		x"3d",	--2557
		x"00",	--2558
		x"b0",	--2559
		x"24",	--2560
		x"0f",	--2561
		x"07",	--2562
		x"0e",	--2563
		x"0f",	--2564
		x"b0",	--2565
		x"6a",	--2566
		x"3a",	--2567
		x"3b",	--2568
		x"30",	--2569
		x"0c",	--2570
		x"3d",	--2571
		x"00",	--2572
		x"0e",	--2573
		x"0f",	--2574
		x"b0",	--2575
		x"10",	--2576
		x"b0",	--2577
		x"6a",	--2578
		x"0e",	--2579
		x"3f",	--2580
		x"00",	--2581
		x"3a",	--2582
		x"3b",	--2583
		x"30",	--2584
		x"0b",	--2585
		x"0a",	--2586
		x"09",	--2587
		x"08",	--2588
		x"07",	--2589
		x"06",	--2590
		x"05",	--2591
		x"04",	--2592
		x"31",	--2593
		x"fa",	--2594
		x"08",	--2595
		x"6b",	--2596
		x"6b",	--2597
		x"67",	--2598
		x"6c",	--2599
		x"6c",	--2600
		x"e9",	--2601
		x"6b",	--2602
		x"02",	--2603
		x"30",	--2604
		x"b2",	--2605
		x"6c",	--2606
		x"e3",	--2607
		x"6c",	--2608
		x"bb",	--2609
		x"6b",	--2610
		x"df",	--2611
		x"91",	--2612
		x"02",	--2613
		x"00",	--2614
		x"1b",	--2615
		x"02",	--2616
		x"14",	--2617
		x"04",	--2618
		x"15",	--2619
		x"06",	--2620
		x"16",	--2621
		x"04",	--2622
		x"17",	--2623
		x"06",	--2624
		x"2c",	--2625
		x"0c",	--2626
		x"09",	--2627
		x"0c",	--2628
		x"bf",	--2629
		x"39",	--2630
		x"20",	--2631
		x"50",	--2632
		x"1c",	--2633
		x"d7",	--2634
		x"81",	--2635
		x"02",	--2636
		x"81",	--2637
		x"04",	--2638
		x"4c",	--2639
		x"7c",	--2640
		x"1f",	--2641
		x"0b",	--2642
		x"0a",	--2643
		x"0b",	--2644
		x"12",	--2645
		x"0b",	--2646
		x"0a",	--2647
		x"7c",	--2648
		x"fb",	--2649
		x"81",	--2650
		x"02",	--2651
		x"81",	--2652
		x"04",	--2653
		x"1c",	--2654
		x"0d",	--2655
		x"79",	--2656
		x"1f",	--2657
		x"04",	--2658
		x"0c",	--2659
		x"0d",	--2660
		x"79",	--2661
		x"fc",	--2662
		x"3c",	--2663
		x"3d",	--2664
		x"0c",	--2665
		x"0d",	--2666
		x"1a",	--2667
		x"0b",	--2668
		x"0c",	--2669
		x"02",	--2670
		x"0d",	--2671
		x"e5",	--2672
		x"16",	--2673
		x"02",	--2674
		x"17",	--2675
		x"04",	--2676
		x"06",	--2677
		x"07",	--2678
		x"5f",	--2679
		x"01",	--2680
		x"5f",	--2681
		x"01",	--2682
		x"28",	--2683
		x"c8",	--2684
		x"01",	--2685
		x"a8",	--2686
		x"02",	--2687
		x"0e",	--2688
		x"0f",	--2689
		x"0e",	--2690
		x"0f",	--2691
		x"88",	--2692
		x"04",	--2693
		x"88",	--2694
		x"06",	--2695
		x"f8",	--2696
		x"03",	--2697
		x"00",	--2698
		x"0f",	--2699
		x"4d",	--2700
		x"0f",	--2701
		x"31",	--2702
		x"06",	--2703
		x"34",	--2704
		x"35",	--2705
		x"36",	--2706
		x"37",	--2707
		x"38",	--2708
		x"39",	--2709
		x"3a",	--2710
		x"3b",	--2711
		x"30",	--2712
		x"2b",	--2713
		x"67",	--2714
		x"81",	--2715
		x"00",	--2716
		x"04",	--2717
		x"05",	--2718
		x"5f",	--2719
		x"01",	--2720
		x"5f",	--2721
		x"01",	--2722
		x"d8",	--2723
		x"4f",	--2724
		x"68",	--2725
		x"0e",	--2726
		x"0f",	--2727
		x"0e",	--2728
		x"0f",	--2729
		x"0f",	--2730
		x"69",	--2731
		x"c8",	--2732
		x"01",	--2733
		x"a8",	--2734
		x"02",	--2735
		x"88",	--2736
		x"04",	--2737
		x"88",	--2738
		x"06",	--2739
		x"0c",	--2740
		x"0d",	--2741
		x"3c",	--2742
		x"3d",	--2743
		x"3d",	--2744
		x"ff",	--2745
		x"05",	--2746
		x"3d",	--2747
		x"00",	--2748
		x"17",	--2749
		x"3c",	--2750
		x"15",	--2751
		x"1b",	--2752
		x"02",	--2753
		x"3b",	--2754
		x"0e",	--2755
		x"0f",	--2756
		x"0a",	--2757
		x"3b",	--2758
		x"0c",	--2759
		x"0d",	--2760
		x"3c",	--2761
		x"3d",	--2762
		x"3d",	--2763
		x"ff",	--2764
		x"f5",	--2765
		x"3c",	--2766
		x"88",	--2767
		x"04",	--2768
		x"88",	--2769
		x"06",	--2770
		x"88",	--2771
		x"02",	--2772
		x"f8",	--2773
		x"03",	--2774
		x"00",	--2775
		x"0f",	--2776
		x"b3",	--2777
		x"0c",	--2778
		x"0d",	--2779
		x"1c",	--2780
		x"0d",	--2781
		x"12",	--2782
		x"0f",	--2783
		x"0e",	--2784
		x"0a",	--2785
		x"0b",	--2786
		x"0a",	--2787
		x"0b",	--2788
		x"88",	--2789
		x"04",	--2790
		x"88",	--2791
		x"06",	--2792
		x"98",	--2793
		x"02",	--2794
		x"0f",	--2795
		x"a1",	--2796
		x"6b",	--2797
		x"9f",	--2798
		x"ad",	--2799
		x"00",	--2800
		x"9d",	--2801
		x"02",	--2802
		x"02",	--2803
		x"9d",	--2804
		x"04",	--2805
		x"04",	--2806
		x"9d",	--2807
		x"06",	--2808
		x"06",	--2809
		x"5e",	--2810
		x"01",	--2811
		x"5e",	--2812
		x"01",	--2813
		x"cd",	--2814
		x"01",	--2815
		x"0f",	--2816
		x"8c",	--2817
		x"06",	--2818
		x"07",	--2819
		x"9a",	--2820
		x"39",	--2821
		x"19",	--2822
		x"39",	--2823
		x"20",	--2824
		x"8f",	--2825
		x"3e",	--2826
		x"3c",	--2827
		x"b6",	--2828
		x"c1",	--2829
		x"0e",	--2830
		x"0f",	--2831
		x"0e",	--2832
		x"0f",	--2833
		x"97",	--2834
		x"0f",	--2835
		x"79",	--2836
		x"d8",	--2837
		x"01",	--2838
		x"a8",	--2839
		x"02",	--2840
		x"3e",	--2841
		x"3f",	--2842
		x"1e",	--2843
		x"0f",	--2844
		x"88",	--2845
		x"04",	--2846
		x"88",	--2847
		x"06",	--2848
		x"92",	--2849
		x"0c",	--2850
		x"7b",	--2851
		x"81",	--2852
		x"00",	--2853
		x"81",	--2854
		x"02",	--2855
		x"81",	--2856
		x"04",	--2857
		x"4d",	--2858
		x"7d",	--2859
		x"1f",	--2860
		x"0c",	--2861
		x"4b",	--2862
		x"0c",	--2863
		x"0d",	--2864
		x"12",	--2865
		x"0d",	--2866
		x"0c",	--2867
		x"7b",	--2868
		x"fb",	--2869
		x"81",	--2870
		x"02",	--2871
		x"81",	--2872
		x"04",	--2873
		x"1c",	--2874
		x"0d",	--2875
		x"79",	--2876
		x"1f",	--2877
		x"04",	--2878
		x"0c",	--2879
		x"0d",	--2880
		x"79",	--2881
		x"fc",	--2882
		x"3c",	--2883
		x"3d",	--2884
		x"0c",	--2885
		x"0d",	--2886
		x"1a",	--2887
		x"0b",	--2888
		x"0c",	--2889
		x"04",	--2890
		x"0d",	--2891
		x"02",	--2892
		x"0a",	--2893
		x"0b",	--2894
		x"14",	--2895
		x"02",	--2896
		x"15",	--2897
		x"04",	--2898
		x"04",	--2899
		x"05",	--2900
		x"49",	--2901
		x"0a",	--2902
		x"0b",	--2903
		x"18",	--2904
		x"6c",	--2905
		x"33",	--2906
		x"df",	--2907
		x"01",	--2908
		x"01",	--2909
		x"2f",	--2910
		x"3f",	--2911
		x"c2",	--2912
		x"2c",	--2913
		x"31",	--2914
		x"e0",	--2915
		x"81",	--2916
		x"04",	--2917
		x"81",	--2918
		x"06",	--2919
		x"81",	--2920
		x"00",	--2921
		x"81",	--2922
		x"02",	--2923
		x"0e",	--2924
		x"3e",	--2925
		x"18",	--2926
		x"0f",	--2927
		x"2f",	--2928
		x"b0",	--2929
		x"2c",	--2930
		x"0e",	--2931
		x"3e",	--2932
		x"10",	--2933
		x"0f",	--2934
		x"b0",	--2935
		x"2c",	--2936
		x"0d",	--2937
		x"3d",	--2938
		x"0e",	--2939
		x"3e",	--2940
		x"10",	--2941
		x"0f",	--2942
		x"3f",	--2943
		x"18",	--2944
		x"b0",	--2945
		x"32",	--2946
		x"b0",	--2947
		x"4e",	--2948
		x"31",	--2949
		x"20",	--2950
		x"30",	--2951
		x"31",	--2952
		x"e0",	--2953
		x"81",	--2954
		x"04",	--2955
		x"81",	--2956
		x"06",	--2957
		x"81",	--2958
		x"00",	--2959
		x"81",	--2960
		x"02",	--2961
		x"0e",	--2962
		x"3e",	--2963
		x"18",	--2964
		x"0f",	--2965
		x"2f",	--2966
		x"b0",	--2967
		x"2c",	--2968
		x"0e",	--2969
		x"3e",	--2970
		x"10",	--2971
		x"0f",	--2972
		x"b0",	--2973
		x"2c",	--2974
		x"d1",	--2975
		x"11",	--2976
		x"0d",	--2977
		x"3d",	--2978
		x"0e",	--2979
		x"3e",	--2980
		x"10",	--2981
		x"0f",	--2982
		x"3f",	--2983
		x"18",	--2984
		x"b0",	--2985
		x"32",	--2986
		x"b0",	--2987
		x"4e",	--2988
		x"31",	--2989
		x"20",	--2990
		x"30",	--2991
		x"0b",	--2992
		x"0a",	--2993
		x"09",	--2994
		x"08",	--2995
		x"07",	--2996
		x"06",	--2997
		x"05",	--2998
		x"04",	--2999
		x"31",	--3000
		x"dc",	--3001
		x"81",	--3002
		x"04",	--3003
		x"81",	--3004
		x"06",	--3005
		x"81",	--3006
		x"00",	--3007
		x"81",	--3008
		x"02",	--3009
		x"0e",	--3010
		x"3e",	--3011
		x"18",	--3012
		x"0f",	--3013
		x"2f",	--3014
		x"b0",	--3015
		x"2c",	--3016
		x"0e",	--3017
		x"3e",	--3018
		x"10",	--3019
		x"0f",	--3020
		x"b0",	--3021
		x"2c",	--3022
		x"5f",	--3023
		x"18",	--3024
		x"6f",	--3025
		x"b6",	--3026
		x"5e",	--3027
		x"10",	--3028
		x"6e",	--3029
		x"d9",	--3030
		x"6f",	--3031
		x"ae",	--3032
		x"6e",	--3033
		x"e2",	--3034
		x"6f",	--3035
		x"ac",	--3036
		x"6e",	--3037
		x"d1",	--3038
		x"14",	--3039
		x"1c",	--3040
		x"15",	--3041
		x"1e",	--3042
		x"18",	--3043
		x"14",	--3044
		x"19",	--3045
		x"16",	--3046
		x"3c",	--3047
		x"20",	--3048
		x"0e",	--3049
		x"0f",	--3050
		x"06",	--3051
		x"07",	--3052
		x"81",	--3053
		x"20",	--3054
		x"81",	--3055
		x"22",	--3056
		x"0a",	--3057
		x"0b",	--3058
		x"81",	--3059
		x"20",	--3060
		x"08",	--3061
		x"08",	--3062
		x"09",	--3063
		x"12",	--3064
		x"05",	--3065
		x"04",	--3066
		x"b1",	--3067
		x"20",	--3068
		x"19",	--3069
		x"14",	--3070
		x"0d",	--3071
		x"0a",	--3072
		x"0b",	--3073
		x"0e",	--3074
		x"0f",	--3075
		x"1c",	--3076
		x"0d",	--3077
		x"0b",	--3078
		x"03",	--3079
		x"0b",	--3080
		x"0c",	--3081
		x"0d",	--3082
		x"0e",	--3083
		x"0f",	--3084
		x"06",	--3085
		x"07",	--3086
		x"09",	--3087
		x"e5",	--3088
		x"16",	--3089
		x"07",	--3090
		x"e2",	--3091
		x"0a",	--3092
		x"f5",	--3093
		x"f2",	--3094
		x"81",	--3095
		x"20",	--3096
		x"81",	--3097
		x"22",	--3098
		x"0c",	--3099
		x"1a",	--3100
		x"1a",	--3101
		x"1a",	--3102
		x"12",	--3103
		x"06",	--3104
		x"26",	--3105
		x"81",	--3106
		x"0a",	--3107
		x"5d",	--3108
		x"d1",	--3109
		x"11",	--3110
		x"19",	--3111
		x"83",	--3112
		x"c1",	--3113
		x"09",	--3114
		x"0c",	--3115
		x"3c",	--3116
		x"3f",	--3117
		x"00",	--3118
		x"18",	--3119
		x"1d",	--3120
		x"0a",	--3121
		x"3d",	--3122
		x"1a",	--3123
		x"20",	--3124
		x"1b",	--3125
		x"22",	--3126
		x"0c",	--3127
		x"0e",	--3128
		x"0f",	--3129
		x"0b",	--3130
		x"2a",	--3131
		x"0a",	--3132
		x"0b",	--3133
		x"3d",	--3134
		x"3f",	--3135
		x"00",	--3136
		x"f5",	--3137
		x"81",	--3138
		x"20",	--3139
		x"81",	--3140
		x"22",	--3141
		x"81",	--3142
		x"0a",	--3143
		x"0c",	--3144
		x"0d",	--3145
		x"3c",	--3146
		x"7f",	--3147
		x"0d",	--3148
		x"3c",	--3149
		x"40",	--3150
		x"44",	--3151
		x"81",	--3152
		x"0c",	--3153
		x"81",	--3154
		x"0e",	--3155
		x"f1",	--3156
		x"03",	--3157
		x"08",	--3158
		x"0f",	--3159
		x"3f",	--3160
		x"b0",	--3161
		x"4e",	--3162
		x"31",	--3163
		x"24",	--3164
		x"34",	--3165
		x"35",	--3166
		x"36",	--3167
		x"37",	--3168
		x"38",	--3169
		x"39",	--3170
		x"3a",	--3171
		x"3b",	--3172
		x"30",	--3173
		x"1e",	--3174
		x"0f",	--3175
		x"d3",	--3176
		x"3a",	--3177
		x"03",	--3178
		x"08",	--3179
		x"1e",	--3180
		x"10",	--3181
		x"1c",	--3182
		x"20",	--3183
		x"1d",	--3184
		x"22",	--3185
		x"12",	--3186
		x"0d",	--3187
		x"0c",	--3188
		x"06",	--3189
		x"07",	--3190
		x"06",	--3191
		x"37",	--3192
		x"00",	--3193
		x"81",	--3194
		x"20",	--3195
		x"81",	--3196
		x"22",	--3197
		x"12",	--3198
		x"0f",	--3199
		x"0e",	--3200
		x"1a",	--3201
		x"0f",	--3202
		x"e7",	--3203
		x"81",	--3204
		x"0a",	--3205
		x"a6",	--3206
		x"6e",	--3207
		x"36",	--3208
		x"5f",	--3209
		x"d1",	--3210
		x"11",	--3211
		x"19",	--3212
		x"20",	--3213
		x"c1",	--3214
		x"19",	--3215
		x"0f",	--3216
		x"3f",	--3217
		x"18",	--3218
		x"c5",	--3219
		x"0d",	--3220
		x"ba",	--3221
		x"0c",	--3222
		x"0d",	--3223
		x"3c",	--3224
		x"80",	--3225
		x"0d",	--3226
		x"0c",	--3227
		x"b3",	--3228
		x"0d",	--3229
		x"b1",	--3230
		x"81",	--3231
		x"20",	--3232
		x"03",	--3233
		x"81",	--3234
		x"22",	--3235
		x"ab",	--3236
		x"3e",	--3237
		x"40",	--3238
		x"0f",	--3239
		x"3e",	--3240
		x"80",	--3241
		x"3f",	--3242
		x"a4",	--3243
		x"4d",	--3244
		x"7b",	--3245
		x"4f",	--3246
		x"de",	--3247
		x"5f",	--3248
		x"d1",	--3249
		x"11",	--3250
		x"19",	--3251
		x"06",	--3252
		x"c1",	--3253
		x"11",	--3254
		x"0f",	--3255
		x"3f",	--3256
		x"10",	--3257
		x"9e",	--3258
		x"4f",	--3259
		x"f8",	--3260
		x"6f",	--3261
		x"f1",	--3262
		x"3f",	--3263
		x"c2",	--3264
		x"97",	--3265
		x"0b",	--3266
		x"0a",	--3267
		x"09",	--3268
		x"08",	--3269
		x"07",	--3270
		x"31",	--3271
		x"e8",	--3272
		x"81",	--3273
		x"04",	--3274
		x"81",	--3275
		x"06",	--3276
		x"81",	--3277
		x"00",	--3278
		x"81",	--3279
		x"02",	--3280
		x"0e",	--3281
		x"3e",	--3282
		x"10",	--3283
		x"0f",	--3284
		x"2f",	--3285
		x"b0",	--3286
		x"2c",	--3287
		x"0e",	--3288
		x"3e",	--3289
		x"0f",	--3290
		x"b0",	--3291
		x"2c",	--3292
		x"5f",	--3293
		x"10",	--3294
		x"6f",	--3295
		x"5d",	--3296
		x"5e",	--3297
		x"08",	--3298
		x"6e",	--3299
		x"82",	--3300
		x"d1",	--3301
		x"09",	--3302
		x"11",	--3303
		x"6f",	--3304
		x"58",	--3305
		x"6f",	--3306
		x"56",	--3307
		x"6e",	--3308
		x"6f",	--3309
		x"6e",	--3310
		x"4c",	--3311
		x"1d",	--3312
		x"12",	--3313
		x"1d",	--3314
		x"0a",	--3315
		x"81",	--3316
		x"12",	--3317
		x"1e",	--3318
		x"14",	--3319
		x"1f",	--3320
		x"16",	--3321
		x"18",	--3322
		x"0c",	--3323
		x"19",	--3324
		x"0e",	--3325
		x"0f",	--3326
		x"1e",	--3327
		x"0e",	--3328
		x"0f",	--3329
		x"3d",	--3330
		x"81",	--3331
		x"12",	--3332
		x"37",	--3333
		x"1f",	--3334
		x"0c",	--3335
		x"3d",	--3336
		x"00",	--3337
		x"0a",	--3338
		x"0b",	--3339
		x"0b",	--3340
		x"0a",	--3341
		x"0b",	--3342
		x"0e",	--3343
		x"0f",	--3344
		x"12",	--3345
		x"0d",	--3346
		x"0c",	--3347
		x"0e",	--3348
		x"0f",	--3349
		x"37",	--3350
		x"0b",	--3351
		x"0f",	--3352
		x"f7",	--3353
		x"f2",	--3354
		x"0e",	--3355
		x"f4",	--3356
		x"ef",	--3357
		x"09",	--3358
		x"e5",	--3359
		x"0e",	--3360
		x"e3",	--3361
		x"dd",	--3362
		x"0c",	--3363
		x"0d",	--3364
		x"3c",	--3365
		x"7f",	--3366
		x"0d",	--3367
		x"3c",	--3368
		x"40",	--3369
		x"1c",	--3370
		x"81",	--3371
		x"14",	--3372
		x"81",	--3373
		x"16",	--3374
		x"0f",	--3375
		x"3f",	--3376
		x"10",	--3377
		x"b0",	--3378
		x"4e",	--3379
		x"31",	--3380
		x"18",	--3381
		x"37",	--3382
		x"38",	--3383
		x"39",	--3384
		x"3a",	--3385
		x"3b",	--3386
		x"30",	--3387
		x"e1",	--3388
		x"10",	--3389
		x"0f",	--3390
		x"3f",	--3391
		x"10",	--3392
		x"f0",	--3393
		x"4f",	--3394
		x"fa",	--3395
		x"3f",	--3396
		x"c2",	--3397
		x"eb",	--3398
		x"0d",	--3399
		x"e2",	--3400
		x"0c",	--3401
		x"0d",	--3402
		x"3c",	--3403
		x"80",	--3404
		x"0d",	--3405
		x"0c",	--3406
		x"db",	--3407
		x"0d",	--3408
		x"d9",	--3409
		x"0e",	--3410
		x"02",	--3411
		x"0f",	--3412
		x"d5",	--3413
		x"3a",	--3414
		x"40",	--3415
		x"0b",	--3416
		x"3a",	--3417
		x"80",	--3418
		x"3b",	--3419
		x"ce",	--3420
		x"81",	--3421
		x"14",	--3422
		x"81",	--3423
		x"16",	--3424
		x"81",	--3425
		x"12",	--3426
		x"0f",	--3427
		x"3f",	--3428
		x"10",	--3429
		x"cb",	--3430
		x"0f",	--3431
		x"3f",	--3432
		x"c8",	--3433
		x"31",	--3434
		x"e8",	--3435
		x"81",	--3436
		x"04",	--3437
		x"81",	--3438
		x"06",	--3439
		x"81",	--3440
		x"00",	--3441
		x"81",	--3442
		x"02",	--3443
		x"0e",	--3444
		x"3e",	--3445
		x"10",	--3446
		x"0f",	--3447
		x"2f",	--3448
		x"b0",	--3449
		x"2c",	--3450
		x"0e",	--3451
		x"3e",	--3452
		x"0f",	--3453
		x"b0",	--3454
		x"2c",	--3455
		x"e1",	--3456
		x"10",	--3457
		x"0d",	--3458
		x"e1",	--3459
		x"08",	--3460
		x"0a",	--3461
		x"0e",	--3462
		x"3e",	--3463
		x"0f",	--3464
		x"3f",	--3465
		x"10",	--3466
		x"b0",	--3467
		x"50",	--3468
		x"31",	--3469
		x"18",	--3470
		x"30",	--3471
		x"3f",	--3472
		x"fb",	--3473
		x"31",	--3474
		x"e8",	--3475
		x"81",	--3476
		x"04",	--3477
		x"81",	--3478
		x"06",	--3479
		x"81",	--3480
		x"00",	--3481
		x"81",	--3482
		x"02",	--3483
		x"0e",	--3484
		x"3e",	--3485
		x"10",	--3486
		x"0f",	--3487
		x"2f",	--3488
		x"b0",	--3489
		x"2c",	--3490
		x"0e",	--3491
		x"3e",	--3492
		x"0f",	--3493
		x"b0",	--3494
		x"2c",	--3495
		x"e1",	--3496
		x"10",	--3497
		x"0d",	--3498
		x"e1",	--3499
		x"08",	--3500
		x"0a",	--3501
		x"0e",	--3502
		x"3e",	--3503
		x"0f",	--3504
		x"3f",	--3505
		x"10",	--3506
		x"b0",	--3507
		x"50",	--3508
		x"31",	--3509
		x"18",	--3510
		x"30",	--3511
		x"3f",	--3512
		x"fb",	--3513
		x"31",	--3514
		x"e8",	--3515
		x"81",	--3516
		x"04",	--3517
		x"81",	--3518
		x"06",	--3519
		x"81",	--3520
		x"00",	--3521
		x"81",	--3522
		x"02",	--3523
		x"0e",	--3524
		x"3e",	--3525
		x"10",	--3526
		x"0f",	--3527
		x"2f",	--3528
		x"b0",	--3529
		x"2c",	--3530
		x"0e",	--3531
		x"3e",	--3532
		x"0f",	--3533
		x"b0",	--3534
		x"2c",	--3535
		x"e1",	--3536
		x"10",	--3537
		x"0d",	--3538
		x"e1",	--3539
		x"08",	--3540
		x"0a",	--3541
		x"0e",	--3542
		x"3e",	--3543
		x"0f",	--3544
		x"3f",	--3545
		x"10",	--3546
		x"b0",	--3547
		x"50",	--3548
		x"31",	--3549
		x"18",	--3550
		x"30",	--3551
		x"1f",	--3552
		x"fb",	--3553
		x"0b",	--3554
		x"0a",	--3555
		x"31",	--3556
		x"f1",	--3557
		x"03",	--3558
		x"00",	--3559
		x"0d",	--3560
		x"0d",	--3561
		x"0d",	--3562
		x"0d",	--3563
		x"4c",	--3564
		x"c1",	--3565
		x"01",	--3566
		x"0e",	--3567
		x"0b",	--3568
		x"0f",	--3569
		x"09",	--3570
		x"e1",	--3571
		x"00",	--3572
		x"0f",	--3573
		x"b0",	--3574
		x"4e",	--3575
		x"31",	--3576
		x"3a",	--3577
		x"3b",	--3578
		x"30",	--3579
		x"b1",	--3580
		x"1e",	--3581
		x"02",	--3582
		x"4c",	--3583
		x"1b",	--3584
		x"0a",	--3585
		x"0b",	--3586
		x"81",	--3587
		x"04",	--3588
		x"81",	--3589
		x"06",	--3590
		x"0e",	--3591
		x"0f",	--3592
		x"b0",	--3593
		x"dc",	--3594
		x"3f",	--3595
		x"1f",	--3596
		x"e7",	--3597
		x"81",	--3598
		x"04",	--3599
		x"81",	--3600
		x"06",	--3601
		x"4e",	--3602
		x"7e",	--3603
		x"1f",	--3604
		x"0f",	--3605
		x"3e",	--3606
		x"1e",	--3607
		x"0e",	--3608
		x"81",	--3609
		x"02",	--3610
		x"d9",	--3611
		x"0e",	--3612
		x"10",	--3613
		x"0a",	--3614
		x"0b",	--3615
		x"3a",	--3616
		x"3b",	--3617
		x"1a",	--3618
		x"0b",	--3619
		x"de",	--3620
		x"91",	--3621
		x"04",	--3622
		x"04",	--3623
		x"91",	--3624
		x"06",	--3625
		x"06",	--3626
		x"7e",	--3627
		x"f8",	--3628
		x"e8",	--3629
		x"3f",	--3630
		x"00",	--3631
		x"ed",	--3632
		x"0e",	--3633
		x"3f",	--3634
		x"00",	--3635
		x"c3",	--3636
		x"31",	--3637
		x"f4",	--3638
		x"81",	--3639
		x"00",	--3640
		x"81",	--3641
		x"02",	--3642
		x"0e",	--3643
		x"2e",	--3644
		x"0f",	--3645
		x"b0",	--3646
		x"2c",	--3647
		x"5f",	--3648
		x"04",	--3649
		x"6f",	--3650
		x"28",	--3651
		x"27",	--3652
		x"6f",	--3653
		x"07",	--3654
		x"1d",	--3655
		x"06",	--3656
		x"0d",	--3657
		x"21",	--3658
		x"3d",	--3659
		x"1f",	--3660
		x"09",	--3661
		x"c1",	--3662
		x"05",	--3663
		x"26",	--3664
		x"3e",	--3665
		x"3f",	--3666
		x"ff",	--3667
		x"31",	--3668
		x"0c",	--3669
		x"30",	--3670
		x"1e",	--3671
		x"08",	--3672
		x"1f",	--3673
		x"0a",	--3674
		x"3c",	--3675
		x"1e",	--3676
		x"4c",	--3677
		x"4d",	--3678
		x"7d",	--3679
		x"1f",	--3680
		x"0f",	--3681
		x"c1",	--3682
		x"05",	--3683
		x"ef",	--3684
		x"3e",	--3685
		x"3f",	--3686
		x"1e",	--3687
		x"0f",	--3688
		x"31",	--3689
		x"0c",	--3690
		x"30",	--3691
		x"0e",	--3692
		x"0f",	--3693
		x"31",	--3694
		x"0c",	--3695
		x"30",	--3696
		x"12",	--3697
		x"0f",	--3698
		x"0e",	--3699
		x"7d",	--3700
		x"fb",	--3701
		x"eb",	--3702
		x"0e",	--3703
		x"3f",	--3704
		x"00",	--3705
		x"31",	--3706
		x"0c",	--3707
		x"30",	--3708
		x"0b",	--3709
		x"0a",	--3710
		x"09",	--3711
		x"08",	--3712
		x"31",	--3713
		x"0a",	--3714
		x"0b",	--3715
		x"c1",	--3716
		x"01",	--3717
		x"0e",	--3718
		x"0d",	--3719
		x"0b",	--3720
		x"0b",	--3721
		x"e1",	--3722
		x"00",	--3723
		x"0f",	--3724
		x"b0",	--3725
		x"4e",	--3726
		x"31",	--3727
		x"38",	--3728
		x"39",	--3729
		x"3a",	--3730
		x"3b",	--3731
		x"30",	--3732
		x"f1",	--3733
		x"03",	--3734
		x"00",	--3735
		x"b1",	--3736
		x"1e",	--3737
		x"02",	--3738
		x"81",	--3739
		x"04",	--3740
		x"81",	--3741
		x"06",	--3742
		x"0e",	--3743
		x"0f",	--3744
		x"b0",	--3745
		x"dc",	--3746
		x"3f",	--3747
		x"0f",	--3748
		x"18",	--3749
		x"e5",	--3750
		x"81",	--3751
		x"04",	--3752
		x"81",	--3753
		x"06",	--3754
		x"4e",	--3755
		x"7e",	--3756
		x"1f",	--3757
		x"06",	--3758
		x"3e",	--3759
		x"1e",	--3760
		x"0e",	--3761
		x"81",	--3762
		x"02",	--3763
		x"d7",	--3764
		x"91",	--3765
		x"04",	--3766
		x"04",	--3767
		x"91",	--3768
		x"06",	--3769
		x"06",	--3770
		x"7e",	--3771
		x"f8",	--3772
		x"f1",	--3773
		x"0e",	--3774
		x"3e",	--3775
		x"1e",	--3776
		x"1c",	--3777
		x"0d",	--3778
		x"48",	--3779
		x"78",	--3780
		x"1f",	--3781
		x"04",	--3782
		x"0c",	--3783
		x"0d",	--3784
		x"78",	--3785
		x"fc",	--3786
		x"3c",	--3787
		x"3d",	--3788
		x"0c",	--3789
		x"0d",	--3790
		x"18",	--3791
		x"09",	--3792
		x"0c",	--3793
		x"04",	--3794
		x"0d",	--3795
		x"02",	--3796
		x"08",	--3797
		x"09",	--3798
		x"7e",	--3799
		x"1f",	--3800
		x"0e",	--3801
		x"0d",	--3802
		x"0e",	--3803
		x"0d",	--3804
		x"0e",	--3805
		x"81",	--3806
		x"04",	--3807
		x"81",	--3808
		x"06",	--3809
		x"3e",	--3810
		x"1e",	--3811
		x"0e",	--3812
		x"81",	--3813
		x"02",	--3814
		x"a4",	--3815
		x"12",	--3816
		x"0b",	--3817
		x"0a",	--3818
		x"7e",	--3819
		x"fb",	--3820
		x"ec",	--3821
		x"0b",	--3822
		x"0a",	--3823
		x"09",	--3824
		x"1f",	--3825
		x"17",	--3826
		x"3e",	--3827
		x"00",	--3828
		x"2c",	--3829
		x"3a",	--3830
		x"18",	--3831
		x"0b",	--3832
		x"39",	--3833
		x"0c",	--3834
		x"0d",	--3835
		x"4f",	--3836
		x"4f",	--3837
		x"17",	--3838
		x"3c",	--3839
		x"ca",	--3840
		x"6e",	--3841
		x"0f",	--3842
		x"0a",	--3843
		x"0b",	--3844
		x"0f",	--3845
		x"39",	--3846
		x"3a",	--3847
		x"3b",	--3848
		x"30",	--3849
		x"3f",	--3850
		x"00",	--3851
		x"0f",	--3852
		x"3a",	--3853
		x"0b",	--3854
		x"39",	--3855
		x"18",	--3856
		x"0c",	--3857
		x"0d",	--3858
		x"4f",	--3859
		x"4f",	--3860
		x"e9",	--3861
		x"12",	--3862
		x"0d",	--3863
		x"0c",	--3864
		x"7f",	--3865
		x"fb",	--3866
		x"e3",	--3867
		x"3a",	--3868
		x"10",	--3869
		x"0b",	--3870
		x"39",	--3871
		x"10",	--3872
		x"ef",	--3873
		x"3a",	--3874
		x"20",	--3875
		x"0b",	--3876
		x"09",	--3877
		x"ea",	--3878
		x"0b",	--3879
		x"0a",	--3880
		x"09",	--3881
		x"08",	--3882
		x"07",	--3883
		x"0d",	--3884
		x"1e",	--3885
		x"04",	--3886
		x"1f",	--3887
		x"06",	--3888
		x"5a",	--3889
		x"01",	--3890
		x"6c",	--3891
		x"6c",	--3892
		x"70",	--3893
		x"6c",	--3894
		x"6a",	--3895
		x"6c",	--3896
		x"36",	--3897
		x"0e",	--3898
		x"32",	--3899
		x"1b",	--3900
		x"02",	--3901
		x"3b",	--3902
		x"82",	--3903
		x"6d",	--3904
		x"3b",	--3905
		x"80",	--3906
		x"5e",	--3907
		x"0c",	--3908
		x"0d",	--3909
		x"3c",	--3910
		x"7f",	--3911
		x"0d",	--3912
		x"3c",	--3913
		x"40",	--3914
		x"40",	--3915
		x"3e",	--3916
		x"3f",	--3917
		x"0f",	--3918
		x"0f",	--3919
		x"4a",	--3920
		x"0d",	--3921
		x"3d",	--3922
		x"7f",	--3923
		x"12",	--3924
		x"0f",	--3925
		x"0e",	--3926
		x"12",	--3927
		x"0f",	--3928
		x"0e",	--3929
		x"12",	--3930
		x"0f",	--3931
		x"0e",	--3932
		x"12",	--3933
		x"0f",	--3934
		x"0e",	--3935
		x"12",	--3936
		x"0f",	--3937
		x"0e",	--3938
		x"12",	--3939
		x"0f",	--3940
		x"0e",	--3941
		x"12",	--3942
		x"0f",	--3943
		x"0e",	--3944
		x"3e",	--3945
		x"3f",	--3946
		x"7f",	--3947
		x"4d",	--3948
		x"05",	--3949
		x"0f",	--3950
		x"cc",	--3951
		x"4d",	--3952
		x"0e",	--3953
		x"0f",	--3954
		x"4d",	--3955
		x"0d",	--3956
		x"0d",	--3957
		x"0d",	--3958
		x"0d",	--3959
		x"0d",	--3960
		x"0d",	--3961
		x"0d",	--3962
		x"0c",	--3963
		x"3c",	--3964
		x"7f",	--3965
		x"0c",	--3966
		x"4f",	--3967
		x"0f",	--3968
		x"0f",	--3969
		x"0f",	--3970
		x"0d",	--3971
		x"0d",	--3972
		x"0f",	--3973
		x"37",	--3974
		x"38",	--3975
		x"39",	--3976
		x"3a",	--3977
		x"3b",	--3978
		x"30",	--3979
		x"0d",	--3980
		x"be",	--3981
		x"0c",	--3982
		x"0d",	--3983
		x"3c",	--3984
		x"80",	--3985
		x"0d",	--3986
		x"0c",	--3987
		x"02",	--3988
		x"0d",	--3989
		x"b8",	--3990
		x"3e",	--3991
		x"40",	--3992
		x"0f",	--3993
		x"b4",	--3994
		x"12",	--3995
		x"0f",	--3996
		x"0e",	--3997
		x"0d",	--3998
		x"3d",	--3999
		x"80",	--4000
		x"b2",	--4001
		x"7d",	--4002
		x"0e",	--4003
		x"0f",	--4004
		x"cd",	--4005
		x"0e",	--4006
		x"3f",	--4007
		x"10",	--4008
		x"3e",	--4009
		x"3f",	--4010
		x"7f",	--4011
		x"7d",	--4012
		x"c5",	--4013
		x"37",	--4014
		x"82",	--4015
		x"07",	--4016
		x"37",	--4017
		x"1a",	--4018
		x"4f",	--4019
		x"0c",	--4020
		x"0d",	--4021
		x"4b",	--4022
		x"7b",	--4023
		x"1f",	--4024
		x"05",	--4025
		x"12",	--4026
		x"0d",	--4027
		x"0c",	--4028
		x"7b",	--4029
		x"fb",	--4030
		x"18",	--4031
		x"09",	--4032
		x"77",	--4033
		x"1f",	--4034
		x"04",	--4035
		x"08",	--4036
		x"09",	--4037
		x"77",	--4038
		x"fc",	--4039
		x"38",	--4040
		x"39",	--4041
		x"08",	--4042
		x"09",	--4043
		x"1e",	--4044
		x"0f",	--4045
		x"08",	--4046
		x"04",	--4047
		x"09",	--4048
		x"02",	--4049
		x"0e",	--4050
		x"0f",	--4051
		x"08",	--4052
		x"09",	--4053
		x"08",	--4054
		x"09",	--4055
		x"0e",	--4056
		x"0f",	--4057
		x"3e",	--4058
		x"7f",	--4059
		x"0f",	--4060
		x"3e",	--4061
		x"40",	--4062
		x"26",	--4063
		x"38",	--4064
		x"3f",	--4065
		x"09",	--4066
		x"0e",	--4067
		x"0f",	--4068
		x"12",	--4069
		x"0f",	--4070
		x"0e",	--4071
		x"12",	--4072
		x"0f",	--4073
		x"0e",	--4074
		x"12",	--4075
		x"0f",	--4076
		x"0e",	--4077
		x"12",	--4078
		x"0f",	--4079
		x"0e",	--4080
		x"12",	--4081
		x"0f",	--4082
		x"0e",	--4083
		x"12",	--4084
		x"0f",	--4085
		x"0e",	--4086
		x"12",	--4087
		x"0f",	--4088
		x"0e",	--4089
		x"3e",	--4090
		x"3f",	--4091
		x"7f",	--4092
		x"5d",	--4093
		x"39",	--4094
		x"00",	--4095
		x"72",	--4096
		x"4d",	--4097
		x"70",	--4098
		x"08",	--4099
		x"09",	--4100
		x"da",	--4101
		x"0f",	--4102
		x"d8",	--4103
		x"0e",	--4104
		x"0f",	--4105
		x"3e",	--4106
		x"80",	--4107
		x"0f",	--4108
		x"0e",	--4109
		x"04",	--4110
		x"38",	--4111
		x"40",	--4112
		x"09",	--4113
		x"d0",	--4114
		x"0f",	--4115
		x"ce",	--4116
		x"f9",	--4117
		x"0b",	--4118
		x"0a",	--4119
		x"2a",	--4120
		x"5b",	--4121
		x"02",	--4122
		x"3b",	--4123
		x"7f",	--4124
		x"1d",	--4125
		x"02",	--4126
		x"12",	--4127
		x"0d",	--4128
		x"12",	--4129
		x"0d",	--4130
		x"12",	--4131
		x"0d",	--4132
		x"12",	--4133
		x"0d",	--4134
		x"12",	--4135
		x"0d",	--4136
		x"12",	--4137
		x"0d",	--4138
		x"12",	--4139
		x"0d",	--4140
		x"4d",	--4141
		x"5f",	--4142
		x"03",	--4143
		x"3f",	--4144
		x"80",	--4145
		x"0f",	--4146
		x"0f",	--4147
		x"ce",	--4148
		x"01",	--4149
		x"0d",	--4150
		x"2d",	--4151
		x"0a",	--4152
		x"51",	--4153
		x"be",	--4154
		x"82",	--4155
		x"02",	--4156
		x"0c",	--4157
		x"0d",	--4158
		x"0c",	--4159
		x"0d",	--4160
		x"0c",	--4161
		x"0d",	--4162
		x"0c",	--4163
		x"0d",	--4164
		x"0c",	--4165
		x"0d",	--4166
		x"0c",	--4167
		x"0d",	--4168
		x"0c",	--4169
		x"0d",	--4170
		x"0c",	--4171
		x"0d",	--4172
		x"fe",	--4173
		x"03",	--4174
		x"00",	--4175
		x"3d",	--4176
		x"00",	--4177
		x"0b",	--4178
		x"3f",	--4179
		x"81",	--4180
		x"0c",	--4181
		x"0d",	--4182
		x"0a",	--4183
		x"3f",	--4184
		x"3d",	--4185
		x"00",	--4186
		x"f9",	--4187
		x"8e",	--4188
		x"02",	--4189
		x"8e",	--4190
		x"04",	--4191
		x"8e",	--4192
		x"06",	--4193
		x"3a",	--4194
		x"3b",	--4195
		x"30",	--4196
		x"3d",	--4197
		x"ff",	--4198
		x"2a",	--4199
		x"3d",	--4200
		x"81",	--4201
		x"8e",	--4202
		x"02",	--4203
		x"fe",	--4204
		x"03",	--4205
		x"00",	--4206
		x"0c",	--4207
		x"0d",	--4208
		x"0c",	--4209
		x"0d",	--4210
		x"0c",	--4211
		x"0d",	--4212
		x"0c",	--4213
		x"0d",	--4214
		x"0c",	--4215
		x"0d",	--4216
		x"0c",	--4217
		x"0d",	--4218
		x"0c",	--4219
		x"0d",	--4220
		x"0c",	--4221
		x"0d",	--4222
		x"0a",	--4223
		x"0b",	--4224
		x"0a",	--4225
		x"3b",	--4226
		x"00",	--4227
		x"8e",	--4228
		x"04",	--4229
		x"8e",	--4230
		x"06",	--4231
		x"3a",	--4232
		x"3b",	--4233
		x"30",	--4234
		x"0b",	--4235
		x"ad",	--4236
		x"ee",	--4237
		x"00",	--4238
		x"3a",	--4239
		x"3b",	--4240
		x"30",	--4241
		x"0a",	--4242
		x"0c",	--4243
		x"0c",	--4244
		x"0d",	--4245
		x"0c",	--4246
		x"3d",	--4247
		x"10",	--4248
		x"0c",	--4249
		x"02",	--4250
		x"0d",	--4251
		x"08",	--4252
		x"de",	--4253
		x"00",	--4254
		x"e4",	--4255
		x"0b",	--4256
		x"f2",	--4257
		x"ee",	--4258
		x"00",	--4259
		x"e3",	--4260
		x"ce",	--4261
		x"00",	--4262
		x"dc",	--4263
		x"0b",	--4264
		x"6d",	--4265
		x"6d",	--4266
		x"12",	--4267
		x"6c",	--4268
		x"6c",	--4269
		x"0f",	--4270
		x"6d",	--4271
		x"41",	--4272
		x"6c",	--4273
		x"11",	--4274
		x"6d",	--4275
		x"0d",	--4276
		x"6c",	--4277
		x"14",	--4278
		x"5d",	--4279
		x"01",	--4280
		x"5d",	--4281
		x"01",	--4282
		x"14",	--4283
		x"4d",	--4284
		x"09",	--4285
		x"1e",	--4286
		x"0f",	--4287
		x"3b",	--4288
		x"30",	--4289
		x"6c",	--4290
		x"28",	--4291
		x"ce",	--4292
		x"01",	--4293
		x"f7",	--4294
		x"3e",	--4295
		x"0f",	--4296
		x"3b",	--4297
		x"30",	--4298
		x"cf",	--4299
		x"01",	--4300
		x"f0",	--4301
		x"3e",	--4302
		x"f8",	--4303
		x"1b",	--4304
		x"02",	--4305
		x"1c",	--4306
		x"02",	--4307
		x"0c",	--4308
		x"e6",	--4309
		x"0b",	--4310
		x"16",	--4311
		x"1b",	--4312
		x"04",	--4313
		x"1f",	--4314
		x"06",	--4315
		x"1c",	--4316
		x"04",	--4317
		x"1e",	--4318
		x"06",	--4319
		x"0e",	--4320
		x"da",	--4321
		x"0f",	--4322
		x"02",	--4323
		x"0c",	--4324
		x"d6",	--4325
		x"0f",	--4326
		x"06",	--4327
		x"0e",	--4328
		x"02",	--4329
		x"0b",	--4330
		x"02",	--4331
		x"0e",	--4332
		x"d1",	--4333
		x"4d",	--4334
		x"ce",	--4335
		x"3e",	--4336
		x"d6",	--4337
		x"6c",	--4338
		x"d7",	--4339
		x"5e",	--4340
		x"01",	--4341
		x"5f",	--4342
		x"01",	--4343
		x"0e",	--4344
		x"c5",	--4345
		x"1e",	--4346
		x"1e",	--4347
		x"1e",	--4348
		x"0b",	--4349
		x"1d",	--4350
		x"1c",	--4351
		x"cd",	--4352
		x"00",	--4353
		x"1d",	--4354
		x"82",	--4355
		x"1c",	--4356
		x"3e",	--4357
		x"82",	--4358
		x"1e",	--4359
		x"30",	--4360
		x"3f",	--4361
		x"30",	--4362
		x"0b",	--4363
		x"0a",	--4364
		x"21",	--4365
		x"81",	--4366
		x"00",	--4367
		x"1a",	--4368
		x"1c",	--4369
		x"1b",	--4370
		x"1e",	--4371
		x"0d",	--4372
		x"0e",	--4373
		x"3f",	--4374
		x"f4",	--4375
		x"b0",	--4376
		x"48",	--4377
		x"0f",	--4378
		x"05",	--4379
		x"0e",	--4380
		x"0e",	--4381
		x"ce",	--4382
		x"ff",	--4383
		x"04",	--4384
		x"1e",	--4385
		x"1c",	--4386
		x"ce",	--4387
		x"00",	--4388
		x"21",	--4389
		x"3a",	--4390
		x"3b",	--4391
		x"30",	--4392
		x"92",	--4393
		x"02",	--4394
		x"1c",	--4395
		x"b2",	--4396
		x"ff",	--4397
		x"1e",	--4398
		x"0e",	--4399
		x"3e",	--4400
		x"06",	--4401
		x"1f",	--4402
		x"04",	--4403
		x"b0",	--4404
		x"16",	--4405
		x"30",	--4406
		x"92",	--4407
		x"02",	--4408
		x"1c",	--4409
		x"92",	--4410
		x"04",	--4411
		x"1e",	--4412
		x"0e",	--4413
		x"3e",	--4414
		x"1f",	--4415
		x"06",	--4416
		x"b0",	--4417
		x"16",	--4418
		x"30",	--4419
		x"0c",	--4420
		x"82",	--4421
		x"1c",	--4422
		x"b2",	--4423
		x"ff",	--4424
		x"1e",	--4425
		x"0e",	--4426
		x"0f",	--4427
		x"b0",	--4428
		x"16",	--4429
		x"30",	--4430
		x"82",	--4431
		x"1c",	--4432
		x"82",	--4433
		x"1e",	--4434
		x"0e",	--4435
		x"0f",	--4436
		x"b0",	--4437
		x"16",	--4438
		x"30",	--4439
		x"0b",	--4440
		x"0a",	--4441
		x"09",	--4442
		x"08",	--4443
		x"07",	--4444
		x"06",	--4445
		x"05",	--4446
		x"04",	--4447
		x"31",	--4448
		x"08",	--4449
		x"81",	--4450
		x"04",	--4451
		x"09",	--4452
		x"1f",	--4453
		x"1a",	--4454
		x"1d",	--4455
		x"1c",	--4456
		x"4c",	--4457
		x"04",	--4458
		x"84",	--4459
		x"45",	--4460
		x"4e",	--4461
		x"7e",	--4462
		x"40",	--4463
		x"11",	--4464
		x"f1",	--4465
		x"30",	--4466
		x"00",	--4467
		x"0e",	--4468
		x"8e",	--4469
		x"5e",	--4470
		x"03",	--4471
		x"7e",	--4472
		x"58",	--4473
		x"02",	--4474
		x"7e",	--4475
		x"78",	--4476
		x"c1",	--4477
		x"01",	--4478
		x"0c",	--4479
		x"2c",	--4480
		x"0f",	--4481
		x"7e",	--4482
		x"20",	--4483
		x"04",	--4484
		x"f1",	--4485
		x"30",	--4486
		x"00",	--4487
		x"04",	--4488
		x"4c",	--4489
		x"05",	--4490
		x"c1",	--4491
		x"00",	--4492
		x"0c",	--4493
		x"1c",	--4494
		x"01",	--4495
		x"0c",	--4496
		x"0a",	--4497
		x"8c",	--4498
		x"8c",	--4499
		x"8c",	--4500
		x"8c",	--4501
		x"0b",	--4502
		x"06",	--4503
		x"0c",	--4504
		x"8c",	--4505
		x"8c",	--4506
		x"8c",	--4507
		x"8c",	--4508
		x"07",	--4509
		x"0a",	--4510
		x"0b",	--4511
		x"0e",	--4512
		x"8e",	--4513
		x"c1",	--4514
		x"02",	--4515
		x"6e",	--4516
		x"02",	--4517
		x"07",	--4518
		x"01",	--4519
		x"37",	--4520
		x"4f",	--4521
		x"7f",	--4522
		x"10",	--4523
		x"3c",	--4524
		x"1d",	--4525
		x"04",	--4526
		x"3d",	--4527
		x"1d",	--4528
		x"cd",	--4529
		x"00",	--4530
		x"fc",	--4531
		x"1d",	--4532
		x"04",	--4533
		x"09",	--4534
		x"02",	--4535
		x"09",	--4536
		x"01",	--4537
		x"09",	--4538
		x"e1",	--4539
		x"02",	--4540
		x"05",	--4541
		x"09",	--4542
		x"02",	--4543
		x"09",	--4544
		x"01",	--4545
		x"09",	--4546
		x"05",	--4547
		x"07",	--4548
		x"01",	--4549
		x"05",	--4550
		x"4f",	--4551
		x"0d",	--4552
		x"f1",	--4553
		x"20",	--4554
		x"06",	--4555
		x"06",	--4556
		x"0b",	--4557
		x"0e",	--4558
		x"0f",	--4559
		x"0f",	--4560
		x"6f",	--4561
		x"8f",	--4562
		x"16",	--4563
		x"88",	--4564
		x"01",	--4565
		x"06",	--4566
		x"06",	--4567
		x"f6",	--4568
		x"0b",	--4569
		x"f1",	--4570
		x"30",	--4571
		x"06",	--4572
		x"05",	--4573
		x"05",	--4574
		x"5f",	--4575
		x"06",	--4576
		x"8f",	--4577
		x"88",	--4578
		x"1b",	--4579
		x"0f",	--4580
		x"0f",	--4581
		x"0f",	--4582
		x"f7",	--4583
		x"0a",	--4584
		x"06",	--4585
		x"0b",	--4586
		x"07",	--4587
		x"1b",	--4588
		x"0f",	--4589
		x"0f",	--4590
		x"6f",	--4591
		x"8f",	--4592
		x"16",	--4593
		x"88",	--4594
		x"06",	--4595
		x"f7",	--4596
		x"e1",	--4597
		x"02",	--4598
		x"02",	--4599
		x"4a",	--4600
		x"08",	--4601
		x"1a",	--4602
		x"04",	--4603
		x"0a",	--4604
		x"0d",	--4605
		x"3f",	--4606
		x"30",	--4607
		x"88",	--4608
		x"7a",	--4609
		x"4a",	--4610
		x"fa",	--4611
		x"44",	--4612
		x"0b",	--4613
		x"f3",	--4614
		x"37",	--4615
		x"8f",	--4616
		x"88",	--4617
		x"1b",	--4618
		x"0f",	--4619
		x"0f",	--4620
		x"6f",	--4621
		x"4f",	--4622
		x"07",	--4623
		x"07",	--4624
		x"f5",	--4625
		x"04",	--4626
		x"3f",	--4627
		x"20",	--4628
		x"88",	--4629
		x"1b",	--4630
		x"0b",	--4631
		x"fa",	--4632
		x"0f",	--4633
		x"31",	--4634
		x"34",	--4635
		x"35",	--4636
		x"36",	--4637
		x"37",	--4638
		x"38",	--4639
		x"39",	--4640
		x"3a",	--4641
		x"3b",	--4642
		x"30",	--4643
		x"0b",	--4644
		x"0a",	--4645
		x"09",	--4646
		x"08",	--4647
		x"07",	--4648
		x"06",	--4649
		x"05",	--4650
		x"04",	--4651
		x"31",	--4652
		x"b6",	--4653
		x"81",	--4654
		x"3a",	--4655
		x"06",	--4656
		x"05",	--4657
		x"81",	--4658
		x"3e",	--4659
		x"c1",	--4660
		x"2f",	--4661
		x"c1",	--4662
		x"2b",	--4663
		x"c1",	--4664
		x"2e",	--4665
		x"c1",	--4666
		x"2a",	--4667
		x"81",	--4668
		x"30",	--4669
		x"81",	--4670
		x"26",	--4671
		x"07",	--4672
		x"81",	--4673
		x"2c",	--4674
		x"0e",	--4675
		x"3e",	--4676
		x"1c",	--4677
		x"81",	--4678
		x"1c",	--4679
		x"30",	--4680
		x"c2",	--4681
		x"0f",	--4682
		x"1f",	--4683
		x"81",	--4684
		x"40",	--4685
		x"07",	--4686
		x"1e",	--4687
		x"7e",	--4688
		x"25",	--4689
		x"13",	--4690
		x"81",	--4691
		x"00",	--4692
		x"81",	--4693
		x"02",	--4694
		x"81",	--4695
		x"3e",	--4696
		x"c1",	--4697
		x"2f",	--4698
		x"c1",	--4699
		x"2b",	--4700
		x"c1",	--4701
		x"2e",	--4702
		x"c1",	--4703
		x"2a",	--4704
		x"81",	--4705
		x"30",	--4706
		x"30",	--4707
		x"b8",	--4708
		x"05",	--4709
		x"8e",	--4710
		x"0f",	--4711
		x"91",	--4712
		x"3c",	--4713
		x"91",	--4714
		x"2c",	--4715
		x"30",	--4716
		x"9e",	--4717
		x"7e",	--4718
		x"63",	--4719
		x"c5",	--4720
		x"7e",	--4721
		x"64",	--4722
		x"27",	--4723
		x"7e",	--4724
		x"30",	--4725
		x"94",	--4726
		x"7e",	--4727
		x"31",	--4728
		x"1a",	--4729
		x"7e",	--4730
		x"2a",	--4731
		x"77",	--4732
		x"7e",	--4733
		x"2b",	--4734
		x"0a",	--4735
		x"7e",	--4736
		x"23",	--4737
		x"42",	--4738
		x"7e",	--4739
		x"25",	--4740
		x"e0",	--4741
		x"7e",	--4742
		x"20",	--4743
		x"32",	--4744
		x"56",	--4745
		x"7e",	--4746
		x"2d",	--4747
		x"49",	--4748
		x"7e",	--4749
		x"2e",	--4750
		x"5b",	--4751
		x"7e",	--4752
		x"2b",	--4753
		x"28",	--4754
		x"47",	--4755
		x"7e",	--4756
		x"3a",	--4757
		x"8c",	--4758
		x"7e",	--4759
		x"58",	--4760
		x"21",	--4761
		x"e9",	--4762
		x"7e",	--4763
		x"6f",	--4764
		x"24",	--4765
		x"7e",	--4766
		x"70",	--4767
		x"0a",	--4768
		x"7e",	--4769
		x"69",	--4770
		x"e3",	--4771
		x"7e",	--4772
		x"6c",	--4773
		x"22",	--4774
		x"7e",	--4775
		x"64",	--4776
		x"11",	--4777
		x"dc",	--4778
		x"7e",	--4779
		x"73",	--4780
		x"98",	--4781
		x"7e",	--4782
		x"74",	--4783
		x"04",	--4784
		x"7e",	--4785
		x"70",	--4786
		x"07",	--4787
		x"b8",	--4788
		x"7e",	--4789
		x"75",	--4790
		x"d1",	--4791
		x"7e",	--4792
		x"78",	--4793
		x"d2",	--4794
		x"19",	--4795
		x"3e",	--4796
		x"18",	--4797
		x"2c",	--4798
		x"08",	--4799
		x"30",	--4800
		x"8c",	--4801
		x"b1",	--4802
		x"28",	--4803
		x"cb",	--4804
		x"f1",	--4805
		x"00",	--4806
		x"30",	--4807
		x"bc",	--4808
		x"69",	--4809
		x"59",	--4810
		x"6e",	--4811
		x"04",	--4812
		x"7e",	--4813
		x"fe",	--4814
		x"6e",	--4815
		x"01",	--4816
		x"5e",	--4817
		x"c1",	--4818
		x"00",	--4819
		x"30",	--4820
		x"bc",	--4821
		x"f1",	--4822
		x"10",	--4823
		x"00",	--4824
		x"30",	--4825
		x"bc",	--4826
		x"f1",	--4827
		x"2b",	--4828
		x"02",	--4829
		x"30",	--4830
		x"bc",	--4831
		x"f1",	--4832
		x"2b",	--4833
		x"02",	--4834
		x"02",	--4835
		x"30",	--4836
		x"bc",	--4837
		x"f1",	--4838
		x"20",	--4839
		x"02",	--4840
		x"30",	--4841
		x"bc",	--4842
		x"c1",	--4843
		x"2a",	--4844
		x"02",	--4845
		x"30",	--4846
		x"a2",	--4847
		x"d1",	--4848
		x"2e",	--4849
		x"30",	--4850
		x"bc",	--4851
		x"0e",	--4852
		x"2e",	--4853
		x"2a",	--4854
		x"0a",	--4855
		x"03",	--4856
		x"81",	--4857
		x"26",	--4858
		x"0d",	--4859
		x"c1",	--4860
		x"2e",	--4861
		x"02",	--4862
		x"30",	--4863
		x"b2",	--4864
		x"f1",	--4865
		x"10",	--4866
		x"00",	--4867
		x"3a",	--4868
		x"81",	--4869
		x"26",	--4870
		x"91",	--4871
		x"26",	--4872
		x"05",	--4873
		x"27",	--4874
		x"81",	--4875
		x"26",	--4876
		x"15",	--4877
		x"c1",	--4878
		x"2e",	--4879
		x"12",	--4880
		x"69",	--4881
		x"79",	--4882
		x"10",	--4883
		x"5e",	--4884
		x"01",	--4885
		x"4e",	--4886
		x"4e",	--4887
		x"0e",	--4888
		x"0e",	--4889
		x"4e",	--4890
		x"6a",	--4891
		x"7a",	--4892
		x"7f",	--4893
		x"4a",	--4894
		x"c1",	--4895
		x"00",	--4896
		x"30",	--4897
		x"bc",	--4898
		x"1a",	--4899
		x"26",	--4900
		x"0a",	--4901
		x"0c",	--4902
		x"0c",	--4903
		x"0c",	--4904
		x"0a",	--4905
		x"81",	--4906
		x"26",	--4907
		x"b1",	--4908
		x"d0",	--4909
		x"26",	--4910
		x"8e",	--4911
		x"81",	--4912
		x"26",	--4913
		x"d1",	--4914
		x"2a",	--4915
		x"30",	--4916
		x"bc",	--4917
		x"07",	--4918
		x"27",	--4919
		x"6e",	--4920
		x"c1",	--4921
		x"2e",	--4922
		x"03",	--4923
		x"c1",	--4924
		x"2a",	--4925
		x"26",	--4926
		x"c1",	--4927
		x"04",	--4928
		x"c1",	--4929
		x"05",	--4930
		x"0e",	--4931
		x"2e",	--4932
		x"03",	--4933
		x"07",	--4934
		x"27",	--4935
		x"2e",	--4936
		x"c1",	--4937
		x"2e",	--4938
		x"07",	--4939
		x"e1",	--4940
		x"01",	--4941
		x"1f",	--4942
		x"26",	--4943
		x"c1",	--4944
		x"03",	--4945
		x"06",	--4946
		x"c1",	--4947
		x"2a",	--4948
		x"03",	--4949
		x"91",	--4950
		x"26",	--4951
		x"30",	--4952
		x"0e",	--4953
		x"02",	--4954
		x"3e",	--4955
		x"ca",	--4956
		x"11",	--4957
		x"04",	--4958
		x"11",	--4959
		x"04",	--4960
		x"1d",	--4961
		x"34",	--4962
		x"1f",	--4963
		x"3e",	--4964
		x"b0",	--4965
		x"b0",	--4966
		x"21",	--4967
		x"81",	--4968
		x"2c",	--4969
		x"05",	--4970
		x"30",	--4971
		x"9e",	--4972
		x"07",	--4973
		x"27",	--4974
		x"29",	--4975
		x"81",	--4976
		x"1e",	--4977
		x"5e",	--4978
		x"09",	--4979
		x"01",	--4980
		x"4e",	--4981
		x"4e",	--4982
		x"4e",	--4983
		x"4e",	--4984
		x"6a",	--4985
		x"7a",	--4986
		x"f7",	--4987
		x"4a",	--4988
		x"c1",	--4989
		x"00",	--4990
		x"05",	--4991
		x"b1",	--4992
		x"10",	--4993
		x"28",	--4994
		x"53",	--4995
		x"d1",	--4996
		x"01",	--4997
		x"06",	--4998
		x"e1",	--4999
		x"00",	--5000
		x"b1",	--5001
		x"0a",	--5002
		x"28",	--5003
		x"03",	--5004
		x"b1",	--5005
		x"10",	--5006
		x"28",	--5007
		x"6b",	--5008
		x"6b",	--5009
		x"24",	--5010
		x"0c",	--5011
		x"3c",	--5012
		x"28",	--5013
		x"17",	--5014
		x"02",	--5015
		x"16",	--5016
		x"04",	--5017
		x"1b",	--5018
		x"06",	--5019
		x"81",	--5020
		x"1e",	--5021
		x"81",	--5022
		x"20",	--5023
		x"81",	--5024
		x"22",	--5025
		x"81",	--5026
		x"24",	--5027
		x"d1",	--5028
		x"2b",	--5029
		x"08",	--5030
		x"06",	--5031
		x"07",	--5032
		x"04",	--5033
		x"06",	--5034
		x"02",	--5035
		x"0b",	--5036
		x"02",	--5037
		x"c1",	--5038
		x"2b",	--5039
		x"0b",	--5040
		x"0b",	--5041
		x"0b",	--5042
		x"c1",	--5043
		x"2f",	--5044
		x"05",	--5045
		x"20",	--5046
		x"5b",	--5047
		x"07",	--5048
		x"0d",	--5049
		x"27",	--5050
		x"28",	--5051
		x"1b",	--5052
		x"02",	--5053
		x"81",	--5054
		x"1e",	--5055
		x"81",	--5056
		x"20",	--5057
		x"d1",	--5058
		x"2b",	--5059
		x"08",	--5060
		x"09",	--5061
		x"06",	--5062
		x"27",	--5063
		x"2b",	--5064
		x"81",	--5065
		x"1e",	--5066
		x"d1",	--5067
		x"2b",	--5068
		x"0b",	--5069
		x"02",	--5070
		x"c1",	--5071
		x"2b",	--5072
		x"0b",	--5073
		x"0b",	--5074
		x"0b",	--5075
		x"c1",	--5076
		x"2f",	--5077
		x"05",	--5078
		x"f1",	--5079
		x"00",	--5080
		x"12",	--5081
		x"c1",	--5082
		x"2b",	--5083
		x"0f",	--5084
		x"68",	--5085
		x"b1",	--5086
		x"10",	--5087
		x"28",	--5088
		x"03",	--5089
		x"78",	--5090
		x"40",	--5091
		x"05",	--5092
		x"b1",	--5093
		x"28",	--5094
		x"04",	--5095
		x"78",	--5096
		x"20",	--5097
		x"c1",	--5098
		x"00",	--5099
		x"68",	--5100
		x"68",	--5101
		x"30",	--5102
		x"c1",	--5103
		x"2f",	--5104
		x"2d",	--5105
		x"f1",	--5106
		x"2d",	--5107
		x"02",	--5108
		x"68",	--5109
		x"11",	--5110
		x"b1",	--5111
		x"1e",	--5112
		x"b1",	--5113
		x"20",	--5114
		x"b1",	--5115
		x"22",	--5116
		x"b1",	--5117
		x"24",	--5118
		x"91",	--5119
		x"1e",	--5120
		x"81",	--5121
		x"20",	--5122
		x"81",	--5123
		x"22",	--5124
		x"81",	--5125
		x"24",	--5126
		x"17",	--5127
		x"58",	--5128
		x"0f",	--5129
		x"1a",	--5130
		x"1e",	--5131
		x"1b",	--5132
		x"20",	--5133
		x"3a",	--5134
		x"3b",	--5135
		x"0e",	--5136
		x"0f",	--5137
		x"1e",	--5138
		x"0f",	--5139
		x"81",	--5140
		x"1e",	--5141
		x"81",	--5142
		x"20",	--5143
		x"06",	--5144
		x"1a",	--5145
		x"1e",	--5146
		x"3a",	--5147
		x"1a",	--5148
		x"81",	--5149
		x"1e",	--5150
		x"c1",	--5151
		x"1b",	--5152
		x"68",	--5153
		x"6a",	--5154
		x"16",	--5155
		x"1e",	--5156
		x"91",	--5157
		x"20",	--5158
		x"3c",	--5159
		x"18",	--5160
		x"22",	--5161
		x"14",	--5162
		x"24",	--5163
		x"07",	--5164
		x"37",	--5165
		x"1a",	--5166
		x"09",	--5167
		x"91",	--5168
		x"28",	--5169
		x"32",	--5170
		x"1b",	--5171
		x"28",	--5172
		x"8b",	--5173
		x"8b",	--5174
		x"8b",	--5175
		x"8b",	--5176
		x"81",	--5177
		x"34",	--5178
		x"81",	--5179
		x"36",	--5180
		x"81",	--5181
		x"38",	--5182
		x"11",	--5183
		x"3a",	--5184
		x"11",	--5185
		x"3a",	--5186
		x"11",	--5187
		x"3a",	--5188
		x"11",	--5189
		x"3a",	--5190
		x"0c",	--5191
		x"1d",	--5192
		x"44",	--5193
		x"0e",	--5194
		x"0f",	--5195
		x"b0",	--5196
		x"52",	--5197
		x"31",	--5198
		x"0b",	--5199
		x"3c",	--5200
		x"0a",	--5201
		x"05",	--5202
		x"7b",	--5203
		x"30",	--5204
		x"c7",	--5205
		x"00",	--5206
		x"0c",	--5207
		x"4b",	--5208
		x"d1",	--5209
		x"01",	--5210
		x"03",	--5211
		x"7a",	--5212
		x"37",	--5213
		x"02",	--5214
		x"7a",	--5215
		x"57",	--5216
		x"4a",	--5217
		x"c7",	--5218
		x"00",	--5219
		x"06",	--5220
		x"36",	--5221
		x"11",	--5222
		x"3a",	--5223
		x"11",	--5224
		x"3a",	--5225
		x"11",	--5226
		x"3a",	--5227
		x"11",	--5228
		x"3a",	--5229
		x"0c",	--5230
		x"1d",	--5231
		x"44",	--5232
		x"0e",	--5233
		x"0f",	--5234
		x"b0",	--5235
		x"2c",	--5236
		x"31",	--5237
		x"09",	--5238
		x"81",	--5239
		x"3c",	--5240
		x"08",	--5241
		x"04",	--5242
		x"37",	--5243
		x"0c",	--5244
		x"b2",	--5245
		x"0d",	--5246
		x"b0",	--5247
		x"0e",	--5248
		x"ae",	--5249
		x"0f",	--5250
		x"ac",	--5251
		x"81",	--5252
		x"1e",	--5253
		x"81",	--5254
		x"20",	--5255
		x"81",	--5256
		x"22",	--5257
		x"81",	--5258
		x"24",	--5259
		x"6c",	--5260
		x"58",	--5261
		x"3e",	--5262
		x"14",	--5263
		x"1e",	--5264
		x"17",	--5265
		x"20",	--5266
		x"08",	--5267
		x"38",	--5268
		x"1a",	--5269
		x"19",	--5270
		x"28",	--5271
		x"89",	--5272
		x"89",	--5273
		x"89",	--5274
		x"89",	--5275
		x"1c",	--5276
		x"28",	--5277
		x"0d",	--5278
		x"0e",	--5279
		x"0f",	--5280
		x"b0",	--5281
		x"56",	--5282
		x"0b",	--5283
		x"3e",	--5284
		x"0a",	--5285
		x"05",	--5286
		x"7b",	--5287
		x"30",	--5288
		x"c8",	--5289
		x"00",	--5290
		x"0c",	--5291
		x"4b",	--5292
		x"d1",	--5293
		x"01",	--5294
		x"03",	--5295
		x"7a",	--5296
		x"37",	--5297
		x"02",	--5298
		x"7a",	--5299
		x"57",	--5300
		x"4a",	--5301
		x"c8",	--5302
		x"00",	--5303
		x"06",	--5304
		x"36",	--5305
		x"1c",	--5306
		x"28",	--5307
		x"0d",	--5308
		x"0e",	--5309
		x"0f",	--5310
		x"b0",	--5311
		x"20",	--5312
		x"04",	--5313
		x"07",	--5314
		x"38",	--5315
		x"0e",	--5316
		x"d0",	--5317
		x"0f",	--5318
		x"ce",	--5319
		x"81",	--5320
		x"1e",	--5321
		x"81",	--5322
		x"20",	--5323
		x"2c",	--5324
		x"17",	--5325
		x"1e",	--5326
		x"08",	--5327
		x"38",	--5328
		x"1a",	--5329
		x"1e",	--5330
		x"28",	--5331
		x"0f",	--5332
		x"b0",	--5333
		x"c6",	--5334
		x"0d",	--5335
		x"3f",	--5336
		x"0a",	--5337
		x"05",	--5338
		x"7d",	--5339
		x"30",	--5340
		x"c8",	--5341
		x"00",	--5342
		x"0c",	--5343
		x"4d",	--5344
		x"d1",	--5345
		x"01",	--5346
		x"03",	--5347
		x"7c",	--5348
		x"37",	--5349
		x"02",	--5350
		x"7c",	--5351
		x"57",	--5352
		x"4c",	--5353
		x"c8",	--5354
		x"00",	--5355
		x"06",	--5356
		x"36",	--5357
		x"1e",	--5358
		x"28",	--5359
		x"0f",	--5360
		x"b0",	--5361
		x"ac",	--5362
		x"07",	--5363
		x"38",	--5364
		x"0f",	--5365
		x"db",	--5366
		x"81",	--5367
		x"1e",	--5368
		x"b1",	--5369
		x"0a",	--5370
		x"28",	--5371
		x"02",	--5372
		x"c1",	--5373
		x"02",	--5374
		x"c1",	--5375
		x"2e",	--5376
		x"2a",	--5377
		x"0f",	--5378
		x"3f",	--5379
		x"1c",	--5380
		x"81",	--5381
		x"42",	--5382
		x"1a",	--5383
		x"1c",	--5384
		x"8a",	--5385
		x"8a",	--5386
		x"8a",	--5387
		x"8a",	--5388
		x"81",	--5389
		x"44",	--5390
		x"81",	--5391
		x"46",	--5392
		x"0a",	--5393
		x"8a",	--5394
		x"8a",	--5395
		x"8a",	--5396
		x"8a",	--5397
		x"81",	--5398
		x"48",	--5399
		x"1c",	--5400
		x"42",	--5401
		x"1d",	--5402
		x"44",	--5403
		x"1c",	--5404
		x"46",	--5405
		x"1d",	--5406
		x"48",	--5407
		x"2c",	--5408
		x"1c",	--5409
		x"26",	--5410
		x"0e",	--5411
		x"e1",	--5412
		x"01",	--5413
		x"5e",	--5414
		x"26",	--5415
		x"4e",	--5416
		x"c1",	--5417
		x"03",	--5418
		x"06",	--5419
		x"c1",	--5420
		x"2a",	--5421
		x"03",	--5422
		x"91",	--5423
		x"26",	--5424
		x"30",	--5425
		x"11",	--5426
		x"04",	--5427
		x"11",	--5428
		x"04",	--5429
		x"1d",	--5430
		x"34",	--5431
		x"0e",	--5432
		x"1e",	--5433
		x"1f",	--5434
		x"3e",	--5435
		x"b0",	--5436
		x"b0",	--5437
		x"21",	--5438
		x"81",	--5439
		x"2c",	--5440
		x"0d",	--5441
		x"7f",	--5442
		x"8f",	--5443
		x"91",	--5444
		x"3c",	--5445
		x"0e",	--5446
		x"0e",	--5447
		x"19",	--5448
		x"40",	--5449
		x"f7",	--5450
		x"81",	--5451
		x"3e",	--5452
		x"81",	--5453
		x"2c",	--5454
		x"07",	--5455
		x"0e",	--5456
		x"91",	--5457
		x"26",	--5458
		x"30",	--5459
		x"d1",	--5460
		x"2e",	--5461
		x"c1",	--5462
		x"2a",	--5463
		x"03",	--5464
		x"05",	--5465
		x"d1",	--5466
		x"2a",	--5467
		x"81",	--5468
		x"26",	--5469
		x"17",	--5470
		x"16",	--5471
		x"40",	--5472
		x"6e",	--5473
		x"4e",	--5474
		x"02",	--5475
		x"30",	--5476
		x"94",	--5477
		x"1f",	--5478
		x"2c",	--5479
		x"31",	--5480
		x"4a",	--5481
		x"34",	--5482
		x"35",	--5483
		x"36",	--5484
		x"37",	--5485
		x"38",	--5486
		x"39",	--5487
		x"3a",	--5488
		x"3b",	--5489
		x"30",	--5490
		x"0d",	--5491
		x"0f",	--5492
		x"04",	--5493
		x"3d",	--5494
		x"03",	--5495
		x"3f",	--5496
		x"1f",	--5497
		x"0e",	--5498
		x"03",	--5499
		x"5d",	--5500
		x"3e",	--5501
		x"1e",	--5502
		x"0d",	--5503
		x"b0",	--5504
		x"ac",	--5505
		x"3d",	--5506
		x"6d",	--5507
		x"02",	--5508
		x"3e",	--5509
		x"1e",	--5510
		x"5d",	--5511
		x"02",	--5512
		x"3f",	--5513
		x"1f",	--5514
		x"30",	--5515
		x"b0",	--5516
		x"e6",	--5517
		x"0f",	--5518
		x"30",	--5519
		x"0b",	--5520
		x"0a",	--5521
		x"09",	--5522
		x"79",	--5523
		x"20",	--5524
		x"0a",	--5525
		x"0b",	--5526
		x"0c",	--5527
		x"0d",	--5528
		x"0e",	--5529
		x"0f",	--5530
		x"0c",	--5531
		x"0d",	--5532
		x"0d",	--5533
		x"06",	--5534
		x"02",	--5535
		x"0c",	--5536
		x"03",	--5537
		x"0c",	--5538
		x"0d",	--5539
		x"1e",	--5540
		x"19",	--5541
		x"f2",	--5542
		x"39",	--5543
		x"3a",	--5544
		x"3b",	--5545
		x"30",	--5546
		x"b0",	--5547
		x"20",	--5548
		x"0e",	--5549
		x"0f",	--5550
		x"30",	--5551
		x"0b",	--5552
		x"0b",	--5553
		x"0f",	--5554
		x"06",	--5555
		x"3b",	--5556
		x"03",	--5557
		x"3e",	--5558
		x"3f",	--5559
		x"1e",	--5560
		x"0f",	--5561
		x"0d",	--5562
		x"05",	--5563
		x"5b",	--5564
		x"3c",	--5565
		x"3d",	--5566
		x"1c",	--5567
		x"0d",	--5568
		x"b0",	--5569
		x"20",	--5570
		x"6b",	--5571
		x"04",	--5572
		x"3c",	--5573
		x"3d",	--5574
		x"1c",	--5575
		x"0d",	--5576
		x"5b",	--5577
		x"04",	--5578
		x"3e",	--5579
		x"3f",	--5580
		x"1e",	--5581
		x"0f",	--5582
		x"3b",	--5583
		x"30",	--5584
		x"b0",	--5585
		x"60",	--5586
		x"0e",	--5587
		x"0f",	--5588
		x"30",	--5589
		x"7c",	--5590
		x"10",	--5591
		x"0d",	--5592
		x"0e",	--5593
		x"0f",	--5594
		x"0e",	--5595
		x"0e",	--5596
		x"02",	--5597
		x"0e",	--5598
		x"1f",	--5599
		x"1c",	--5600
		x"f8",	--5601
		x"30",	--5602
		x"b0",	--5603
		x"ac",	--5604
		x"0f",	--5605
		x"30",	--5606
		x"07",	--5607
		x"06",	--5608
		x"05",	--5609
		x"04",	--5610
		x"30",	--5611
		x"40",	--5612
		x"04",	--5613
		x"05",	--5614
		x"06",	--5615
		x"07",	--5616
		x"08",	--5617
		x"09",	--5618
		x"0a",	--5619
		x"0b",	--5620
		x"0c",	--5621
		x"0d",	--5622
		x"0e",	--5623
		x"0f",	--5624
		x"08",	--5625
		x"09",	--5626
		x"0a",	--5627
		x"0b",	--5628
		x"0b",	--5629
		x"0e",	--5630
		x"08",	--5631
		x"0a",	--5632
		x"0b",	--5633
		x"05",	--5634
		x"09",	--5635
		x"08",	--5636
		x"02",	--5637
		x"08",	--5638
		x"05",	--5639
		x"08",	--5640
		x"09",	--5641
		x"0a",	--5642
		x"0b",	--5643
		x"1c",	--5644
		x"91",	--5645
		x"00",	--5646
		x"e5",	--5647
		x"21",	--5648
		x"34",	--5649
		x"35",	--5650
		x"36",	--5651
		x"37",	--5652
		x"30",	--5653
		x"0b",	--5654
		x"0a",	--5655
		x"09",	--5656
		x"08",	--5657
		x"18",	--5658
		x"0a",	--5659
		x"19",	--5660
		x"0c",	--5661
		x"1a",	--5662
		x"0e",	--5663
		x"1b",	--5664
		x"10",	--5665
		x"b0",	--5666
		x"ce",	--5667
		x"38",	--5668
		x"39",	--5669
		x"3a",	--5670
		x"3b",	--5671
		x"30",	--5672
		x"0b",	--5673
		x"0a",	--5674
		x"09",	--5675
		x"08",	--5676
		x"18",	--5677
		x"0a",	--5678
		x"19",	--5679
		x"0c",	--5680
		x"1a",	--5681
		x"0e",	--5682
		x"1b",	--5683
		x"10",	--5684
		x"b0",	--5685
		x"ce",	--5686
		x"0c",	--5687
		x"0d",	--5688
		x"0e",	--5689
		x"0f",	--5690
		x"38",	--5691
		x"39",	--5692
		x"3a",	--5693
		x"3b",	--5694
		x"30",	--5695
		x"0b",	--5696
		x"0a",	--5697
		x"09",	--5698
		x"08",	--5699
		x"07",	--5700
		x"18",	--5701
		x"0c",	--5702
		x"19",	--5703
		x"0e",	--5704
		x"1a",	--5705
		x"10",	--5706
		x"1b",	--5707
		x"12",	--5708
		x"b0",	--5709
		x"ce",	--5710
		x"17",	--5711
		x"14",	--5712
		x"87",	--5713
		x"00",	--5714
		x"87",	--5715
		x"02",	--5716
		x"87",	--5717
		x"04",	--5718
		x"87",	--5719
		x"06",	--5720
		x"37",	--5721
		x"38",	--5722
		x"39",	--5723
		x"3a",	--5724
		x"3b",	--5725
		x"30",	--5726
		x"00",	--5727
		x"32",	--5728
		x"f0",	--5729
		x"fd",	--5730
		x"53",	--5731
		x"6f",	--5732
		x"0d",	--5733
		x"00",	--5734
		x"6f",	--5735
		x"72",	--5736
		x"63",	--5737
		x"20",	--5738
		x"73",	--5739
		x"67",	--5740
		x"3a",	--5741
		x"0a",	--5742
		x"09",	--5743
		x"63",	--5744
		x"4c",	--5745
		x"46",	--5746
		x"20",	--5747
		x"49",	--5748
		x"48",	--5749
		x"20",	--5750
		x"54",	--5751
		x"4d",	--5752
		x"4f",	--5753
		x"54",	--5754
		x"0d",	--5755
		x"00",	--5756
		x"64",	--5757
		x"25",	--5758
		x"0d",	--5759
		x"00",	--5760
		x"6f",	--5761
		x"20",	--5762
		x"6d",	--5763
		x"6c",	--5764
		x"6d",	--5765
		x"6e",	--5766
		x"65",	--5767
		x"20",	--5768
		x"65",	--5769
		x"0d",	--5770
		x"00",	--5771
		x"61",	--5772
		x"74",	--5773
		x"6e",	--5774
		x"20",	--5775
		x"6f",	--5776
		x"20",	--5777
		x"20",	--5778
		x"65",	--5779
		x"20",	--5780
		x"62",	--5781
		x"6e",	--5782
		x"66",	--5783
		x"6c",	--5784
		x"0d",	--5785
		x"00",	--5786
		x"65",	--5787
		x"73",	--5788
		x"6f",	--5789
		x"6c",	--5790
		x"20",	--5791
		x"6f",	--5792
		x"20",	--5793
		x"65",	--5794
		x"20",	--5795
		x"68",	--5796
		x"74",	--5797
		x"0a",	--5798
		x"53",	--5799
		x"6f",	--5800
		x"0d",	--5801
		x"00",	--5802
		x"72",	--5803
		x"6f",	--5804
		x"3a",	--5805
		x"6d",	--5806
		x"73",	--5807
		x"69",	--5808
		x"67",	--5809
		x"61",	--5810
		x"67",	--5811
		x"6d",	--5812
		x"6e",	--5813
		x"0d",	--5814
		x"00",	--5815
		x"6f",	--5816
		x"72",	--5817
		x"63",	--5818
		x"20",	--5819
		x"73",	--5820
		x"67",	--5821
		x"3a",	--5822
		x"0a",	--5823
		x"09",	--5824
		x"73",	--5825
		x"4c",	--5826
		x"46",	--5827
		x"20",	--5828
		x"49",	--5829
		x"48",	--5830
		x"20",	--5831
		x"54",	--5832
		x"4d",	--5833
		x"4f",	--5834
		x"54",	--5835
		x"0d",	--5836
		x"00",	--5837
		x"64",	--5838
		x"25",	--5839
		x"0d",	--5840
		x"00",	--5841
		x"6c",	--5842
		x"20",	--5843
		x"6c",	--5844
		x"00",	--5845
		x"73",	--5846
		x"0a",	--5847
		x"25",	--5848
		x"20",	--5849
		x"64",	--5850
		x"0a",	--5851
		x"46",	--5852
		x"6e",	--5853
		x"74",	--5854
		x"7c",	--5855
		x"84",	--5856
		x"8c",	--5857
		x"5e",	--5858
		x"66",	--5859
		x"0d",	--5860
		x"3d",	--5861
		x"3d",	--5862
		x"3d",	--5863
		x"20",	--5864
		x"61",	--5865
		x"63",	--5866
		x"6c",	--5867
		x"4d",	--5868
		x"55",	--5869
		x"3d",	--5870
		x"3d",	--5871
		x"3d",	--5872
		x"0d",	--5873
		x"00",	--5874
		x"6e",	--5875
		x"65",	--5876
		x"61",	--5877
		x"74",	--5878
		x"76",	--5879
		x"20",	--5880
		x"6f",	--5881
		x"65",	--5882
		x"77",	--5883
		x"69",	--5884
		x"65",	--5885
		x"72",	--5886
		x"61",	--5887
		x"00",	--5888
		x"75",	--5889
		x"7a",	--5890
		x"72",	--5891
		x"70",	--5892
		x"6d",	--5893
		x"65",	--5894
		x"63",	--5895
		x"64",	--5896
		x"72",	--5897
		x"73",	--5898
		x"65",	--5899
		x"64",	--5900
		x"63",	--5901
		x"6e",	--5902
		x"72",	--5903
		x"6c",	--5904
		x"65",	--5905
		x"00",	--5906
		x"70",	--5907
		x"65",	--5908
		x"20",	--5909
		x"6f",	--5910
		x"66",	--5911
		x"67",	--5912
		x"72",	--5913
		x"74",	--5914
		x"6f",	--5915
		x"00",	--5916
		x"6f",	--5917
		x"74",	--5918
		x"6f",	--5919
		x"64",	--5920
		x"72",	--5921
		x"0d",	--5922
		x"00",	--5923
		x"20",	--5924
		x"00",	--5925
		x"63",	--5926
		x"55",	--5927
		x"0d",	--5928
		x"00",	--5929
		x"4f",	--5930
		x"4e",	--5931
		x"0a",	--5932
		x"52",	--5933
		x"47",	--5934
		x"54",	--5935
		x"0a",	--5936
		x"4c",	--5937
		x"46",	--5938
		x"0d",	--5939
		x"00",	--5940
		x"77",	--5941
		x"69",	--5942
		x"65",	--5943
		x"0d",	--5944
		x"65",	--5945
		x"72",	--5946
		x"72",	--5947
		x"20",	--5948
		x"69",	--5949
		x"73",	--5950
		x"6e",	--5951
		x"20",	--5952
		x"72",	--5953
		x"75",	--5954
		x"65",	--5955
		x"74",	--5956
		x"0a",	--5957
		x"63",	--5958
		x"72",	--5959
		x"65",	--5960
		x"74",	--5961
		x"75",	--5962
		x"61",	--5963
		x"65",	--5964
		x"0d",	--5965
		x"00",	--5966
		x"25",	--5967
		x"20",	--5968
		x"45",	--5969
		x"49",	--5970
		x"54",	--5971
		x"52",	--5972
		x"56",	--5973
		x"4c",	--5974
		x"45",	--5975
		x"0a",	--5976
		x"72",	--5977
		x"25",	--5978
		x"20",	--5979
		x"3d",	--5980
		x"64",	--5981
		x"0a",	--5982
		x"09",	--5983
		x"73",	--5984
		x"52",	--5985
		x"47",	--5986
		x"53",	--5987
		x"45",	--5988
		x"0d",	--5989
		x"00",	--5990
		x"65",	--5991
		x"64",	--5992
		x"0d",	--5993
		x"25",	--5994
		x"20",	--5995
		x"73",	--5996
		x"6e",	--5997
		x"74",	--5998
		x"61",	--5999
		x"6e",	--6000
		x"6d",	--6001
		x"65",	--6002
		x"0d",	--6003
		x"00",	--6004
		x"63",	--6005
		x"25",	--6006
		x"0d",	--6007
		x"00",	--6008
		x"63",	--6009
		x"20",	--6010
		x"6f",	--6011
		x"73",	--6012
		x"63",	--6013
		x"20",	--6014
		x"6f",	--6015
		x"6d",	--6016
		x"6e",	--6017
		x"0d",	--6018
		x"00",	--6019
		x"2e",	--6020
		x"5c",	--6021
		x"5c",	--6022
		x"5c",	--6023
		x"5c",	--6024
		x"5c",	--6025
		x"5c",	--6026
		x"5c",	--6027
		x"5c",	--6028
		x"5c",	--6029
		x"5c",	--6030
		x"5c",	--6031
		x"5c",	--6032
		x"5c",	--6033
		x"5c",	--6034
		x"5c",	--6035
		x"5c",	--6036
		x"5c",	--6037
		x"5c",	--6038
		x"5c",	--6039
		x"5c",	--6040
		x"5c",	--6041
		x"5c",	--6042
		x"5c",	--6043
		x"5c",	--6044
		x"5c",	--6045
		x"5c",	--6046
		x"5c",	--6047
		x"5c",	--6048
		x"20",	--6049
		x"5c",	--6050
		x"5c",	--6051
		x"5c",	--6052
		x"5c",	--6053
		x"5c",	--6054
		x"5c",	--6055
		x"5c",	--6056
		x"5c",	--6057
		x"5c",	--6058
		x"5c",	--6059
		x"5c",	--6060
		x"5c",	--6061
		x"5c",	--6062
		x"5c",	--6063
		x"5c",	--6064
		x"5c",	--6065
		x"5c",	--6066
		x"5c",	--6067
		x"5c",	--6068
		x"5c",	--6069
		x"5c",	--6070
		x"5c",	--6071
		x"5c",	--6072
		x"5c",	--6073
		x"5c",	--6074
		x"5c",	--6075
		x"5c",	--6076
		x"5c",	--6077
		x"5c",	--6078
		x"5c",	--6079
		x"5c",	--6080
		x"12",	--6081
		x"04",	--6082
		x"f6",	--6083
		x"5c",	--6084
		x"5c",	--6085
		x"5c",	--6086
		x"5c",	--6087
		x"5c",	--6088
		x"5c",	--6089
		x"5c",	--6090
		x"de",	--6091
		x"5c",	--6092
		x"cc",	--6093
		x"5c",	--6094
		x"5c",	--6095
		x"5c",	--6096
		x"5c",	--6097
		x"b0",	--6098
		x"5c",	--6099
		x"5c",	--6100
		x"5c",	--6101
		x"a2",	--6102
		x"90",	--6103
		x"30",	--6104
		x"32",	--6105
		x"34",	--6106
		x"36",	--6107
		x"38",	--6108
		x"61",	--6109
		x"63",	--6110
		x"65",	--6111
		x"00",	--6112
		x"00",	--6113
		x"00",	--6114
		x"00",	--6115
		x"00",	--6116
		x"00",	--6117
		x"02",	--6118
		x"03",	--6119
		x"03",	--6120
		x"04",	--6121
		x"04",	--6122
		x"04",	--6123
		x"04",	--6124
		x"05",	--6125
		x"05",	--6126
		x"05",	--6127
		x"05",	--6128
		x"05",	--6129
		x"05",	--6130
		x"05",	--6131
		x"05",	--6132
		x"06",	--6133
		x"06",	--6134
		x"06",	--6135
		x"06",	--6136
		x"06",	--6137
		x"06",	--6138
		x"06",	--6139
		x"06",	--6140
		x"06",	--6141
		x"06",	--6142
		x"06",	--6143
		x"06",	--6144
		x"06",	--6145
		x"06",	--6146
		x"06",	--6147
		x"06",	--6148
		x"07",	--6149
		x"07",	--6150
		x"07",	--6151
		x"07",	--6152
		x"07",	--6153
		x"07",	--6154
		x"07",	--6155
		x"07",	--6156
		x"07",	--6157
		x"07",	--6158
		x"07",	--6159
		x"07",	--6160
		x"07",	--6161
		x"07",	--6162
		x"07",	--6163
		x"07",	--6164
		x"07",	--6165
		x"07",	--6166
		x"07",	--6167
		x"07",	--6168
		x"07",	--6169
		x"07",	--6170
		x"07",	--6171
		x"07",	--6172
		x"07",	--6173
		x"07",	--6174
		x"07",	--6175
		x"07",	--6176
		x"07",	--6177
		x"07",	--6178
		x"07",	--6179
		x"07",	--6180
		x"08",	--6181
		x"08",	--6182
		x"08",	--6183
		x"08",	--6184
		x"08",	--6185
		x"08",	--6186
		x"08",	--6187
		x"08",	--6188
		x"08",	--6189
		x"08",	--6190
		x"08",	--6191
		x"08",	--6192
		x"08",	--6193
		x"08",	--6194
		x"08",	--6195
		x"08",	--6196
		x"08",	--6197
		x"08",	--6198
		x"08",	--6199
		x"08",	--6200
		x"08",	--6201
		x"08",	--6202
		x"08",	--6203
		x"08",	--6204
		x"08",	--6205
		x"08",	--6206
		x"08",	--6207
		x"08",	--6208
		x"08",	--6209
		x"08",	--6210
		x"08",	--6211
		x"08",	--6212
		x"08",	--6213
		x"08",	--6214
		x"08",	--6215
		x"08",	--6216
		x"08",	--6217
		x"08",	--6218
		x"08",	--6219
		x"08",	--6220
		x"08",	--6221
		x"08",	--6222
		x"08",	--6223
		x"08",	--6224
		x"08",	--6225
		x"08",	--6226
		x"08",	--6227
		x"08",	--6228
		x"08",	--6229
		x"08",	--6230
		x"08",	--6231
		x"08",	--6232
		x"08",	--6233
		x"08",	--6234
		x"08",	--6235
		x"08",	--6236
		x"08",	--6237
		x"08",	--6238
		x"08",	--6239
		x"08",	--6240
		x"08",	--6241
		x"08",	--6242
		x"08",	--6243
		x"08",	--6244
		x"28",	--6245
		x"75",	--6246
		x"6c",	--6247
		x"00",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"68",	--6252
		x"6c",	--6253
		x"00",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"3c",	--8176
		x"3c",	--8177
		x"3c",	--8178
		x"3c",	--8179
		x"3c",	--8180
		x"3c",	--8181
		x"3c",	--8182
		x"38",	--8183
		x"8a",	--8184
		x"3c",	--8185
		x"3c",	--8186
		x"3c",	--8187
		x"3c",	--8188
		x"3c",	--8189
		x"3c",	--8190
		x"00");	--8191
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"f0",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"d3",	--44
		x"12",	--45
		x"cd",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"ed",	--50
		x"12",	--51
		x"d2",	--52
		x"53",	--53
		x"40",	--54
		x"ed",	--55
		x"40",	--56
		x"c9",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"ce",	--61
		x"40",	--62
		x"ed",	--63
		x"40",	--64
		x"ca",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"ce",	--69
		x"40",	--70
		x"ed",	--71
		x"40",	--72
		x"cb",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"ce",	--77
		x"40",	--78
		x"ee",	--79
		x"40",	--80
		x"c3",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"ce",	--85
		x"40",	--86
		x"ee",	--87
		x"40",	--88
		x"c6",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"ce",	--93
		x"40",	--94
		x"ee",	--95
		x"40",	--96
		x"c8",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"ce",	--101
		x"40",	--102
		x"ee",	--103
		x"40",	--104
		x"c3",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"ce",	--109
		x"40",	--110
		x"ee",	--111
		x"40",	--112
		x"c5",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"ce",	--117
		x"40",	--118
		x"ee",	--119
		x"40",	--120
		x"c5",	--121
		x"40",	--122
		x"00",	--123
		x"12",	--124
		x"ce",	--125
		x"43",	--126
		x"43",	--127
		x"12",	--128
		x"cd",	--129
		x"43",	--130
		x"40",	--131
		x"4e",	--132
		x"40",	--133
		x"01",	--134
		x"41",	--135
		x"50",	--136
		x"00",	--137
		x"12",	--138
		x"cc",	--139
		x"41",	--140
		x"50",	--141
		x"00",	--142
		x"12",	--143
		x"cd",	--144
		x"43",	--145
		x"40",	--146
		x"4e",	--147
		x"40",	--148
		x"01",	--149
		x"41",	--150
		x"50",	--151
		x"00",	--152
		x"12",	--153
		x"cc",	--154
		x"41",	--155
		x"50",	--156
		x"00",	--157
		x"12",	--158
		x"cd",	--159
		x"41",	--160
		x"50",	--161
		x"00",	--162
		x"41",	--163
		x"50",	--164
		x"00",	--165
		x"12",	--166
		x"c6",	--167
		x"40",	--168
		x"01",	--169
		x"41",	--170
		x"52",	--171
		x"12",	--172
		x"d0",	--173
		x"40",	--174
		x"01",	--175
		x"41",	--176
		x"53",	--177
		x"12",	--178
		x"d0",	--179
		x"41",	--180
		x"53",	--181
		x"41",	--182
		x"52",	--183
		x"12",	--184
		x"c7",	--185
		x"41",	--186
		x"50",	--187
		x"00",	--188
		x"41",	--189
		x"50",	--190
		x"00",	--191
		x"12",	--192
		x"c7",	--193
		x"12",	--194
		x"ce",	--195
		x"40",	--196
		x"01",	--197
		x"41",	--198
		x"12",	--199
		x"d0",	--200
		x"41",	--201
		x"12",	--202
		x"c3",	--203
		x"40",	--204
		x"00",	--205
		x"40",	--206
		x"11",	--207
		x"41",	--208
		x"12",	--209
		x"d0",	--210
		x"12",	--211
		x"12",	--212
		x"12",	--213
		x"39",	--214
		x"12",	--215
		x"b7",	--216
		x"12",	--217
		x"3a",	--218
		x"12",	--219
		x"49",	--220
		x"40",	--221
		x"00",	--222
		x"41",	--223
		x"50",	--224
		x"00",	--225
		x"41",	--226
		x"50",	--227
		x"00",	--228
		x"41",	--229
		x"50",	--230
		x"00",	--231
		x"12",	--232
		x"c5",	--233
		x"50",	--234
		x"00",	--235
		x"12",	--236
		x"12",	--237
		x"12",	--238
		x"39",	--239
		x"12",	--240
		x"b7",	--241
		x"12",	--242
		x"3a",	--243
		x"12",	--244
		x"49",	--245
		x"40",	--246
		x"00",	--247
		x"41",	--248
		x"50",	--249
		x"00",	--250
		x"41",	--251
		x"50",	--252
		x"00",	--253
		x"41",	--254
		x"50",	--255
		x"00",	--256
		x"12",	--257
		x"c5",	--258
		x"50",	--259
		x"00",	--260
		x"41",	--261
		x"50",	--262
		x"00",	--263
		x"41",	--264
		x"50",	--265
		x"00",	--266
		x"12",	--267
		x"c3",	--268
		x"12",	--269
		x"c3",	--270
		x"40",	--271
		x"ff",	--272
		x"00",	--273
		x"d2",	--274
		x"43",	--275
		x"43",	--276
		x"3c",	--277
		x"43",	--278
		x"3c",	--279
		x"43",	--280
		x"3c",	--281
		x"43",	--282
		x"12",	--283
		x"d3",	--284
		x"93",	--285
		x"27",	--286
		x"12",	--287
		x"d3",	--288
		x"93",	--289
		x"20",	--290
		x"90",	--291
		x"00",	--292
		x"24",	--293
		x"90",	--294
		x"00",	--295
		x"27",	--296
		x"92",	--297
		x"20",	--298
		x"3c",	--299
		x"12",	--300
		x"ee",	--301
		x"12",	--302
		x"d2",	--303
		x"53",	--304
		x"40",	--305
		x"00",	--306
		x"51",	--307
		x"5f",	--308
		x"43",	--309
		x"00",	--310
		x"4f",	--311
		x"41",	--312
		x"00",	--313
		x"12",	--314
		x"ce",	--315
		x"43",	--316
		x"3f",	--317
		x"93",	--318
		x"27",	--319
		x"53",	--320
		x"12",	--321
		x"ee",	--322
		x"12",	--323
		x"d2",	--324
		x"53",	--325
		x"3f",	--326
		x"90",	--327
		x"00",	--328
		x"2f",	--329
		x"93",	--330
		x"02",	--331
		x"24",	--332
		x"4f",	--333
		x"11",	--334
		x"12",	--335
		x"12",	--336
		x"ee",	--337
		x"4f",	--338
		x"00",	--339
		x"12",	--340
		x"d2",	--341
		x"52",	--342
		x"41",	--343
		x"00",	--344
		x"40",	--345
		x"00",	--346
		x"51",	--347
		x"5a",	--348
		x"4f",	--349
		x"00",	--350
		x"53",	--351
		x"3f",	--352
		x"93",	--353
		x"20",	--354
		x"90",	--355
		x"00",	--356
		x"23",	--357
		x"3f",	--358
		x"93",	--359
		x"23",	--360
		x"90",	--361
		x"00",	--362
		x"24",	--363
		x"90",	--364
		x"00",	--365
		x"34",	--366
		x"90",	--367
		x"00",	--368
		x"23",	--369
		x"3c",	--370
		x"90",	--371
		x"00",	--372
		x"24",	--373
		x"90",	--374
		x"00",	--375
		x"23",	--376
		x"3c",	--377
		x"12",	--378
		x"ee",	--379
		x"12",	--380
		x"d2",	--381
		x"53",	--382
		x"12",	--383
		x"c4",	--384
		x"43",	--385
		x"3f",	--386
		x"12",	--387
		x"ee",	--388
		x"12",	--389
		x"d2",	--390
		x"53",	--391
		x"12",	--392
		x"c4",	--393
		x"43",	--394
		x"3f",	--395
		x"12",	--396
		x"ee",	--397
		x"12",	--398
		x"d2",	--399
		x"53",	--400
		x"12",	--401
		x"c4",	--402
		x"43",	--403
		x"3f",	--404
		x"12",	--405
		x"ee",	--406
		x"12",	--407
		x"d2",	--408
		x"53",	--409
		x"12",	--410
		x"c4",	--411
		x"43",	--412
		x"3f",	--413
		x"40",	--414
		x"ec",	--415
		x"4f",	--416
		x"02",	--417
		x"41",	--418
		x"12",	--419
		x"12",	--420
		x"82",	--421
		x"4f",	--422
		x"4e",	--423
		x"93",	--424
		x"38",	--425
		x"41",	--426
		x"4b",	--427
		x"00",	--428
		x"12",	--429
		x"cb",	--430
		x"4f",	--431
		x"93",	--432
		x"24",	--433
		x"41",	--434
		x"4b",	--435
		x"00",	--436
		x"4d",	--437
		x"00",	--438
		x"12",	--439
		x"cb",	--440
		x"4f",	--441
		x"41",	--442
		x"00",	--443
		x"42",	--444
		x"02",	--445
		x"12",	--446
		x"d0",	--447
		x"43",	--448
		x"52",	--449
		x"41",	--450
		x"41",	--451
		x"41",	--452
		x"40",	--453
		x"00",	--454
		x"40",	--455
		x"11",	--456
		x"3f",	--457
		x"40",	--458
		x"11",	--459
		x"3f",	--460
		x"43",	--461
		x"42",	--462
		x"02",	--463
		x"12",	--464
		x"c6",	--465
		x"43",	--466
		x"42",	--467
		x"02",	--468
		x"12",	--469
		x"c6",	--470
		x"12",	--471
		x"ec",	--472
		x"12",	--473
		x"d2",	--474
		x"53",	--475
		x"41",	--476
		x"93",	--477
		x"02",	--478
		x"24",	--479
		x"42",	--480
		x"02",	--481
		x"12",	--482
		x"c6",	--483
		x"42",	--484
		x"02",	--485
		x"12",	--486
		x"c6",	--487
		x"41",	--488
		x"43",	--489
		x"40",	--490
		x"c3",	--491
		x"12",	--492
		x"cf",	--493
		x"4f",	--494
		x"02",	--495
		x"3f",	--496
		x"4f",	--497
		x"02",	--498
		x"4e",	--499
		x"02",	--500
		x"41",	--501
		x"12",	--502
		x"12",	--503
		x"83",	--504
		x"4e",	--505
		x"90",	--506
		x"00",	--507
		x"38",	--508
		x"20",	--509
		x"41",	--510
		x"4b",	--511
		x"00",	--512
		x"12",	--513
		x"cc",	--514
		x"4f",	--515
		x"41",	--516
		x"4b",	--517
		x"00",	--518
		x"12",	--519
		x"cc",	--520
		x"4f",	--521
		x"12",	--522
		x"12",	--523
		x"12",	--524
		x"ec",	--525
		x"12",	--526
		x"d2",	--527
		x"50",	--528
		x"00",	--529
		x"4a",	--530
		x"42",	--531
		x"02",	--532
		x"12",	--533
		x"c6",	--534
		x"4b",	--535
		x"42",	--536
		x"02",	--537
		x"12",	--538
		x"c6",	--539
		x"43",	--540
		x"53",	--541
		x"41",	--542
		x"41",	--543
		x"41",	--544
		x"41",	--545
		x"4b",	--546
		x"00",	--547
		x"12",	--548
		x"cb",	--549
		x"43",	--550
		x"4f",	--551
		x"42",	--552
		x"02",	--553
		x"12",	--554
		x"cf",	--555
		x"3f",	--556
		x"12",	--557
		x"ec",	--558
		x"12",	--559
		x"d2",	--560
		x"4b",	--561
		x"00",	--562
		x"12",	--563
		x"ec",	--564
		x"12",	--565
		x"d2",	--566
		x"52",	--567
		x"43",	--568
		x"3f",	--569
		x"40",	--570
		x"ff",	--571
		x"42",	--572
		x"02",	--573
		x"12",	--574
		x"c6",	--575
		x"40",	--576
		x"00",	--577
		x"42",	--578
		x"02",	--579
		x"12",	--580
		x"c6",	--581
		x"43",	--582
		x"40",	--583
		x"00",	--584
		x"42",	--585
		x"02",	--586
		x"12",	--587
		x"cf",	--588
		x"41",	--589
		x"40",	--590
		x"00",	--591
		x"42",	--592
		x"02",	--593
		x"12",	--594
		x"c6",	--595
		x"40",	--596
		x"ff",	--597
		x"42",	--598
		x"02",	--599
		x"12",	--600
		x"c6",	--601
		x"43",	--602
		x"40",	--603
		x"00",	--604
		x"42",	--605
		x"02",	--606
		x"12",	--607
		x"cf",	--608
		x"41",	--609
		x"40",	--610
		x"ff",	--611
		x"42",	--612
		x"02",	--613
		x"12",	--614
		x"c6",	--615
		x"40",	--616
		x"ff",	--617
		x"42",	--618
		x"02",	--619
		x"12",	--620
		x"c6",	--621
		x"43",	--622
		x"40",	--623
		x"00",	--624
		x"42",	--625
		x"02",	--626
		x"12",	--627
		x"cf",	--628
		x"41",	--629
		x"40",	--630
		x"00",	--631
		x"42",	--632
		x"02",	--633
		x"12",	--634
		x"c6",	--635
		x"40",	--636
		x"00",	--637
		x"42",	--638
		x"02",	--639
		x"12",	--640
		x"c6",	--641
		x"43",	--642
		x"40",	--643
		x"00",	--644
		x"42",	--645
		x"02",	--646
		x"12",	--647
		x"cf",	--648
		x"41",	--649
		x"12",	--650
		x"ed",	--651
		x"12",	--652
		x"d2",	--653
		x"53",	--654
		x"43",	--655
		x"41",	--656
		x"40",	--657
		x"c0",	--658
		x"01",	--659
		x"40",	--660
		x"00",	--661
		x"01",	--662
		x"40",	--663
		x"02",	--664
		x"01",	--665
		x"12",	--666
		x"ed",	--667
		x"12",	--668
		x"d2",	--669
		x"43",	--670
		x"01",	--671
		x"40",	--672
		x"ed",	--673
		x"00",	--674
		x"12",	--675
		x"d2",	--676
		x"53",	--677
		x"43",	--678
		x"41",	--679
		x"12",	--680
		x"12",	--681
		x"12",	--682
		x"4f",	--683
		x"4f",	--684
		x"00",	--685
		x"12",	--686
		x"d0",	--687
		x"4e",	--688
		x"4f",	--689
		x"89",	--690
		x"00",	--691
		x"79",	--692
		x"00",	--693
		x"12",	--694
		x"db",	--695
		x"4a",	--696
		x"00",	--697
		x"4b",	--698
		x"00",	--699
		x"4e",	--700
		x"4f",	--701
		x"49",	--702
		x"12",	--703
		x"ca",	--704
		x"43",	--705
		x"40",	--706
		x"3f",	--707
		x"12",	--708
		x"d6",	--709
		x"4e",	--710
		x"4f",	--711
		x"40",	--712
		x"66",	--713
		x"40",	--714
		x"3f",	--715
		x"12",	--716
		x"da",	--717
		x"93",	--718
		x"24",	--719
		x"34",	--720
		x"40",	--721
		x"cc",	--722
		x"40",	--723
		x"3d",	--724
		x"4a",	--725
		x"4b",	--726
		x"12",	--727
		x"db",	--728
		x"93",	--729
		x"34",	--730
		x"40",	--731
		x"cc",	--732
		x"40",	--733
		x"3d",	--734
		x"4a",	--735
		x"4b",	--736
		x"49",	--737
		x"00",	--738
		x"12",	--739
		x"cd",	--740
		x"41",	--741
		x"41",	--742
		x"41",	--743
		x"41",	--744
		x"40",	--745
		x"66",	--746
		x"40",	--747
		x"3f",	--748
		x"3f",	--749
		x"12",	--750
		x"12",	--751
		x"4f",	--752
		x"4c",	--753
		x"4e",	--754
		x"00",	--755
		x"4d",	--756
		x"00",	--757
		x"12",	--758
		x"00",	--759
		x"12",	--760
		x"00",	--761
		x"12",	--762
		x"00",	--763
		x"12",	--764
		x"00",	--765
		x"41",	--766
		x"00",	--767
		x"41",	--768
		x"00",	--769
		x"12",	--770
		x"c9",	--771
		x"52",	--772
		x"4a",	--773
		x"00",	--774
		x"4b",	--775
		x"40",	--776
		x"c5",	--777
		x"12",	--778
		x"cf",	--779
		x"4f",	--780
		x"00",	--781
		x"41",	--782
		x"41",	--783
		x"41",	--784
		x"12",	--785
		x"4f",	--786
		x"4f",	--787
		x"00",	--788
		x"12",	--789
		x"d0",	--790
		x"4e",	--791
		x"00",	--792
		x"4f",	--793
		x"00",	--794
		x"43",	--795
		x"4b",	--796
		x"00",	--797
		x"4b",	--798
		x"00",	--799
		x"12",	--800
		x"cf",	--801
		x"41",	--802
		x"41",	--803
		x"12",	--804
		x"4f",	--805
		x"43",	--806
		x"40",	--807
		x"3f",	--808
		x"4f",	--809
		x"00",	--810
		x"12",	--811
		x"cd",	--812
		x"4b",	--813
		x"00",	--814
		x"12",	--815
		x"cf",	--816
		x"41",	--817
		x"41",	--818
		x"12",	--819
		x"4f",	--820
		x"4e",	--821
		x"10",	--822
		x"11",	--823
		x"10",	--824
		x"11",	--825
		x"4d",	--826
		x"12",	--827
		x"db",	--828
		x"4e",	--829
		x"4f",	--830
		x"4b",	--831
		x"12",	--832
		x"ca",	--833
		x"41",	--834
		x"41",	--835
		x"12",	--836
		x"12",	--837
		x"43",	--838
		x"40",	--839
		x"3f",	--840
		x"4a",	--841
		x"4b",	--842
		x"42",	--843
		x"02",	--844
		x"12",	--845
		x"cd",	--846
		x"4a",	--847
		x"4b",	--848
		x"42",	--849
		x"02",	--850
		x"12",	--851
		x"cd",	--852
		x"12",	--853
		x"ed",	--854
		x"12",	--855
		x"d2",	--856
		x"53",	--857
		x"41",	--858
		x"41",	--859
		x"41",	--860
		x"4f",	--861
		x"02",	--862
		x"4e",	--863
		x"02",	--864
		x"41",	--865
		x"12",	--866
		x"12",	--867
		x"83",	--868
		x"4f",	--869
		x"4e",	--870
		x"93",	--871
		x"02",	--872
		x"24",	--873
		x"90",	--874
		x"00",	--875
		x"38",	--876
		x"20",	--877
		x"41",	--878
		x"4b",	--879
		x"00",	--880
		x"12",	--881
		x"cb",	--882
		x"4f",	--883
		x"41",	--884
		x"4b",	--885
		x"00",	--886
		x"12",	--887
		x"cb",	--888
		x"4f",	--889
		x"12",	--890
		x"12",	--891
		x"12",	--892
		x"ed",	--893
		x"12",	--894
		x"d2",	--895
		x"50",	--896
		x"00",	--897
		x"4a",	--898
		x"43",	--899
		x"12",	--900
		x"dc",	--901
		x"43",	--902
		x"40",	--903
		x"42",	--904
		x"12",	--905
		x"d9",	--906
		x"4e",	--907
		x"4f",	--908
		x"43",	--909
		x"40",	--910
		x"3f",	--911
		x"12",	--912
		x"d7",	--913
		x"4e",	--914
		x"4f",	--915
		x"42",	--916
		x"02",	--917
		x"12",	--918
		x"cd",	--919
		x"4b",	--920
		x"43",	--921
		x"12",	--922
		x"dc",	--923
		x"43",	--924
		x"40",	--925
		x"42",	--926
		x"12",	--927
		x"d9",	--928
		x"4e",	--929
		x"4f",	--930
		x"42",	--931
		x"02",	--932
		x"12",	--933
		x"cd",	--934
		x"43",	--935
		x"53",	--936
		x"41",	--937
		x"41",	--938
		x"41",	--939
		x"41",	--940
		x"4b",	--941
		x"00",	--942
		x"12",	--943
		x"cb",	--944
		x"43",	--945
		x"4f",	--946
		x"42",	--947
		x"02",	--948
		x"12",	--949
		x"cf",	--950
		x"3f",	--951
		x"43",	--952
		x"40",	--953
		x"c6",	--954
		x"12",	--955
		x"cf",	--956
		x"4f",	--957
		x"02",	--958
		x"3f",	--959
		x"12",	--960
		x"ed",	--961
		x"12",	--962
		x"d2",	--963
		x"40",	--964
		x"ed",	--965
		x"00",	--966
		x"12",	--967
		x"d2",	--968
		x"4b",	--969
		x"00",	--970
		x"12",	--971
		x"ed",	--972
		x"12",	--973
		x"d2",	--974
		x"52",	--975
		x"43",	--976
		x"3f",	--977
		x"12",	--978
		x"12",	--979
		x"42",	--980
		x"02",	--981
		x"12",	--982
		x"d0",	--983
		x"4e",	--984
		x"4f",	--985
		x"42",	--986
		x"02",	--987
		x"12",	--988
		x"d0",	--989
		x"12",	--990
		x"12",	--991
		x"e3",	--992
		x"e3",	--993
		x"53",	--994
		x"63",	--995
		x"12",	--996
		x"12",	--997
		x"12",	--998
		x"ed",	--999
		x"12",	--1000
		x"02",	--1001
		x"12",	--1002
		x"e2",	--1003
		x"50",	--1004
		x"00",	--1005
		x"12",	--1006
		x"02",	--1007
		x"12",	--1008
		x"ed",	--1009
		x"12",	--1010
		x"d2",	--1011
		x"52",	--1012
		x"41",	--1013
		x"41",	--1014
		x"41",	--1015
		x"4f",	--1016
		x"02",	--1017
		x"4e",	--1018
		x"02",	--1019
		x"41",	--1020
		x"4f",	--1021
		x"02",	--1022
		x"4e",	--1023
		x"02",	--1024
		x"41",	--1025
		x"12",	--1026
		x"12",	--1027
		x"12",	--1028
		x"12",	--1029
		x"83",	--1030
		x"4f",	--1031
		x"4e",	--1032
		x"43",	--1033
		x"00",	--1034
		x"93",	--1035
		x"24",	--1036
		x"93",	--1037
		x"02",	--1038
		x"24",	--1039
		x"43",	--1040
		x"02",	--1041
		x"41",	--1042
		x"4b",	--1043
		x"00",	--1044
		x"12",	--1045
		x"cb",	--1046
		x"4f",	--1047
		x"90",	--1048
		x"00",	--1049
		x"34",	--1050
		x"43",	--1051
		x"49",	--1052
		x"48",	--1053
		x"42",	--1054
		x"02",	--1055
		x"12",	--1056
		x"cf",	--1057
		x"43",	--1058
		x"53",	--1059
		x"41",	--1060
		x"41",	--1061
		x"41",	--1062
		x"41",	--1063
		x"41",	--1064
		x"93",	--1065
		x"02",	--1066
		x"24",	--1067
		x"43",	--1068
		x"02",	--1069
		x"42",	--1070
		x"02",	--1071
		x"12",	--1072
		x"cf",	--1073
		x"43",	--1074
		x"53",	--1075
		x"41",	--1076
		x"41",	--1077
		x"41",	--1078
		x"41",	--1079
		x"41",	--1080
		x"41",	--1081
		x"4b",	--1082
		x"00",	--1083
		x"12",	--1084
		x"cb",	--1085
		x"4f",	--1086
		x"90",	--1087
		x"00",	--1088
		x"3b",	--1089
		x"41",	--1090
		x"4b",	--1091
		x"00",	--1092
		x"12",	--1093
		x"cb",	--1094
		x"4f",	--1095
		x"41",	--1096
		x"4b",	--1097
		x"00",	--1098
		x"12",	--1099
		x"cb",	--1100
		x"4f",	--1101
		x"12",	--1102
		x"12",	--1103
		x"12",	--1104
		x"ed",	--1105
		x"12",	--1106
		x"d2",	--1107
		x"50",	--1108
		x"00",	--1109
		x"4a",	--1110
		x"43",	--1111
		x"12",	--1112
		x"dc",	--1113
		x"43",	--1114
		x"40",	--1115
		x"42",	--1116
		x"12",	--1117
		x"d9",	--1118
		x"4e",	--1119
		x"4f",	--1120
		x"42",	--1121
		x"02",	--1122
		x"12",	--1123
		x"cd",	--1124
		x"4b",	--1125
		x"43",	--1126
		x"12",	--1127
		x"dc",	--1128
		x"43",	--1129
		x"40",	--1130
		x"42",	--1131
		x"12",	--1132
		x"d9",	--1133
		x"4e",	--1134
		x"4f",	--1135
		x"42",	--1136
		x"02",	--1137
		x"12",	--1138
		x"cd",	--1139
		x"3f",	--1140
		x"43",	--1141
		x"12",	--1142
		x"c7",	--1143
		x"43",	--1144
		x"53",	--1145
		x"41",	--1146
		x"41",	--1147
		x"41",	--1148
		x"41",	--1149
		x"41",	--1150
		x"43",	--1151
		x"40",	--1152
		x"c7",	--1153
		x"12",	--1154
		x"cf",	--1155
		x"4f",	--1156
		x"02",	--1157
		x"3f",	--1158
		x"43",	--1159
		x"93",	--1160
		x"02",	--1161
		x"24",	--1162
		x"43",	--1163
		x"4f",	--1164
		x"02",	--1165
		x"43",	--1166
		x"41",	--1167
		x"42",	--1168
		x"00",	--1169
		x"4e",	--1170
		x"be",	--1171
		x"20",	--1172
		x"df",	--1173
		x"00",	--1174
		x"41",	--1175
		x"cf",	--1176
		x"00",	--1177
		x"41",	--1178
		x"42",	--1179
		x"02",	--1180
		x"92",	--1181
		x"2c",	--1182
		x"4e",	--1183
		x"5f",	--1184
		x"4f",	--1185
		x"ed",	--1186
		x"43",	--1187
		x"00",	--1188
		x"90",	--1189
		x"00",	--1190
		x"38",	--1191
		x"43",	--1192
		x"02",	--1193
		x"41",	--1194
		x"53",	--1195
		x"4e",	--1196
		x"02",	--1197
		x"41",	--1198
		x"40",	--1199
		x"00",	--1200
		x"00",	--1201
		x"3f",	--1202
		x"40",	--1203
		x"00",	--1204
		x"00",	--1205
		x"3f",	--1206
		x"42",	--1207
		x"00",	--1208
		x"3f",	--1209
		x"40",	--1210
		x"00",	--1211
		x"00",	--1212
		x"3f",	--1213
		x"40",	--1214
		x"00",	--1215
		x"00",	--1216
		x"3f",	--1217
		x"40",	--1218
		x"00",	--1219
		x"00",	--1220
		x"3f",	--1221
		x"40",	--1222
		x"00",	--1223
		x"00",	--1224
		x"3f",	--1225
		x"4d",	--1226
		x"00",	--1227
		x"4e",	--1228
		x"00",	--1229
		x"41",	--1230
		x"00",	--1231
		x"00",	--1232
		x"41",	--1233
		x"00",	--1234
		x"00",	--1235
		x"41",	--1236
		x"00",	--1237
		x"00",	--1238
		x"41",	--1239
		x"00",	--1240
		x"00",	--1241
		x"43",	--1242
		x"00",	--1243
		x"43",	--1244
		x"00",	--1245
		x"43",	--1246
		x"00",	--1247
		x"43",	--1248
		x"00",	--1249
		x"43",	--1250
		x"00",	--1251
		x"43",	--1252
		x"00",	--1253
		x"41",	--1254
		x"43",	--1255
		x"00",	--1256
		x"43",	--1257
		x"00",	--1258
		x"43",	--1259
		x"00",	--1260
		x"43",	--1261
		x"00",	--1262
		x"43",	--1263
		x"00",	--1264
		x"43",	--1265
		x"00",	--1266
		x"41",	--1267
		x"4d",	--1268
		x"00",	--1269
		x"4e",	--1270
		x"00",	--1271
		x"41",	--1272
		x"4d",	--1273
		x"00",	--1274
		x"4e",	--1275
		x"00",	--1276
		x"41",	--1277
		x"4d",	--1278
		x"00",	--1279
		x"4e",	--1280
		x"00",	--1281
		x"41",	--1282
		x"4d",	--1283
		x"00",	--1284
		x"4e",	--1285
		x"00",	--1286
		x"41",	--1287
		x"12",	--1288
		x"12",	--1289
		x"12",	--1290
		x"12",	--1291
		x"12",	--1292
		x"12",	--1293
		x"12",	--1294
		x"4f",	--1295
		x"4d",	--1296
		x"4e",	--1297
		x"4f",	--1298
		x"00",	--1299
		x"4f",	--1300
		x"00",	--1301
		x"12",	--1302
		x"d7",	--1303
		x"4e",	--1304
		x"4f",	--1305
		x"4b",	--1306
		x"00",	--1307
		x"4b",	--1308
		x"00",	--1309
		x"12",	--1310
		x"d6",	--1311
		x"4e",	--1312
		x"4f",	--1313
		x"4e",	--1314
		x"00",	--1315
		x"4f",	--1316
		x"00",	--1317
		x"4b",	--1318
		x"4b",	--1319
		x"00",	--1320
		x"48",	--1321
		x"49",	--1322
		x"12",	--1323
		x"d7",	--1324
		x"4e",	--1325
		x"4f",	--1326
		x"4b",	--1327
		x"00",	--1328
		x"4b",	--1329
		x"00",	--1330
		x"46",	--1331
		x"47",	--1332
		x"12",	--1333
		x"d7",	--1334
		x"44",	--1335
		x"45",	--1336
		x"12",	--1337
		x"d6",	--1338
		x"4e",	--1339
		x"4f",	--1340
		x"4b",	--1341
		x"00",	--1342
		x"4b",	--1343
		x"00",	--1344
		x"48",	--1345
		x"49",	--1346
		x"12",	--1347
		x"d7",	--1348
		x"4b",	--1349
		x"00",	--1350
		x"4b",	--1351
		x"00",	--1352
		x"12",	--1353
		x"d7",	--1354
		x"46",	--1355
		x"47",	--1356
		x"12",	--1357
		x"d6",	--1358
		x"41",	--1359
		x"41",	--1360
		x"41",	--1361
		x"41",	--1362
		x"41",	--1363
		x"41",	--1364
		x"41",	--1365
		x"41",	--1366
		x"12",	--1367
		x"12",	--1368
		x"83",	--1369
		x"4f",	--1370
		x"4e",	--1371
		x"12",	--1372
		x"ee",	--1373
		x"12",	--1374
		x"d2",	--1375
		x"53",	--1376
		x"90",	--1377
		x"00",	--1378
		x"38",	--1379
		x"41",	--1380
		x"4b",	--1381
		x"00",	--1382
		x"12",	--1383
		x"cb",	--1384
		x"4f",	--1385
		x"41",	--1386
		x"4b",	--1387
		x"00",	--1388
		x"12",	--1389
		x"cb",	--1390
		x"4f",	--1391
		x"12",	--1392
		x"12",	--1393
		x"12",	--1394
		x"ee",	--1395
		x"12",	--1396
		x"d2",	--1397
		x"50",	--1398
		x"00",	--1399
		x"4b",	--1400
		x"00",	--1401
		x"43",	--1402
		x"53",	--1403
		x"41",	--1404
		x"41",	--1405
		x"41",	--1406
		x"12",	--1407
		x"ee",	--1408
		x"12",	--1409
		x"d2",	--1410
		x"40",	--1411
		x"ee",	--1412
		x"00",	--1413
		x"12",	--1414
		x"d2",	--1415
		x"4b",	--1416
		x"00",	--1417
		x"12",	--1418
		x"ee",	--1419
		x"12",	--1420
		x"d2",	--1421
		x"52",	--1422
		x"43",	--1423
		x"3f",	--1424
		x"12",	--1425
		x"83",	--1426
		x"4e",	--1427
		x"93",	--1428
		x"24",	--1429
		x"38",	--1430
		x"12",	--1431
		x"ee",	--1432
		x"12",	--1433
		x"d2",	--1434
		x"53",	--1435
		x"41",	--1436
		x"4b",	--1437
		x"00",	--1438
		x"12",	--1439
		x"cb",	--1440
		x"12",	--1441
		x"12",	--1442
		x"12",	--1443
		x"ee",	--1444
		x"12",	--1445
		x"d2",	--1446
		x"50",	--1447
		x"00",	--1448
		x"43",	--1449
		x"53",	--1450
		x"41",	--1451
		x"41",	--1452
		x"12",	--1453
		x"ee",	--1454
		x"12",	--1455
		x"d2",	--1456
		x"40",	--1457
		x"ee",	--1458
		x"00",	--1459
		x"12",	--1460
		x"d2",	--1461
		x"4b",	--1462
		x"00",	--1463
		x"12",	--1464
		x"ee",	--1465
		x"12",	--1466
		x"d2",	--1467
		x"52",	--1468
		x"43",	--1469
		x"3f",	--1470
		x"12",	--1471
		x"12",	--1472
		x"43",	--1473
		x"00",	--1474
		x"4f",	--1475
		x"93",	--1476
		x"24",	--1477
		x"53",	--1478
		x"43",	--1479
		x"43",	--1480
		x"3c",	--1481
		x"90",	--1482
		x"00",	--1483
		x"2c",	--1484
		x"5c",	--1485
		x"5c",	--1486
		x"5c",	--1487
		x"5c",	--1488
		x"11",	--1489
		x"5d",	--1490
		x"50",	--1491
		x"ff",	--1492
		x"43",	--1493
		x"4f",	--1494
		x"93",	--1495
		x"24",	--1496
		x"90",	--1497
		x"00",	--1498
		x"24",	--1499
		x"4d",	--1500
		x"50",	--1501
		x"ff",	--1502
		x"93",	--1503
		x"23",	--1504
		x"90",	--1505
		x"00",	--1506
		x"2c",	--1507
		x"5c",	--1508
		x"4c",	--1509
		x"5b",	--1510
		x"5b",	--1511
		x"5b",	--1512
		x"11",	--1513
		x"5d",	--1514
		x"50",	--1515
		x"ff",	--1516
		x"4f",	--1517
		x"93",	--1518
		x"23",	--1519
		x"43",	--1520
		x"00",	--1521
		x"4c",	--1522
		x"41",	--1523
		x"41",	--1524
		x"41",	--1525
		x"43",	--1526
		x"3f",	--1527
		x"4d",	--1528
		x"50",	--1529
		x"ff",	--1530
		x"90",	--1531
		x"00",	--1532
		x"2c",	--1533
		x"5c",	--1534
		x"5c",	--1535
		x"5c",	--1536
		x"5c",	--1537
		x"11",	--1538
		x"5d",	--1539
		x"50",	--1540
		x"ff",	--1541
		x"43",	--1542
		x"3f",	--1543
		x"4d",	--1544
		x"50",	--1545
		x"ff",	--1546
		x"90",	--1547
		x"00",	--1548
		x"2c",	--1549
		x"5c",	--1550
		x"5c",	--1551
		x"5c",	--1552
		x"5c",	--1553
		x"11",	--1554
		x"5d",	--1555
		x"50",	--1556
		x"ff",	--1557
		x"43",	--1558
		x"3f",	--1559
		x"11",	--1560
		x"12",	--1561
		x"12",	--1562
		x"ee",	--1563
		x"12",	--1564
		x"d2",	--1565
		x"52",	--1566
		x"43",	--1567
		x"4c",	--1568
		x"41",	--1569
		x"41",	--1570
		x"41",	--1571
		x"43",	--1572
		x"3f",	--1573
		x"12",	--1574
		x"12",	--1575
		x"43",	--1576
		x"00",	--1577
		x"4f",	--1578
		x"93",	--1579
		x"24",	--1580
		x"53",	--1581
		x"43",	--1582
		x"43",	--1583
		x"3c",	--1584
		x"4b",	--1585
		x"50",	--1586
		x"ff",	--1587
		x"90",	--1588
		x"00",	--1589
		x"2c",	--1590
		x"5c",	--1591
		x"4c",	--1592
		x"5d",	--1593
		x"5d",	--1594
		x"5d",	--1595
		x"11",	--1596
		x"5b",	--1597
		x"50",	--1598
		x"ff",	--1599
		x"4f",	--1600
		x"93",	--1601
		x"24",	--1602
		x"90",	--1603
		x"00",	--1604
		x"23",	--1605
		x"43",	--1606
		x"4f",	--1607
		x"93",	--1608
		x"23",	--1609
		x"12",	--1610
		x"c2",	--1611
		x"43",	--1612
		x"4a",	--1613
		x"01",	--1614
		x"4c",	--1615
		x"01",	--1616
		x"42",	--1617
		x"01",	--1618
		x"41",	--1619
		x"43",	--1620
		x"00",	--1621
		x"41",	--1622
		x"41",	--1623
		x"41",	--1624
		x"11",	--1625
		x"12",	--1626
		x"12",	--1627
		x"ee",	--1628
		x"12",	--1629
		x"d2",	--1630
		x"52",	--1631
		x"43",	--1632
		x"41",	--1633
		x"41",	--1634
		x"41",	--1635
		x"43",	--1636
		x"3f",	--1637
		x"12",	--1638
		x"12",	--1639
		x"4e",	--1640
		x"4c",	--1641
		x"4e",	--1642
		x"00",	--1643
		x"4d",	--1644
		x"00",	--1645
		x"4c",	--1646
		x"00",	--1647
		x"4d",	--1648
		x"43",	--1649
		x"40",	--1650
		x"36",	--1651
		x"40",	--1652
		x"01",	--1653
		x"12",	--1654
		x"eb",	--1655
		x"4e",	--1656
		x"00",	--1657
		x"12",	--1658
		x"c2",	--1659
		x"43",	--1660
		x"4a",	--1661
		x"01",	--1662
		x"40",	--1663
		x"00",	--1664
		x"01",	--1665
		x"42",	--1666
		x"01",	--1667
		x"00",	--1668
		x"41",	--1669
		x"43",	--1670
		x"41",	--1671
		x"41",	--1672
		x"41",	--1673
		x"12",	--1674
		x"12",	--1675
		x"12",	--1676
		x"43",	--1677
		x"00",	--1678
		x"40",	--1679
		x"3f",	--1680
		x"00",	--1681
		x"4f",	--1682
		x"4b",	--1683
		x"00",	--1684
		x"43",	--1685
		x"12",	--1686
		x"dc",	--1687
		x"43",	--1688
		x"40",	--1689
		x"3f",	--1690
		x"12",	--1691
		x"d7",	--1692
		x"4e",	--1693
		x"4f",	--1694
		x"4b",	--1695
		x"00",	--1696
		x"43",	--1697
		x"12",	--1698
		x"dc",	--1699
		x"4e",	--1700
		x"4f",	--1701
		x"48",	--1702
		x"49",	--1703
		x"12",	--1704
		x"d7",	--1705
		x"12",	--1706
		x"d3",	--1707
		x"4e",	--1708
		x"00",	--1709
		x"43",	--1710
		x"00",	--1711
		x"41",	--1712
		x"41",	--1713
		x"41",	--1714
		x"41",	--1715
		x"12",	--1716
		x"12",	--1717
		x"12",	--1718
		x"4d",	--1719
		x"4e",	--1720
		x"4d",	--1721
		x"00",	--1722
		x"4e",	--1723
		x"00",	--1724
		x"4f",	--1725
		x"49",	--1726
		x"00",	--1727
		x"43",	--1728
		x"12",	--1729
		x"dc",	--1730
		x"4e",	--1731
		x"4f",	--1732
		x"4a",	--1733
		x"4b",	--1734
		x"12",	--1735
		x"d7",	--1736
		x"4e",	--1737
		x"4f",	--1738
		x"49",	--1739
		x"00",	--1740
		x"43",	--1741
		x"12",	--1742
		x"dc",	--1743
		x"4e",	--1744
		x"4f",	--1745
		x"4a",	--1746
		x"4b",	--1747
		x"12",	--1748
		x"d7",	--1749
		x"12",	--1750
		x"d3",	--1751
		x"4e",	--1752
		x"00",	--1753
		x"41",	--1754
		x"41",	--1755
		x"41",	--1756
		x"41",	--1757
		x"4f",	--1758
		x"4e",	--1759
		x"00",	--1760
		x"41",	--1761
		x"12",	--1762
		x"12",	--1763
		x"93",	--1764
		x"02",	--1765
		x"38",	--1766
		x"40",	--1767
		x"02",	--1768
		x"43",	--1769
		x"12",	--1770
		x"4b",	--1771
		x"ff",	--1772
		x"11",	--1773
		x"12",	--1774
		x"12",	--1775
		x"ee",	--1776
		x"12",	--1777
		x"d2",	--1778
		x"50",	--1779
		x"00",	--1780
		x"53",	--1781
		x"50",	--1782
		x"00",	--1783
		x"92",	--1784
		x"02",	--1785
		x"3b",	--1786
		x"43",	--1787
		x"41",	--1788
		x"41",	--1789
		x"41",	--1790
		x"42",	--1791
		x"02",	--1792
		x"90",	--1793
		x"00",	--1794
		x"34",	--1795
		x"4e",	--1796
		x"5f",	--1797
		x"5e",	--1798
		x"5f",	--1799
		x"50",	--1800
		x"02",	--1801
		x"40",	--1802
		x"00",	--1803
		x"00",	--1804
		x"40",	--1805
		x"cd",	--1806
		x"00",	--1807
		x"40",	--1808
		x"02",	--1809
		x"00",	--1810
		x"53",	--1811
		x"4e",	--1812
		x"02",	--1813
		x"41",	--1814
		x"12",	--1815
		x"42",	--1816
		x"02",	--1817
		x"90",	--1818
		x"00",	--1819
		x"34",	--1820
		x"4b",	--1821
		x"5c",	--1822
		x"5b",	--1823
		x"5c",	--1824
		x"50",	--1825
		x"02",	--1826
		x"4f",	--1827
		x"00",	--1828
		x"4e",	--1829
		x"00",	--1830
		x"4d",	--1831
		x"00",	--1832
		x"53",	--1833
		x"4b",	--1834
		x"02",	--1835
		x"43",	--1836
		x"41",	--1837
		x"41",	--1838
		x"43",	--1839
		x"3f",	--1840
		x"12",	--1841
		x"50",	--1842
		x"ff",	--1843
		x"42",	--1844
		x"02",	--1845
		x"93",	--1846
		x"38",	--1847
		x"92",	--1848
		x"02",	--1849
		x"24",	--1850
		x"40",	--1851
		x"02",	--1852
		x"43",	--1853
		x"3c",	--1854
		x"50",	--1855
		x"00",	--1856
		x"9f",	--1857
		x"ff",	--1858
		x"24",	--1859
		x"53",	--1860
		x"9b",	--1861
		x"23",	--1862
		x"12",	--1863
		x"ee",	--1864
		x"12",	--1865
		x"d2",	--1866
		x"53",	--1867
		x"43",	--1868
		x"50",	--1869
		x"00",	--1870
		x"41",	--1871
		x"41",	--1872
		x"43",	--1873
		x"4e",	--1874
		x"00",	--1875
		x"4e",	--1876
		x"93",	--1877
		x"24",	--1878
		x"53",	--1879
		x"43",	--1880
		x"3c",	--1881
		x"4e",	--1882
		x"93",	--1883
		x"24",	--1884
		x"53",	--1885
		x"92",	--1886
		x"34",	--1887
		x"90",	--1888
		x"00",	--1889
		x"23",	--1890
		x"43",	--1891
		x"ff",	--1892
		x"4f",	--1893
		x"5d",	--1894
		x"51",	--1895
		x"4e",	--1896
		x"00",	--1897
		x"53",	--1898
		x"4e",	--1899
		x"93",	--1900
		x"23",	--1901
		x"4c",	--1902
		x"5e",	--1903
		x"5e",	--1904
		x"5c",	--1905
		x"50",	--1906
		x"02",	--1907
		x"41",	--1908
		x"12",	--1909
		x"00",	--1910
		x"50",	--1911
		x"00",	--1912
		x"41",	--1913
		x"41",	--1914
		x"43",	--1915
		x"3f",	--1916
		x"d0",	--1917
		x"02",	--1918
		x"01",	--1919
		x"40",	--1920
		x"0b",	--1921
		x"01",	--1922
		x"43",	--1923
		x"41",	--1924
		x"12",	--1925
		x"4f",	--1926
		x"42",	--1927
		x"02",	--1928
		x"90",	--1929
		x"00",	--1930
		x"34",	--1931
		x"4f",	--1932
		x"5c",	--1933
		x"4c",	--1934
		x"5d",	--1935
		x"5d",	--1936
		x"5d",	--1937
		x"8c",	--1938
		x"50",	--1939
		x"03",	--1940
		x"43",	--1941
		x"00",	--1942
		x"43",	--1943
		x"00",	--1944
		x"43",	--1945
		x"00",	--1946
		x"4b",	--1947
		x"00",	--1948
		x"4e",	--1949
		x"00",	--1950
		x"4f",	--1951
		x"53",	--1952
		x"4e",	--1953
		x"02",	--1954
		x"41",	--1955
		x"41",	--1956
		x"43",	--1957
		x"3f",	--1958
		x"5f",	--1959
		x"4f",	--1960
		x"5c",	--1961
		x"5c",	--1962
		x"5c",	--1963
		x"8f",	--1964
		x"50",	--1965
		x"03",	--1966
		x"43",	--1967
		x"00",	--1968
		x"4e",	--1969
		x"00",	--1970
		x"43",	--1971
		x"00",	--1972
		x"4d",	--1973
		x"00",	--1974
		x"43",	--1975
		x"00",	--1976
		x"43",	--1977
		x"41",	--1978
		x"5f",	--1979
		x"4f",	--1980
		x"5e",	--1981
		x"5e",	--1982
		x"5e",	--1983
		x"8f",	--1984
		x"43",	--1985
		x"03",	--1986
		x"43",	--1987
		x"41",	--1988
		x"12",	--1989
		x"12",	--1990
		x"12",	--1991
		x"12",	--1992
		x"12",	--1993
		x"12",	--1994
		x"12",	--1995
		x"12",	--1996
		x"12",	--1997
		x"93",	--1998
		x"02",	--1999
		x"38",	--2000
		x"40",	--2001
		x"03",	--2002
		x"4a",	--2003
		x"53",	--2004
		x"4a",	--2005
		x"52",	--2006
		x"4a",	--2007
		x"50",	--2008
		x"00",	--2009
		x"43",	--2010
		x"3c",	--2011
		x"53",	--2012
		x"4f",	--2013
		x"00",	--2014
		x"53",	--2015
		x"50",	--2016
		x"00",	--2017
		x"50",	--2018
		x"00",	--2019
		x"50",	--2020
		x"00",	--2021
		x"50",	--2022
		x"00",	--2023
		x"92",	--2024
		x"02",	--2025
		x"34",	--2026
		x"93",	--2027
		x"00",	--2028
		x"27",	--2029
		x"4b",	--2030
		x"9b",	--2031
		x"00",	--2032
		x"2b",	--2033
		x"43",	--2034
		x"00",	--2035
		x"4b",	--2036
		x"00",	--2037
		x"12",	--2038
		x"00",	--2039
		x"93",	--2040
		x"00",	--2041
		x"27",	--2042
		x"47",	--2043
		x"53",	--2044
		x"4f",	--2045
		x"00",	--2046
		x"98",	--2047
		x"2b",	--2048
		x"43",	--2049
		x"00",	--2050
		x"3f",	--2051
		x"f0",	--2052
		x"ff",	--2053
		x"01",	--2054
		x"41",	--2055
		x"41",	--2056
		x"41",	--2057
		x"41",	--2058
		x"41",	--2059
		x"41",	--2060
		x"41",	--2061
		x"41",	--2062
		x"41",	--2063
		x"13",	--2064
		x"4e",	--2065
		x"00",	--2066
		x"43",	--2067
		x"41",	--2068
		x"4f",	--2069
		x"4f",	--2070
		x"4f",	--2071
		x"00",	--2072
		x"41",	--2073
		x"43",	--2074
		x"00",	--2075
		x"41",	--2076
		x"4e",	--2077
		x"00",	--2078
		x"40",	--2079
		x"d0",	--2080
		x"12",	--2081
		x"cf",	--2082
		x"4f",	--2083
		x"02",	--2084
		x"43",	--2085
		x"41",	--2086
		x"4d",	--2087
		x"4f",	--2088
		x"4e",	--2089
		x"00",	--2090
		x"43",	--2091
		x"4c",	--2092
		x"42",	--2093
		x"02",	--2094
		x"12",	--2095
		x"cf",	--2096
		x"41",	--2097
		x"42",	--2098
		x"00",	--2099
		x"f2",	--2100
		x"23",	--2101
		x"4f",	--2102
		x"00",	--2103
		x"43",	--2104
		x"41",	--2105
		x"f0",	--2106
		x"00",	--2107
		x"4f",	--2108
		x"ef",	--2109
		x"11",	--2110
		x"12",	--2111
		x"d0",	--2112
		x"41",	--2113
		x"12",	--2114
		x"4f",	--2115
		x"4f",	--2116
		x"11",	--2117
		x"11",	--2118
		x"11",	--2119
		x"11",	--2120
		x"4e",	--2121
		x"12",	--2122
		x"d0",	--2123
		x"4b",	--2124
		x"12",	--2125
		x"d0",	--2126
		x"41",	--2127
		x"41",	--2128
		x"12",	--2129
		x"12",	--2130
		x"4f",	--2131
		x"40",	--2132
		x"00",	--2133
		x"4a",	--2134
		x"4b",	--2135
		x"f0",	--2136
		x"00",	--2137
		x"24",	--2138
		x"11",	--2139
		x"53",	--2140
		x"23",	--2141
		x"f3",	--2142
		x"24",	--2143
		x"40",	--2144
		x"00",	--2145
		x"12",	--2146
		x"d0",	--2147
		x"53",	--2148
		x"93",	--2149
		x"23",	--2150
		x"41",	--2151
		x"41",	--2152
		x"41",	--2153
		x"40",	--2154
		x"00",	--2155
		x"3f",	--2156
		x"12",	--2157
		x"4f",	--2158
		x"4f",	--2159
		x"10",	--2160
		x"11",	--2161
		x"4e",	--2162
		x"12",	--2163
		x"d0",	--2164
		x"4b",	--2165
		x"12",	--2166
		x"d0",	--2167
		x"41",	--2168
		x"41",	--2169
		x"12",	--2170
		x"12",	--2171
		x"4e",	--2172
		x"4f",	--2173
		x"4f",	--2174
		x"10",	--2175
		x"11",	--2176
		x"4d",	--2177
		x"12",	--2178
		x"d0",	--2179
		x"4b",	--2180
		x"12",	--2181
		x"d0",	--2182
		x"4b",	--2183
		x"4a",	--2184
		x"10",	--2185
		x"10",	--2186
		x"ec",	--2187
		x"ec",	--2188
		x"4d",	--2189
		x"12",	--2190
		x"d0",	--2191
		x"4a",	--2192
		x"12",	--2193
		x"d0",	--2194
		x"41",	--2195
		x"41",	--2196
		x"41",	--2197
		x"12",	--2198
		x"12",	--2199
		x"12",	--2200
		x"4f",	--2201
		x"93",	--2202
		x"24",	--2203
		x"4e",	--2204
		x"53",	--2205
		x"43",	--2206
		x"4a",	--2207
		x"5b",	--2208
		x"4d",	--2209
		x"11",	--2210
		x"12",	--2211
		x"d0",	--2212
		x"99",	--2213
		x"24",	--2214
		x"53",	--2215
		x"b0",	--2216
		x"00",	--2217
		x"20",	--2218
		x"40",	--2219
		x"00",	--2220
		x"12",	--2221
		x"d0",	--2222
		x"3f",	--2223
		x"40",	--2224
		x"00",	--2225
		x"12",	--2226
		x"d0",	--2227
		x"3f",	--2228
		x"41",	--2229
		x"41",	--2230
		x"41",	--2231
		x"41",	--2232
		x"12",	--2233
		x"12",	--2234
		x"12",	--2235
		x"4f",	--2236
		x"93",	--2237
		x"24",	--2238
		x"4e",	--2239
		x"53",	--2240
		x"43",	--2241
		x"4a",	--2242
		x"11",	--2243
		x"12",	--2244
		x"d0",	--2245
		x"99",	--2246
		x"24",	--2247
		x"53",	--2248
		x"b0",	--2249
		x"00",	--2250
		x"23",	--2251
		x"40",	--2252
		x"00",	--2253
		x"12",	--2254
		x"d0",	--2255
		x"4a",	--2256
		x"11",	--2257
		x"12",	--2258
		x"d0",	--2259
		x"99",	--2260
		x"23",	--2261
		x"41",	--2262
		x"41",	--2263
		x"41",	--2264
		x"41",	--2265
		x"12",	--2266
		x"12",	--2267
		x"12",	--2268
		x"50",	--2269
		x"ff",	--2270
		x"4f",	--2271
		x"93",	--2272
		x"38",	--2273
		x"90",	--2274
		x"00",	--2275
		x"38",	--2276
		x"43",	--2277
		x"41",	--2278
		x"59",	--2279
		x"40",	--2280
		x"00",	--2281
		x"4b",	--2282
		x"12",	--2283
		x"eb",	--2284
		x"50",	--2285
		x"00",	--2286
		x"4f",	--2287
		x"00",	--2288
		x"53",	--2289
		x"40",	--2290
		x"00",	--2291
		x"4b",	--2292
		x"12",	--2293
		x"ea",	--2294
		x"4f",	--2295
		x"90",	--2296
		x"00",	--2297
		x"37",	--2298
		x"49",	--2299
		x"53",	--2300
		x"51",	--2301
		x"40",	--2302
		x"00",	--2303
		x"4b",	--2304
		x"12",	--2305
		x"eb",	--2306
		x"50",	--2307
		x"00",	--2308
		x"4f",	--2309
		x"00",	--2310
		x"53",	--2311
		x"41",	--2312
		x"5a",	--2313
		x"4f",	--2314
		x"11",	--2315
		x"12",	--2316
		x"d0",	--2317
		x"93",	--2318
		x"23",	--2319
		x"50",	--2320
		x"00",	--2321
		x"41",	--2322
		x"41",	--2323
		x"41",	--2324
		x"41",	--2325
		x"40",	--2326
		x"00",	--2327
		x"12",	--2328
		x"d0",	--2329
		x"e3",	--2330
		x"53",	--2331
		x"3f",	--2332
		x"43",	--2333
		x"43",	--2334
		x"3f",	--2335
		x"12",	--2336
		x"12",	--2337
		x"12",	--2338
		x"41",	--2339
		x"52",	--2340
		x"4b",	--2341
		x"49",	--2342
		x"93",	--2343
		x"20",	--2344
		x"3c",	--2345
		x"11",	--2346
		x"12",	--2347
		x"d0",	--2348
		x"49",	--2349
		x"4a",	--2350
		x"53",	--2351
		x"4a",	--2352
		x"00",	--2353
		x"93",	--2354
		x"24",	--2355
		x"90",	--2356
		x"00",	--2357
		x"23",	--2358
		x"49",	--2359
		x"53",	--2360
		x"49",	--2361
		x"00",	--2362
		x"50",	--2363
		x"ff",	--2364
		x"90",	--2365
		x"00",	--2366
		x"2f",	--2367
		x"4f",	--2368
		x"5f",	--2369
		x"4f",	--2370
		x"ef",	--2371
		x"41",	--2372
		x"41",	--2373
		x"41",	--2374
		x"41",	--2375
		x"4b",	--2376
		x"52",	--2377
		x"4b",	--2378
		x"00",	--2379
		x"4b",	--2380
		x"12",	--2381
		x"d1",	--2382
		x"49",	--2383
		x"3f",	--2384
		x"4b",	--2385
		x"53",	--2386
		x"4b",	--2387
		x"12",	--2388
		x"d0",	--2389
		x"49",	--2390
		x"3f",	--2391
		x"4b",	--2392
		x"53",	--2393
		x"4f",	--2394
		x"49",	--2395
		x"93",	--2396
		x"27",	--2397
		x"53",	--2398
		x"11",	--2399
		x"12",	--2400
		x"d0",	--2401
		x"49",	--2402
		x"93",	--2403
		x"23",	--2404
		x"3f",	--2405
		x"4b",	--2406
		x"52",	--2407
		x"4b",	--2408
		x"00",	--2409
		x"4b",	--2410
		x"12",	--2411
		x"d1",	--2412
		x"49",	--2413
		x"3f",	--2414
		x"4b",	--2415
		x"53",	--2416
		x"4b",	--2417
		x"4e",	--2418
		x"10",	--2419
		x"11",	--2420
		x"10",	--2421
		x"11",	--2422
		x"12",	--2423
		x"d0",	--2424
		x"49",	--2425
		x"3f",	--2426
		x"4b",	--2427
		x"53",	--2428
		x"4b",	--2429
		x"12",	--2430
		x"d1",	--2431
		x"49",	--2432
		x"3f",	--2433
		x"4b",	--2434
		x"53",	--2435
		x"4b",	--2436
		x"12",	--2437
		x"d0",	--2438
		x"49",	--2439
		x"3f",	--2440
		x"4b",	--2441
		x"53",	--2442
		x"4b",	--2443
		x"12",	--2444
		x"d0",	--2445
		x"49",	--2446
		x"3f",	--2447
		x"4b",	--2448
		x"53",	--2449
		x"4b",	--2450
		x"12",	--2451
		x"d0",	--2452
		x"49",	--2453
		x"3f",	--2454
		x"40",	--2455
		x"00",	--2456
		x"12",	--2457
		x"d0",	--2458
		x"3f",	--2459
		x"12",	--2460
		x"12",	--2461
		x"42",	--2462
		x"02",	--2463
		x"42",	--2464
		x"00",	--2465
		x"04",	--2466
		x"42",	--2467
		x"02",	--2468
		x"90",	--2469
		x"00",	--2470
		x"34",	--2471
		x"53",	--2472
		x"02",	--2473
		x"42",	--2474
		x"02",	--2475
		x"42",	--2476
		x"02",	--2477
		x"9f",	--2478
		x"20",	--2479
		x"53",	--2480
		x"02",	--2481
		x"40",	--2482
		x"00",	--2483
		x"00",	--2484
		x"41",	--2485
		x"41",	--2486
		x"c0",	--2487
		x"00",	--2488
		x"00",	--2489
		x"13",	--2490
		x"43",	--2491
		x"02",	--2492
		x"3f",	--2493
		x"4e",	--2494
		x"4f",	--2495
		x"40",	--2496
		x"36",	--2497
		x"40",	--2498
		x"01",	--2499
		x"12",	--2500
		x"eb",	--2501
		x"53",	--2502
		x"4e",	--2503
		x"00",	--2504
		x"40",	--2505
		x"00",	--2506
		x"00",	--2507
		x"41",	--2508
		x"42",	--2509
		x"02",	--2510
		x"42",	--2511
		x"02",	--2512
		x"9f",	--2513
		x"38",	--2514
		x"42",	--2515
		x"02",	--2516
		x"82",	--2517
		x"02",	--2518
		x"41",	--2519
		x"42",	--2520
		x"02",	--2521
		x"42",	--2522
		x"02",	--2523
		x"40",	--2524
		x"00",	--2525
		x"8d",	--2526
		x"8e",	--2527
		x"41",	--2528
		x"42",	--2529
		x"02",	--2530
		x"4f",	--2531
		x"04",	--2532
		x"42",	--2533
		x"02",	--2534
		x"42",	--2535
		x"02",	--2536
		x"9e",	--2537
		x"24",	--2538
		x"42",	--2539
		x"02",	--2540
		x"90",	--2541
		x"00",	--2542
		x"38",	--2543
		x"43",	--2544
		x"02",	--2545
		x"41",	--2546
		x"53",	--2547
		x"02",	--2548
		x"41",	--2549
		x"43",	--2550
		x"41",	--2551
		x"12",	--2552
		x"12",	--2553
		x"4e",	--2554
		x"4f",	--2555
		x"43",	--2556
		x"40",	--2557
		x"4f",	--2558
		x"12",	--2559
		x"db",	--2560
		x"93",	--2561
		x"34",	--2562
		x"4a",	--2563
		x"4b",	--2564
		x"12",	--2565
		x"dc",	--2566
		x"41",	--2567
		x"41",	--2568
		x"41",	--2569
		x"43",	--2570
		x"40",	--2571
		x"4f",	--2572
		x"4a",	--2573
		x"4b",	--2574
		x"12",	--2575
		x"d7",	--2576
		x"12",	--2577
		x"dc",	--2578
		x"53",	--2579
		x"60",	--2580
		x"80",	--2581
		x"41",	--2582
		x"41",	--2583
		x"41",	--2584
		x"12",	--2585
		x"12",	--2586
		x"12",	--2587
		x"12",	--2588
		x"12",	--2589
		x"12",	--2590
		x"12",	--2591
		x"12",	--2592
		x"50",	--2593
		x"ff",	--2594
		x"4d",	--2595
		x"4f",	--2596
		x"93",	--2597
		x"28",	--2598
		x"4e",	--2599
		x"93",	--2600
		x"28",	--2601
		x"92",	--2602
		x"20",	--2603
		x"40",	--2604
		x"d6",	--2605
		x"92",	--2606
		x"24",	--2607
		x"93",	--2608
		x"24",	--2609
		x"93",	--2610
		x"24",	--2611
		x"4f",	--2612
		x"00",	--2613
		x"00",	--2614
		x"4e",	--2615
		x"00",	--2616
		x"4f",	--2617
		x"00",	--2618
		x"4f",	--2619
		x"00",	--2620
		x"4e",	--2621
		x"00",	--2622
		x"4e",	--2623
		x"00",	--2624
		x"41",	--2625
		x"8b",	--2626
		x"4c",	--2627
		x"93",	--2628
		x"38",	--2629
		x"90",	--2630
		x"00",	--2631
		x"34",	--2632
		x"93",	--2633
		x"38",	--2634
		x"46",	--2635
		x"00",	--2636
		x"47",	--2637
		x"00",	--2638
		x"49",	--2639
		x"f0",	--2640
		x"00",	--2641
		x"24",	--2642
		x"46",	--2643
		x"47",	--2644
		x"c3",	--2645
		x"10",	--2646
		x"10",	--2647
		x"53",	--2648
		x"23",	--2649
		x"4a",	--2650
		x"00",	--2651
		x"4b",	--2652
		x"00",	--2653
		x"43",	--2654
		x"43",	--2655
		x"f0",	--2656
		x"00",	--2657
		x"24",	--2658
		x"5c",	--2659
		x"6d",	--2660
		x"53",	--2661
		x"23",	--2662
		x"53",	--2663
		x"63",	--2664
		x"f6",	--2665
		x"f7",	--2666
		x"43",	--2667
		x"43",	--2668
		x"93",	--2669
		x"20",	--2670
		x"93",	--2671
		x"24",	--2672
		x"41",	--2673
		x"00",	--2674
		x"41",	--2675
		x"00",	--2676
		x"da",	--2677
		x"db",	--2678
		x"4f",	--2679
		x"00",	--2680
		x"9e",	--2681
		x"00",	--2682
		x"20",	--2683
		x"4f",	--2684
		x"00",	--2685
		x"41",	--2686
		x"00",	--2687
		x"46",	--2688
		x"47",	--2689
		x"54",	--2690
		x"65",	--2691
		x"4e",	--2692
		x"00",	--2693
		x"4f",	--2694
		x"00",	--2695
		x"40",	--2696
		x"00",	--2697
		x"00",	--2698
		x"93",	--2699
		x"38",	--2700
		x"48",	--2701
		x"50",	--2702
		x"00",	--2703
		x"41",	--2704
		x"41",	--2705
		x"41",	--2706
		x"41",	--2707
		x"41",	--2708
		x"41",	--2709
		x"41",	--2710
		x"41",	--2711
		x"41",	--2712
		x"91",	--2713
		x"38",	--2714
		x"4b",	--2715
		x"00",	--2716
		x"43",	--2717
		x"43",	--2718
		x"4f",	--2719
		x"00",	--2720
		x"9e",	--2721
		x"00",	--2722
		x"27",	--2723
		x"93",	--2724
		x"24",	--2725
		x"46",	--2726
		x"47",	--2727
		x"84",	--2728
		x"75",	--2729
		x"93",	--2730
		x"38",	--2731
		x"43",	--2732
		x"00",	--2733
		x"41",	--2734
		x"00",	--2735
		x"4e",	--2736
		x"00",	--2737
		x"4f",	--2738
		x"00",	--2739
		x"4e",	--2740
		x"4f",	--2741
		x"53",	--2742
		x"63",	--2743
		x"90",	--2744
		x"3f",	--2745
		x"28",	--2746
		x"90",	--2747
		x"40",	--2748
		x"2c",	--2749
		x"93",	--2750
		x"2c",	--2751
		x"48",	--2752
		x"00",	--2753
		x"53",	--2754
		x"5e",	--2755
		x"6f",	--2756
		x"4b",	--2757
		x"53",	--2758
		x"4e",	--2759
		x"4f",	--2760
		x"53",	--2761
		x"63",	--2762
		x"90",	--2763
		x"3f",	--2764
		x"2b",	--2765
		x"24",	--2766
		x"4e",	--2767
		x"00",	--2768
		x"4f",	--2769
		x"00",	--2770
		x"4a",	--2771
		x"00",	--2772
		x"40",	--2773
		x"00",	--2774
		x"00",	--2775
		x"93",	--2776
		x"37",	--2777
		x"4e",	--2778
		x"4f",	--2779
		x"f3",	--2780
		x"f3",	--2781
		x"c3",	--2782
		x"10",	--2783
		x"10",	--2784
		x"4c",	--2785
		x"4d",	--2786
		x"de",	--2787
		x"df",	--2788
		x"4a",	--2789
		x"00",	--2790
		x"4b",	--2791
		x"00",	--2792
		x"53",	--2793
		x"00",	--2794
		x"48",	--2795
		x"3f",	--2796
		x"93",	--2797
		x"23",	--2798
		x"4f",	--2799
		x"00",	--2800
		x"4f",	--2801
		x"00",	--2802
		x"00",	--2803
		x"4f",	--2804
		x"00",	--2805
		x"00",	--2806
		x"4f",	--2807
		x"00",	--2808
		x"00",	--2809
		x"4e",	--2810
		x"00",	--2811
		x"ff",	--2812
		x"00",	--2813
		x"4e",	--2814
		x"00",	--2815
		x"4d",	--2816
		x"3f",	--2817
		x"43",	--2818
		x"43",	--2819
		x"3f",	--2820
		x"e3",	--2821
		x"53",	--2822
		x"90",	--2823
		x"00",	--2824
		x"37",	--2825
		x"3f",	--2826
		x"93",	--2827
		x"2b",	--2828
		x"3f",	--2829
		x"44",	--2830
		x"45",	--2831
		x"86",	--2832
		x"77",	--2833
		x"3f",	--2834
		x"4e",	--2835
		x"3f",	--2836
		x"43",	--2837
		x"00",	--2838
		x"41",	--2839
		x"00",	--2840
		x"e3",	--2841
		x"e3",	--2842
		x"53",	--2843
		x"63",	--2844
		x"4e",	--2845
		x"00",	--2846
		x"4f",	--2847
		x"00",	--2848
		x"3f",	--2849
		x"93",	--2850
		x"27",	--2851
		x"59",	--2852
		x"00",	--2853
		x"44",	--2854
		x"00",	--2855
		x"45",	--2856
		x"00",	--2857
		x"49",	--2858
		x"f0",	--2859
		x"00",	--2860
		x"24",	--2861
		x"4d",	--2862
		x"44",	--2863
		x"45",	--2864
		x"c3",	--2865
		x"10",	--2866
		x"10",	--2867
		x"53",	--2868
		x"23",	--2869
		x"4c",	--2870
		x"00",	--2871
		x"4d",	--2872
		x"00",	--2873
		x"43",	--2874
		x"43",	--2875
		x"f0",	--2876
		x"00",	--2877
		x"24",	--2878
		x"5c",	--2879
		x"6d",	--2880
		x"53",	--2881
		x"23",	--2882
		x"53",	--2883
		x"63",	--2884
		x"f4",	--2885
		x"f5",	--2886
		x"43",	--2887
		x"43",	--2888
		x"93",	--2889
		x"20",	--2890
		x"93",	--2891
		x"20",	--2892
		x"43",	--2893
		x"43",	--2894
		x"41",	--2895
		x"00",	--2896
		x"41",	--2897
		x"00",	--2898
		x"da",	--2899
		x"db",	--2900
		x"3f",	--2901
		x"43",	--2902
		x"43",	--2903
		x"3f",	--2904
		x"92",	--2905
		x"23",	--2906
		x"9e",	--2907
		x"00",	--2908
		x"00",	--2909
		x"27",	--2910
		x"40",	--2911
		x"ef",	--2912
		x"3f",	--2913
		x"50",	--2914
		x"ff",	--2915
		x"4e",	--2916
		x"00",	--2917
		x"4f",	--2918
		x"00",	--2919
		x"4c",	--2920
		x"00",	--2921
		x"4d",	--2922
		x"00",	--2923
		x"41",	--2924
		x"50",	--2925
		x"00",	--2926
		x"41",	--2927
		x"52",	--2928
		x"12",	--2929
		x"e0",	--2930
		x"41",	--2931
		x"50",	--2932
		x"00",	--2933
		x"41",	--2934
		x"12",	--2935
		x"e0",	--2936
		x"41",	--2937
		x"52",	--2938
		x"41",	--2939
		x"50",	--2940
		x"00",	--2941
		x"41",	--2942
		x"50",	--2943
		x"00",	--2944
		x"12",	--2945
		x"d4",	--2946
		x"12",	--2947
		x"de",	--2948
		x"50",	--2949
		x"00",	--2950
		x"41",	--2951
		x"50",	--2952
		x"ff",	--2953
		x"4e",	--2954
		x"00",	--2955
		x"4f",	--2956
		x"00",	--2957
		x"4c",	--2958
		x"00",	--2959
		x"4d",	--2960
		x"00",	--2961
		x"41",	--2962
		x"50",	--2963
		x"00",	--2964
		x"41",	--2965
		x"52",	--2966
		x"12",	--2967
		x"e0",	--2968
		x"41",	--2969
		x"50",	--2970
		x"00",	--2971
		x"41",	--2972
		x"12",	--2973
		x"e0",	--2974
		x"e3",	--2975
		x"00",	--2976
		x"41",	--2977
		x"52",	--2978
		x"41",	--2979
		x"50",	--2980
		x"00",	--2981
		x"41",	--2982
		x"50",	--2983
		x"00",	--2984
		x"12",	--2985
		x"d4",	--2986
		x"12",	--2987
		x"de",	--2988
		x"50",	--2989
		x"00",	--2990
		x"41",	--2991
		x"12",	--2992
		x"12",	--2993
		x"12",	--2994
		x"12",	--2995
		x"12",	--2996
		x"12",	--2997
		x"12",	--2998
		x"12",	--2999
		x"50",	--3000
		x"ff",	--3001
		x"4e",	--3002
		x"00",	--3003
		x"4f",	--3004
		x"00",	--3005
		x"4c",	--3006
		x"00",	--3007
		x"4d",	--3008
		x"00",	--3009
		x"41",	--3010
		x"50",	--3011
		x"00",	--3012
		x"41",	--3013
		x"52",	--3014
		x"12",	--3015
		x"e0",	--3016
		x"41",	--3017
		x"50",	--3018
		x"00",	--3019
		x"41",	--3020
		x"12",	--3021
		x"e0",	--3022
		x"41",	--3023
		x"00",	--3024
		x"93",	--3025
		x"28",	--3026
		x"41",	--3027
		x"00",	--3028
		x"93",	--3029
		x"28",	--3030
		x"92",	--3031
		x"24",	--3032
		x"92",	--3033
		x"24",	--3034
		x"93",	--3035
		x"24",	--3036
		x"93",	--3037
		x"24",	--3038
		x"41",	--3039
		x"00",	--3040
		x"41",	--3041
		x"00",	--3042
		x"41",	--3043
		x"00",	--3044
		x"41",	--3045
		x"00",	--3046
		x"40",	--3047
		x"00",	--3048
		x"43",	--3049
		x"43",	--3050
		x"43",	--3051
		x"43",	--3052
		x"43",	--3053
		x"00",	--3054
		x"43",	--3055
		x"00",	--3056
		x"43",	--3057
		x"43",	--3058
		x"4c",	--3059
		x"00",	--3060
		x"3c",	--3061
		x"58",	--3062
		x"69",	--3063
		x"c3",	--3064
		x"10",	--3065
		x"10",	--3066
		x"53",	--3067
		x"00",	--3068
		x"24",	--3069
		x"b3",	--3070
		x"24",	--3071
		x"58",	--3072
		x"69",	--3073
		x"56",	--3074
		x"67",	--3075
		x"43",	--3076
		x"43",	--3077
		x"99",	--3078
		x"28",	--3079
		x"24",	--3080
		x"43",	--3081
		x"43",	--3082
		x"5c",	--3083
		x"6d",	--3084
		x"56",	--3085
		x"67",	--3086
		x"93",	--3087
		x"37",	--3088
		x"d3",	--3089
		x"d3",	--3090
		x"3f",	--3091
		x"98",	--3092
		x"2b",	--3093
		x"3f",	--3094
		x"4a",	--3095
		x"00",	--3096
		x"4b",	--3097
		x"00",	--3098
		x"4f",	--3099
		x"41",	--3100
		x"00",	--3101
		x"51",	--3102
		x"00",	--3103
		x"4a",	--3104
		x"53",	--3105
		x"46",	--3106
		x"00",	--3107
		x"43",	--3108
		x"91",	--3109
		x"00",	--3110
		x"00",	--3111
		x"24",	--3112
		x"4d",	--3113
		x"00",	--3114
		x"93",	--3115
		x"38",	--3116
		x"90",	--3117
		x"40",	--3118
		x"2c",	--3119
		x"41",	--3120
		x"00",	--3121
		x"53",	--3122
		x"41",	--3123
		x"00",	--3124
		x"41",	--3125
		x"00",	--3126
		x"4d",	--3127
		x"5e",	--3128
		x"6f",	--3129
		x"93",	--3130
		x"38",	--3131
		x"5a",	--3132
		x"6b",	--3133
		x"53",	--3134
		x"90",	--3135
		x"40",	--3136
		x"2b",	--3137
		x"4a",	--3138
		x"00",	--3139
		x"4b",	--3140
		x"00",	--3141
		x"4c",	--3142
		x"00",	--3143
		x"4e",	--3144
		x"4f",	--3145
		x"f0",	--3146
		x"00",	--3147
		x"f3",	--3148
		x"90",	--3149
		x"00",	--3150
		x"24",	--3151
		x"4e",	--3152
		x"00",	--3153
		x"4f",	--3154
		x"00",	--3155
		x"40",	--3156
		x"00",	--3157
		x"00",	--3158
		x"41",	--3159
		x"52",	--3160
		x"12",	--3161
		x"de",	--3162
		x"50",	--3163
		x"00",	--3164
		x"41",	--3165
		x"41",	--3166
		x"41",	--3167
		x"41",	--3168
		x"41",	--3169
		x"41",	--3170
		x"41",	--3171
		x"41",	--3172
		x"41",	--3173
		x"d3",	--3174
		x"d3",	--3175
		x"3f",	--3176
		x"50",	--3177
		x"00",	--3178
		x"4a",	--3179
		x"b3",	--3180
		x"24",	--3181
		x"41",	--3182
		x"00",	--3183
		x"41",	--3184
		x"00",	--3185
		x"c3",	--3186
		x"10",	--3187
		x"10",	--3188
		x"4c",	--3189
		x"4d",	--3190
		x"d3",	--3191
		x"d0",	--3192
		x"80",	--3193
		x"46",	--3194
		x"00",	--3195
		x"47",	--3196
		x"00",	--3197
		x"c3",	--3198
		x"10",	--3199
		x"10",	--3200
		x"53",	--3201
		x"93",	--3202
		x"3b",	--3203
		x"48",	--3204
		x"00",	--3205
		x"3f",	--3206
		x"93",	--3207
		x"24",	--3208
		x"43",	--3209
		x"91",	--3210
		x"00",	--3211
		x"00",	--3212
		x"24",	--3213
		x"4f",	--3214
		x"00",	--3215
		x"41",	--3216
		x"50",	--3217
		x"00",	--3218
		x"3f",	--3219
		x"93",	--3220
		x"23",	--3221
		x"4e",	--3222
		x"4f",	--3223
		x"f0",	--3224
		x"00",	--3225
		x"f3",	--3226
		x"93",	--3227
		x"23",	--3228
		x"93",	--3229
		x"23",	--3230
		x"93",	--3231
		x"00",	--3232
		x"20",	--3233
		x"93",	--3234
		x"00",	--3235
		x"27",	--3236
		x"50",	--3237
		x"00",	--3238
		x"63",	--3239
		x"f0",	--3240
		x"ff",	--3241
		x"f3",	--3242
		x"3f",	--3243
		x"43",	--3244
		x"3f",	--3245
		x"43",	--3246
		x"3f",	--3247
		x"43",	--3248
		x"91",	--3249
		x"00",	--3250
		x"00",	--3251
		x"24",	--3252
		x"4f",	--3253
		x"00",	--3254
		x"41",	--3255
		x"50",	--3256
		x"00",	--3257
		x"3f",	--3258
		x"43",	--3259
		x"3f",	--3260
		x"93",	--3261
		x"23",	--3262
		x"40",	--3263
		x"ef",	--3264
		x"3f",	--3265
		x"12",	--3266
		x"12",	--3267
		x"12",	--3268
		x"12",	--3269
		x"12",	--3270
		x"50",	--3271
		x"ff",	--3272
		x"4e",	--3273
		x"00",	--3274
		x"4f",	--3275
		x"00",	--3276
		x"4c",	--3277
		x"00",	--3278
		x"4d",	--3279
		x"00",	--3280
		x"41",	--3281
		x"50",	--3282
		x"00",	--3283
		x"41",	--3284
		x"52",	--3285
		x"12",	--3286
		x"e0",	--3287
		x"41",	--3288
		x"52",	--3289
		x"41",	--3290
		x"12",	--3291
		x"e0",	--3292
		x"41",	--3293
		x"00",	--3294
		x"93",	--3295
		x"28",	--3296
		x"41",	--3297
		x"00",	--3298
		x"93",	--3299
		x"28",	--3300
		x"e1",	--3301
		x"00",	--3302
		x"00",	--3303
		x"92",	--3304
		x"24",	--3305
		x"93",	--3306
		x"24",	--3307
		x"92",	--3308
		x"24",	--3309
		x"93",	--3310
		x"24",	--3311
		x"41",	--3312
		x"00",	--3313
		x"81",	--3314
		x"00",	--3315
		x"4d",	--3316
		x"00",	--3317
		x"41",	--3318
		x"00",	--3319
		x"41",	--3320
		x"00",	--3321
		x"41",	--3322
		x"00",	--3323
		x"41",	--3324
		x"00",	--3325
		x"99",	--3326
		x"2c",	--3327
		x"5e",	--3328
		x"6f",	--3329
		x"53",	--3330
		x"4d",	--3331
		x"00",	--3332
		x"40",	--3333
		x"00",	--3334
		x"43",	--3335
		x"40",	--3336
		x"40",	--3337
		x"43",	--3338
		x"43",	--3339
		x"3c",	--3340
		x"dc",	--3341
		x"dd",	--3342
		x"88",	--3343
		x"79",	--3344
		x"c3",	--3345
		x"10",	--3346
		x"10",	--3347
		x"5e",	--3348
		x"6f",	--3349
		x"53",	--3350
		x"24",	--3351
		x"99",	--3352
		x"2b",	--3353
		x"23",	--3354
		x"98",	--3355
		x"2b",	--3356
		x"3f",	--3357
		x"9f",	--3358
		x"2b",	--3359
		x"98",	--3360
		x"2f",	--3361
		x"3f",	--3362
		x"4a",	--3363
		x"4b",	--3364
		x"f0",	--3365
		x"00",	--3366
		x"f3",	--3367
		x"90",	--3368
		x"00",	--3369
		x"24",	--3370
		x"4a",	--3371
		x"00",	--3372
		x"4b",	--3373
		x"00",	--3374
		x"41",	--3375
		x"50",	--3376
		x"00",	--3377
		x"12",	--3378
		x"de",	--3379
		x"50",	--3380
		x"00",	--3381
		x"41",	--3382
		x"41",	--3383
		x"41",	--3384
		x"41",	--3385
		x"41",	--3386
		x"41",	--3387
		x"42",	--3388
		x"00",	--3389
		x"41",	--3390
		x"50",	--3391
		x"00",	--3392
		x"3f",	--3393
		x"9e",	--3394
		x"23",	--3395
		x"40",	--3396
		x"ef",	--3397
		x"3f",	--3398
		x"93",	--3399
		x"23",	--3400
		x"4a",	--3401
		x"4b",	--3402
		x"f0",	--3403
		x"00",	--3404
		x"f3",	--3405
		x"93",	--3406
		x"23",	--3407
		x"93",	--3408
		x"23",	--3409
		x"93",	--3410
		x"20",	--3411
		x"93",	--3412
		x"27",	--3413
		x"50",	--3414
		x"00",	--3415
		x"63",	--3416
		x"f0",	--3417
		x"ff",	--3418
		x"f3",	--3419
		x"3f",	--3420
		x"43",	--3421
		x"00",	--3422
		x"43",	--3423
		x"00",	--3424
		x"43",	--3425
		x"00",	--3426
		x"41",	--3427
		x"50",	--3428
		x"00",	--3429
		x"3f",	--3430
		x"41",	--3431
		x"52",	--3432
		x"3f",	--3433
		x"50",	--3434
		x"ff",	--3435
		x"4e",	--3436
		x"00",	--3437
		x"4f",	--3438
		x"00",	--3439
		x"4c",	--3440
		x"00",	--3441
		x"4d",	--3442
		x"00",	--3443
		x"41",	--3444
		x"50",	--3445
		x"00",	--3446
		x"41",	--3447
		x"52",	--3448
		x"12",	--3449
		x"e0",	--3450
		x"41",	--3451
		x"52",	--3452
		x"41",	--3453
		x"12",	--3454
		x"e0",	--3455
		x"93",	--3456
		x"00",	--3457
		x"28",	--3458
		x"93",	--3459
		x"00",	--3460
		x"28",	--3461
		x"41",	--3462
		x"52",	--3463
		x"41",	--3464
		x"50",	--3465
		x"00",	--3466
		x"12",	--3467
		x"e1",	--3468
		x"50",	--3469
		x"00",	--3470
		x"41",	--3471
		x"43",	--3472
		x"3f",	--3473
		x"50",	--3474
		x"ff",	--3475
		x"4e",	--3476
		x"00",	--3477
		x"4f",	--3478
		x"00",	--3479
		x"4c",	--3480
		x"00",	--3481
		x"4d",	--3482
		x"00",	--3483
		x"41",	--3484
		x"50",	--3485
		x"00",	--3486
		x"41",	--3487
		x"52",	--3488
		x"12",	--3489
		x"e0",	--3490
		x"41",	--3491
		x"52",	--3492
		x"41",	--3493
		x"12",	--3494
		x"e0",	--3495
		x"93",	--3496
		x"00",	--3497
		x"28",	--3498
		x"93",	--3499
		x"00",	--3500
		x"28",	--3501
		x"41",	--3502
		x"52",	--3503
		x"41",	--3504
		x"50",	--3505
		x"00",	--3506
		x"12",	--3507
		x"e1",	--3508
		x"50",	--3509
		x"00",	--3510
		x"41",	--3511
		x"43",	--3512
		x"3f",	--3513
		x"50",	--3514
		x"ff",	--3515
		x"4e",	--3516
		x"00",	--3517
		x"4f",	--3518
		x"00",	--3519
		x"4c",	--3520
		x"00",	--3521
		x"4d",	--3522
		x"00",	--3523
		x"41",	--3524
		x"50",	--3525
		x"00",	--3526
		x"41",	--3527
		x"52",	--3528
		x"12",	--3529
		x"e0",	--3530
		x"41",	--3531
		x"52",	--3532
		x"41",	--3533
		x"12",	--3534
		x"e0",	--3535
		x"93",	--3536
		x"00",	--3537
		x"28",	--3538
		x"93",	--3539
		x"00",	--3540
		x"28",	--3541
		x"41",	--3542
		x"52",	--3543
		x"41",	--3544
		x"50",	--3545
		x"00",	--3546
		x"12",	--3547
		x"e1",	--3548
		x"50",	--3549
		x"00",	--3550
		x"41",	--3551
		x"43",	--3552
		x"3f",	--3553
		x"12",	--3554
		x"12",	--3555
		x"82",	--3556
		x"40",	--3557
		x"00",	--3558
		x"00",	--3559
		x"4f",	--3560
		x"5d",	--3561
		x"43",	--3562
		x"6d",	--3563
		x"4d",	--3564
		x"4d",	--3565
		x"00",	--3566
		x"93",	--3567
		x"20",	--3568
		x"93",	--3569
		x"20",	--3570
		x"43",	--3571
		x"00",	--3572
		x"41",	--3573
		x"12",	--3574
		x"de",	--3575
		x"52",	--3576
		x"41",	--3577
		x"41",	--3578
		x"41",	--3579
		x"40",	--3580
		x"00",	--3581
		x"00",	--3582
		x"93",	--3583
		x"20",	--3584
		x"4e",	--3585
		x"4f",	--3586
		x"4a",	--3587
		x"00",	--3588
		x"4b",	--3589
		x"00",	--3590
		x"4a",	--3591
		x"4b",	--3592
		x"12",	--3593
		x"dd",	--3594
		x"53",	--3595
		x"93",	--3596
		x"3b",	--3597
		x"4a",	--3598
		x"00",	--3599
		x"4b",	--3600
		x"00",	--3601
		x"4f",	--3602
		x"f0",	--3603
		x"00",	--3604
		x"20",	--3605
		x"40",	--3606
		x"00",	--3607
		x"8f",	--3608
		x"4e",	--3609
		x"00",	--3610
		x"3f",	--3611
		x"93",	--3612
		x"24",	--3613
		x"4e",	--3614
		x"4f",	--3615
		x"e3",	--3616
		x"e3",	--3617
		x"53",	--3618
		x"63",	--3619
		x"3f",	--3620
		x"51",	--3621
		x"00",	--3622
		x"00",	--3623
		x"61",	--3624
		x"00",	--3625
		x"00",	--3626
		x"53",	--3627
		x"23",	--3628
		x"3f",	--3629
		x"90",	--3630
		x"80",	--3631
		x"23",	--3632
		x"43",	--3633
		x"40",	--3634
		x"cf",	--3635
		x"3f",	--3636
		x"50",	--3637
		x"ff",	--3638
		x"4e",	--3639
		x"00",	--3640
		x"4f",	--3641
		x"00",	--3642
		x"41",	--3643
		x"52",	--3644
		x"41",	--3645
		x"12",	--3646
		x"e0",	--3647
		x"41",	--3648
		x"00",	--3649
		x"93",	--3650
		x"24",	--3651
		x"28",	--3652
		x"92",	--3653
		x"24",	--3654
		x"41",	--3655
		x"00",	--3656
		x"93",	--3657
		x"38",	--3658
		x"90",	--3659
		x"00",	--3660
		x"38",	--3661
		x"93",	--3662
		x"00",	--3663
		x"20",	--3664
		x"43",	--3665
		x"40",	--3666
		x"7f",	--3667
		x"50",	--3668
		x"00",	--3669
		x"41",	--3670
		x"41",	--3671
		x"00",	--3672
		x"41",	--3673
		x"00",	--3674
		x"40",	--3675
		x"00",	--3676
		x"8d",	--3677
		x"4c",	--3678
		x"f0",	--3679
		x"00",	--3680
		x"20",	--3681
		x"93",	--3682
		x"00",	--3683
		x"27",	--3684
		x"e3",	--3685
		x"e3",	--3686
		x"53",	--3687
		x"63",	--3688
		x"50",	--3689
		x"00",	--3690
		x"41",	--3691
		x"43",	--3692
		x"43",	--3693
		x"50",	--3694
		x"00",	--3695
		x"41",	--3696
		x"c3",	--3697
		x"10",	--3698
		x"10",	--3699
		x"53",	--3700
		x"23",	--3701
		x"3f",	--3702
		x"43",	--3703
		x"40",	--3704
		x"80",	--3705
		x"50",	--3706
		x"00",	--3707
		x"41",	--3708
		x"12",	--3709
		x"12",	--3710
		x"12",	--3711
		x"12",	--3712
		x"82",	--3713
		x"4e",	--3714
		x"4f",	--3715
		x"43",	--3716
		x"00",	--3717
		x"93",	--3718
		x"20",	--3719
		x"93",	--3720
		x"20",	--3721
		x"43",	--3722
		x"00",	--3723
		x"41",	--3724
		x"12",	--3725
		x"de",	--3726
		x"52",	--3727
		x"41",	--3728
		x"41",	--3729
		x"41",	--3730
		x"41",	--3731
		x"41",	--3732
		x"40",	--3733
		x"00",	--3734
		x"00",	--3735
		x"40",	--3736
		x"00",	--3737
		x"00",	--3738
		x"4a",	--3739
		x"00",	--3740
		x"4b",	--3741
		x"00",	--3742
		x"4a",	--3743
		x"4b",	--3744
		x"12",	--3745
		x"dd",	--3746
		x"53",	--3747
		x"93",	--3748
		x"38",	--3749
		x"27",	--3750
		x"4a",	--3751
		x"00",	--3752
		x"4b",	--3753
		x"00",	--3754
		x"4f",	--3755
		x"f0",	--3756
		x"00",	--3757
		x"20",	--3758
		x"40",	--3759
		x"00",	--3760
		x"8f",	--3761
		x"4e",	--3762
		x"00",	--3763
		x"3f",	--3764
		x"51",	--3765
		x"00",	--3766
		x"00",	--3767
		x"61",	--3768
		x"00",	--3769
		x"00",	--3770
		x"53",	--3771
		x"23",	--3772
		x"3f",	--3773
		x"4f",	--3774
		x"e3",	--3775
		x"53",	--3776
		x"43",	--3777
		x"43",	--3778
		x"4e",	--3779
		x"f0",	--3780
		x"00",	--3781
		x"24",	--3782
		x"5c",	--3783
		x"6d",	--3784
		x"53",	--3785
		x"23",	--3786
		x"53",	--3787
		x"63",	--3788
		x"fa",	--3789
		x"fb",	--3790
		x"43",	--3791
		x"43",	--3792
		x"93",	--3793
		x"20",	--3794
		x"93",	--3795
		x"20",	--3796
		x"43",	--3797
		x"43",	--3798
		x"f0",	--3799
		x"00",	--3800
		x"20",	--3801
		x"48",	--3802
		x"49",	--3803
		x"da",	--3804
		x"db",	--3805
		x"4d",	--3806
		x"00",	--3807
		x"4e",	--3808
		x"00",	--3809
		x"40",	--3810
		x"00",	--3811
		x"8f",	--3812
		x"4e",	--3813
		x"00",	--3814
		x"3f",	--3815
		x"c3",	--3816
		x"10",	--3817
		x"10",	--3818
		x"53",	--3819
		x"23",	--3820
		x"3f",	--3821
		x"12",	--3822
		x"12",	--3823
		x"12",	--3824
		x"93",	--3825
		x"2c",	--3826
		x"90",	--3827
		x"01",	--3828
		x"28",	--3829
		x"40",	--3830
		x"00",	--3831
		x"43",	--3832
		x"42",	--3833
		x"4e",	--3834
		x"4f",	--3835
		x"49",	--3836
		x"93",	--3837
		x"20",	--3838
		x"50",	--3839
		x"ef",	--3840
		x"4c",	--3841
		x"43",	--3842
		x"8e",	--3843
		x"7f",	--3844
		x"4a",	--3845
		x"41",	--3846
		x"41",	--3847
		x"41",	--3848
		x"41",	--3849
		x"90",	--3850
		x"01",	--3851
		x"28",	--3852
		x"42",	--3853
		x"43",	--3854
		x"40",	--3855
		x"00",	--3856
		x"4e",	--3857
		x"4f",	--3858
		x"49",	--3859
		x"93",	--3860
		x"27",	--3861
		x"c3",	--3862
		x"10",	--3863
		x"10",	--3864
		x"53",	--3865
		x"23",	--3866
		x"3f",	--3867
		x"40",	--3868
		x"00",	--3869
		x"43",	--3870
		x"40",	--3871
		x"00",	--3872
		x"3f",	--3873
		x"40",	--3874
		x"00",	--3875
		x"43",	--3876
		x"43",	--3877
		x"3f",	--3878
		x"12",	--3879
		x"12",	--3880
		x"12",	--3881
		x"12",	--3882
		x"12",	--3883
		x"4f",	--3884
		x"4f",	--3885
		x"00",	--3886
		x"4f",	--3887
		x"00",	--3888
		x"4d",	--3889
		x"00",	--3890
		x"4d",	--3891
		x"93",	--3892
		x"28",	--3893
		x"92",	--3894
		x"24",	--3895
		x"93",	--3896
		x"24",	--3897
		x"93",	--3898
		x"24",	--3899
		x"4d",	--3900
		x"00",	--3901
		x"90",	--3902
		x"ff",	--3903
		x"38",	--3904
		x"90",	--3905
		x"00",	--3906
		x"34",	--3907
		x"4e",	--3908
		x"4f",	--3909
		x"f0",	--3910
		x"00",	--3911
		x"f3",	--3912
		x"90",	--3913
		x"00",	--3914
		x"24",	--3915
		x"50",	--3916
		x"00",	--3917
		x"63",	--3918
		x"93",	--3919
		x"38",	--3920
		x"4b",	--3921
		x"50",	--3922
		x"00",	--3923
		x"c3",	--3924
		x"10",	--3925
		x"10",	--3926
		x"c3",	--3927
		x"10",	--3928
		x"10",	--3929
		x"c3",	--3930
		x"10",	--3931
		x"10",	--3932
		x"c3",	--3933
		x"10",	--3934
		x"10",	--3935
		x"c3",	--3936
		x"10",	--3937
		x"10",	--3938
		x"c3",	--3939
		x"10",	--3940
		x"10",	--3941
		x"c3",	--3942
		x"10",	--3943
		x"10",	--3944
		x"f3",	--3945
		x"f0",	--3946
		x"00",	--3947
		x"4d",	--3948
		x"3c",	--3949
		x"93",	--3950
		x"23",	--3951
		x"43",	--3952
		x"43",	--3953
		x"43",	--3954
		x"4d",	--3955
		x"5d",	--3956
		x"5d",	--3957
		x"5d",	--3958
		x"5d",	--3959
		x"5d",	--3960
		x"5d",	--3961
		x"5d",	--3962
		x"4f",	--3963
		x"f0",	--3964
		x"00",	--3965
		x"dd",	--3966
		x"4a",	--3967
		x"11",	--3968
		x"43",	--3969
		x"10",	--3970
		x"4c",	--3971
		x"df",	--3972
		x"4d",	--3973
		x"41",	--3974
		x"41",	--3975
		x"41",	--3976
		x"41",	--3977
		x"41",	--3978
		x"41",	--3979
		x"93",	--3980
		x"23",	--3981
		x"4e",	--3982
		x"4f",	--3983
		x"f0",	--3984
		x"00",	--3985
		x"f3",	--3986
		x"93",	--3987
		x"20",	--3988
		x"93",	--3989
		x"27",	--3990
		x"50",	--3991
		x"00",	--3992
		x"63",	--3993
		x"3f",	--3994
		x"c3",	--3995
		x"10",	--3996
		x"10",	--3997
		x"4b",	--3998
		x"50",	--3999
		x"00",	--4000
		x"3f",	--4001
		x"43",	--4002
		x"43",	--4003
		x"43",	--4004
		x"3f",	--4005
		x"d3",	--4006
		x"d0",	--4007
		x"00",	--4008
		x"f3",	--4009
		x"f0",	--4010
		x"00",	--4011
		x"43",	--4012
		x"3f",	--4013
		x"40",	--4014
		x"ff",	--4015
		x"8b",	--4016
		x"90",	--4017
		x"00",	--4018
		x"34",	--4019
		x"4e",	--4020
		x"4f",	--4021
		x"47",	--4022
		x"f0",	--4023
		x"00",	--4024
		x"24",	--4025
		x"c3",	--4026
		x"10",	--4027
		x"10",	--4028
		x"53",	--4029
		x"23",	--4030
		x"43",	--4031
		x"43",	--4032
		x"f0",	--4033
		x"00",	--4034
		x"24",	--4035
		x"58",	--4036
		x"69",	--4037
		x"53",	--4038
		x"23",	--4039
		x"53",	--4040
		x"63",	--4041
		x"fe",	--4042
		x"ff",	--4043
		x"43",	--4044
		x"43",	--4045
		x"93",	--4046
		x"20",	--4047
		x"93",	--4048
		x"20",	--4049
		x"43",	--4050
		x"43",	--4051
		x"4e",	--4052
		x"4f",	--4053
		x"dc",	--4054
		x"dd",	--4055
		x"48",	--4056
		x"49",	--4057
		x"f0",	--4058
		x"00",	--4059
		x"f3",	--4060
		x"90",	--4061
		x"00",	--4062
		x"24",	--4063
		x"50",	--4064
		x"00",	--4065
		x"63",	--4066
		x"48",	--4067
		x"49",	--4068
		x"c3",	--4069
		x"10",	--4070
		x"10",	--4071
		x"c3",	--4072
		x"10",	--4073
		x"10",	--4074
		x"c3",	--4075
		x"10",	--4076
		x"10",	--4077
		x"c3",	--4078
		x"10",	--4079
		x"10",	--4080
		x"c3",	--4081
		x"10",	--4082
		x"10",	--4083
		x"c3",	--4084
		x"10",	--4085
		x"10",	--4086
		x"c3",	--4087
		x"10",	--4088
		x"10",	--4089
		x"f3",	--4090
		x"f0",	--4091
		x"00",	--4092
		x"43",	--4093
		x"90",	--4094
		x"40",	--4095
		x"2f",	--4096
		x"43",	--4097
		x"3f",	--4098
		x"43",	--4099
		x"43",	--4100
		x"3f",	--4101
		x"93",	--4102
		x"23",	--4103
		x"48",	--4104
		x"49",	--4105
		x"f0",	--4106
		x"00",	--4107
		x"f3",	--4108
		x"93",	--4109
		x"24",	--4110
		x"50",	--4111
		x"00",	--4112
		x"63",	--4113
		x"3f",	--4114
		x"93",	--4115
		x"27",	--4116
		x"3f",	--4117
		x"12",	--4118
		x"12",	--4119
		x"4f",	--4120
		x"4f",	--4121
		x"00",	--4122
		x"f0",	--4123
		x"00",	--4124
		x"4f",	--4125
		x"00",	--4126
		x"c3",	--4127
		x"10",	--4128
		x"c3",	--4129
		x"10",	--4130
		x"c3",	--4131
		x"10",	--4132
		x"c3",	--4133
		x"10",	--4134
		x"c3",	--4135
		x"10",	--4136
		x"c3",	--4137
		x"10",	--4138
		x"c3",	--4139
		x"10",	--4140
		x"4d",	--4141
		x"4f",	--4142
		x"00",	--4143
		x"b0",	--4144
		x"00",	--4145
		x"43",	--4146
		x"6f",	--4147
		x"4f",	--4148
		x"00",	--4149
		x"93",	--4150
		x"20",	--4151
		x"93",	--4152
		x"24",	--4153
		x"40",	--4154
		x"ff",	--4155
		x"00",	--4156
		x"4a",	--4157
		x"4b",	--4158
		x"5c",	--4159
		x"6d",	--4160
		x"5c",	--4161
		x"6d",	--4162
		x"5c",	--4163
		x"6d",	--4164
		x"5c",	--4165
		x"6d",	--4166
		x"5c",	--4167
		x"6d",	--4168
		x"5c",	--4169
		x"6d",	--4170
		x"5c",	--4171
		x"6d",	--4172
		x"40",	--4173
		x"00",	--4174
		x"00",	--4175
		x"90",	--4176
		x"40",	--4177
		x"2c",	--4178
		x"40",	--4179
		x"ff",	--4180
		x"5c",	--4181
		x"6d",	--4182
		x"4f",	--4183
		x"53",	--4184
		x"90",	--4185
		x"40",	--4186
		x"2b",	--4187
		x"4a",	--4188
		x"00",	--4189
		x"4c",	--4190
		x"00",	--4191
		x"4d",	--4192
		x"00",	--4193
		x"41",	--4194
		x"41",	--4195
		x"41",	--4196
		x"90",	--4197
		x"00",	--4198
		x"24",	--4199
		x"50",	--4200
		x"ff",	--4201
		x"4d",	--4202
		x"00",	--4203
		x"40",	--4204
		x"00",	--4205
		x"00",	--4206
		x"4a",	--4207
		x"4b",	--4208
		x"5c",	--4209
		x"6d",	--4210
		x"5c",	--4211
		x"6d",	--4212
		x"5c",	--4213
		x"6d",	--4214
		x"5c",	--4215
		x"6d",	--4216
		x"5c",	--4217
		x"6d",	--4218
		x"5c",	--4219
		x"6d",	--4220
		x"5c",	--4221
		x"6d",	--4222
		x"4c",	--4223
		x"4d",	--4224
		x"d3",	--4225
		x"d0",	--4226
		x"40",	--4227
		x"4a",	--4228
		x"00",	--4229
		x"4b",	--4230
		x"00",	--4231
		x"41",	--4232
		x"41",	--4233
		x"41",	--4234
		x"93",	--4235
		x"23",	--4236
		x"43",	--4237
		x"00",	--4238
		x"41",	--4239
		x"41",	--4240
		x"41",	--4241
		x"93",	--4242
		x"24",	--4243
		x"4a",	--4244
		x"4b",	--4245
		x"f3",	--4246
		x"f0",	--4247
		x"00",	--4248
		x"93",	--4249
		x"20",	--4250
		x"93",	--4251
		x"24",	--4252
		x"43",	--4253
		x"00",	--4254
		x"3f",	--4255
		x"93",	--4256
		x"23",	--4257
		x"42",	--4258
		x"00",	--4259
		x"3f",	--4260
		x"43",	--4261
		x"00",	--4262
		x"3f",	--4263
		x"12",	--4264
		x"4f",	--4265
		x"93",	--4266
		x"28",	--4267
		x"4e",	--4268
		x"93",	--4269
		x"28",	--4270
		x"92",	--4271
		x"24",	--4272
		x"92",	--4273
		x"24",	--4274
		x"93",	--4275
		x"24",	--4276
		x"93",	--4277
		x"24",	--4278
		x"4f",	--4279
		x"00",	--4280
		x"9e",	--4281
		x"00",	--4282
		x"24",	--4283
		x"93",	--4284
		x"20",	--4285
		x"43",	--4286
		x"4e",	--4287
		x"41",	--4288
		x"41",	--4289
		x"93",	--4290
		x"24",	--4291
		x"93",	--4292
		x"00",	--4293
		x"23",	--4294
		x"43",	--4295
		x"4e",	--4296
		x"41",	--4297
		x"41",	--4298
		x"93",	--4299
		x"00",	--4300
		x"27",	--4301
		x"43",	--4302
		x"3f",	--4303
		x"4f",	--4304
		x"00",	--4305
		x"4e",	--4306
		x"00",	--4307
		x"9b",	--4308
		x"3b",	--4309
		x"9c",	--4310
		x"38",	--4311
		x"4f",	--4312
		x"00",	--4313
		x"4f",	--4314
		x"00",	--4315
		x"4e",	--4316
		x"00",	--4317
		x"4e",	--4318
		x"00",	--4319
		x"9f",	--4320
		x"2b",	--4321
		x"9e",	--4322
		x"28",	--4323
		x"9b",	--4324
		x"2b",	--4325
		x"9e",	--4326
		x"28",	--4327
		x"9f",	--4328
		x"28",	--4329
		x"9c",	--4330
		x"28",	--4331
		x"43",	--4332
		x"3f",	--4333
		x"93",	--4334
		x"23",	--4335
		x"43",	--4336
		x"3f",	--4337
		x"92",	--4338
		x"23",	--4339
		x"4e",	--4340
		x"00",	--4341
		x"4f",	--4342
		x"00",	--4343
		x"8f",	--4344
		x"3f",	--4345
		x"42",	--4346
		x"02",	--4347
		x"93",	--4348
		x"38",	--4349
		x"42",	--4350
		x"02",	--4351
		x"4f",	--4352
		x"00",	--4353
		x"53",	--4354
		x"4d",	--4355
		x"02",	--4356
		x"53",	--4357
		x"4e",	--4358
		x"02",	--4359
		x"41",	--4360
		x"43",	--4361
		x"41",	--4362
		x"12",	--4363
		x"12",	--4364
		x"83",	--4365
		x"4e",	--4366
		x"00",	--4367
		x"42",	--4368
		x"02",	--4369
		x"42",	--4370
		x"02",	--4371
		x"4e",	--4372
		x"4f",	--4373
		x"40",	--4374
		x"e1",	--4375
		x"12",	--4376
		x"e4",	--4377
		x"9b",	--4378
		x"38",	--4379
		x"4a",	--4380
		x"5b",	--4381
		x"43",	--4382
		x"ff",	--4383
		x"3c",	--4384
		x"42",	--4385
		x"02",	--4386
		x"43",	--4387
		x"00",	--4388
		x"53",	--4389
		x"41",	--4390
		x"41",	--4391
		x"41",	--4392
		x"41",	--4393
		x"00",	--4394
		x"02",	--4395
		x"40",	--4396
		x"7f",	--4397
		x"02",	--4398
		x"41",	--4399
		x"50",	--4400
		x"00",	--4401
		x"41",	--4402
		x"00",	--4403
		x"12",	--4404
		x"e2",	--4405
		x"41",	--4406
		x"41",	--4407
		x"00",	--4408
		x"02",	--4409
		x"41",	--4410
		x"00",	--4411
		x"02",	--4412
		x"41",	--4413
		x"52",	--4414
		x"41",	--4415
		x"00",	--4416
		x"12",	--4417
		x"e2",	--4418
		x"41",	--4419
		x"4e",	--4420
		x"4f",	--4421
		x"02",	--4422
		x"40",	--4423
		x"7f",	--4424
		x"02",	--4425
		x"4d",	--4426
		x"4c",	--4427
		x"12",	--4428
		x"e2",	--4429
		x"41",	--4430
		x"4f",	--4431
		x"02",	--4432
		x"4e",	--4433
		x"02",	--4434
		x"4c",	--4435
		x"4d",	--4436
		x"12",	--4437
		x"e2",	--4438
		x"41",	--4439
		x"12",	--4440
		x"12",	--4441
		x"12",	--4442
		x"12",	--4443
		x"12",	--4444
		x"12",	--4445
		x"12",	--4446
		x"12",	--4447
		x"82",	--4448
		x"4f",	--4449
		x"4e",	--4450
		x"00",	--4451
		x"4d",	--4452
		x"41",	--4453
		x"00",	--4454
		x"41",	--4455
		x"00",	--4456
		x"4d",	--4457
		x"4d",	--4458
		x"10",	--4459
		x"44",	--4460
		x"4f",	--4461
		x"b0",	--4462
		x"00",	--4463
		x"24",	--4464
		x"40",	--4465
		x"00",	--4466
		x"00",	--4467
		x"4f",	--4468
		x"10",	--4469
		x"f3",	--4470
		x"24",	--4471
		x"40",	--4472
		x"00",	--4473
		x"3c",	--4474
		x"40",	--4475
		x"00",	--4476
		x"4e",	--4477
		x"00",	--4478
		x"41",	--4479
		x"53",	--4480
		x"3c",	--4481
		x"f0",	--4482
		x"00",	--4483
		x"24",	--4484
		x"40",	--4485
		x"00",	--4486
		x"00",	--4487
		x"3c",	--4488
		x"93",	--4489
		x"24",	--4490
		x"4d",	--4491
		x"00",	--4492
		x"41",	--4493
		x"53",	--4494
		x"3c",	--4495
		x"41",	--4496
		x"4c",	--4497
		x"10",	--4498
		x"11",	--4499
		x"10",	--4500
		x"11",	--4501
		x"4c",	--4502
		x"41",	--4503
		x"41",	--4504
		x"10",	--4505
		x"11",	--4506
		x"10",	--4507
		x"11",	--4508
		x"4c",	--4509
		x"86",	--4510
		x"77",	--4511
		x"4f",	--4512
		x"10",	--4513
		x"4e",	--4514
		x"00",	--4515
		x"f2",	--4516
		x"24",	--4517
		x"45",	--4518
		x"3c",	--4519
		x"43",	--4520
		x"4f",	--4521
		x"b0",	--4522
		x"00",	--4523
		x"20",	--4524
		x"41",	--4525
		x"00",	--4526
		x"53",	--4527
		x"53",	--4528
		x"93",	--4529
		x"00",	--4530
		x"23",	--4531
		x"81",	--4532
		x"00",	--4533
		x"9a",	--4534
		x"28",	--4535
		x"8a",	--4536
		x"3c",	--4537
		x"43",	--4538
		x"b3",	--4539
		x"00",	--4540
		x"24",	--4541
		x"95",	--4542
		x"28",	--4543
		x"85",	--4544
		x"3c",	--4545
		x"43",	--4546
		x"4d",	--4547
		x"9d",	--4548
		x"2c",	--4549
		x"47",	--4550
		x"93",	--4551
		x"38",	--4552
		x"40",	--4553
		x"00",	--4554
		x"00",	--4555
		x"43",	--4556
		x"43",	--4557
		x"3c",	--4558
		x"41",	--4559
		x"56",	--4560
		x"4f",	--4561
		x"11",	--4562
		x"53",	--4563
		x"12",	--4564
		x"3c",	--4565
		x"43",	--4566
		x"9a",	--4567
		x"3b",	--4568
		x"4a",	--4569
		x"40",	--4570
		x"00",	--4571
		x"00",	--4572
		x"8b",	--4573
		x"3c",	--4574
		x"41",	--4575
		x"00",	--4576
		x"11",	--4577
		x"12",	--4578
		x"53",	--4579
		x"45",	--4580
		x"5b",	--4581
		x"99",	--4582
		x"2b",	--4583
		x"3c",	--4584
		x"43",	--4585
		x"43",	--4586
		x"3c",	--4587
		x"53",	--4588
		x"41",	--4589
		x"56",	--4590
		x"4f",	--4591
		x"11",	--4592
		x"53",	--4593
		x"12",	--4594
		x"9a",	--4595
		x"3b",	--4596
		x"b3",	--4597
		x"00",	--4598
		x"24",	--4599
		x"44",	--4600
		x"3c",	--4601
		x"41",	--4602
		x"00",	--4603
		x"8b",	--4604
		x"3c",	--4605
		x"40",	--4606
		x"00",	--4607
		x"12",	--4608
		x"53",	--4609
		x"93",	--4610
		x"23",	--4611
		x"44",	--4612
		x"54",	--4613
		x"3f",	--4614
		x"53",	--4615
		x"11",	--4616
		x"12",	--4617
		x"53",	--4618
		x"4a",	--4619
		x"5b",	--4620
		x"4f",	--4621
		x"93",	--4622
		x"24",	--4623
		x"93",	--4624
		x"23",	--4625
		x"3c",	--4626
		x"40",	--4627
		x"00",	--4628
		x"12",	--4629
		x"53",	--4630
		x"99",	--4631
		x"2b",	--4632
		x"4b",	--4633
		x"52",	--4634
		x"41",	--4635
		x"41",	--4636
		x"41",	--4637
		x"41",	--4638
		x"41",	--4639
		x"41",	--4640
		x"41",	--4641
		x"41",	--4642
		x"41",	--4643
		x"12",	--4644
		x"12",	--4645
		x"12",	--4646
		x"12",	--4647
		x"12",	--4648
		x"12",	--4649
		x"12",	--4650
		x"12",	--4651
		x"50",	--4652
		x"ff",	--4653
		x"4f",	--4654
		x"00",	--4655
		x"4e",	--4656
		x"4d",	--4657
		x"4e",	--4658
		x"00",	--4659
		x"43",	--4660
		x"00",	--4661
		x"43",	--4662
		x"00",	--4663
		x"43",	--4664
		x"00",	--4665
		x"43",	--4666
		x"00",	--4667
		x"43",	--4668
		x"00",	--4669
		x"43",	--4670
		x"00",	--4671
		x"43",	--4672
		x"43",	--4673
		x"00",	--4674
		x"41",	--4675
		x"50",	--4676
		x"00",	--4677
		x"4e",	--4678
		x"00",	--4679
		x"40",	--4680
		x"ea",	--4681
		x"46",	--4682
		x"53",	--4683
		x"4f",	--4684
		x"00",	--4685
		x"93",	--4686
		x"20",	--4687
		x"90",	--4688
		x"00",	--4689
		x"20",	--4690
		x"43",	--4691
		x"00",	--4692
		x"43",	--4693
		x"00",	--4694
		x"46",	--4695
		x"00",	--4696
		x"43",	--4697
		x"00",	--4698
		x"43",	--4699
		x"00",	--4700
		x"43",	--4701
		x"00",	--4702
		x"43",	--4703
		x"00",	--4704
		x"43",	--4705
		x"00",	--4706
		x"40",	--4707
		x"ea",	--4708
		x"47",	--4709
		x"11",	--4710
		x"4e",	--4711
		x"12",	--4712
		x"00",	--4713
		x"53",	--4714
		x"00",	--4715
		x"40",	--4716
		x"ea",	--4717
		x"90",	--4718
		x"00",	--4719
		x"24",	--4720
		x"90",	--4721
		x"00",	--4722
		x"34",	--4723
		x"90",	--4724
		x"00",	--4725
		x"24",	--4726
		x"90",	--4727
		x"00",	--4728
		x"34",	--4729
		x"90",	--4730
		x"00",	--4731
		x"24",	--4732
		x"90",	--4733
		x"00",	--4734
		x"34",	--4735
		x"90",	--4736
		x"00",	--4737
		x"24",	--4738
		x"90",	--4739
		x"00",	--4740
		x"27",	--4741
		x"90",	--4742
		x"00",	--4743
		x"20",	--4744
		x"3c",	--4745
		x"90",	--4746
		x"00",	--4747
		x"24",	--4748
		x"90",	--4749
		x"00",	--4750
		x"24",	--4751
		x"90",	--4752
		x"00",	--4753
		x"20",	--4754
		x"3c",	--4755
		x"90",	--4756
		x"00",	--4757
		x"38",	--4758
		x"90",	--4759
		x"00",	--4760
		x"20",	--4761
		x"3c",	--4762
		x"90",	--4763
		x"00",	--4764
		x"24",	--4765
		x"90",	--4766
		x"00",	--4767
		x"34",	--4768
		x"90",	--4769
		x"00",	--4770
		x"24",	--4771
		x"90",	--4772
		x"00",	--4773
		x"24",	--4774
		x"90",	--4775
		x"00",	--4776
		x"20",	--4777
		x"3c",	--4778
		x"90",	--4779
		x"00",	--4780
		x"24",	--4781
		x"90",	--4782
		x"00",	--4783
		x"34",	--4784
		x"90",	--4785
		x"00",	--4786
		x"20",	--4787
		x"3c",	--4788
		x"90",	--4789
		x"00",	--4790
		x"24",	--4791
		x"90",	--4792
		x"00",	--4793
		x"24",	--4794
		x"41",	--4795
		x"00",	--4796
		x"41",	--4797
		x"00",	--4798
		x"89",	--4799
		x"40",	--4800
		x"ea",	--4801
		x"42",	--4802
		x"00",	--4803
		x"3c",	--4804
		x"d2",	--4805
		x"00",	--4806
		x"40",	--4807
		x"ea",	--4808
		x"41",	--4809
		x"f3",	--4810
		x"41",	--4811
		x"24",	--4812
		x"f0",	--4813
		x"ff",	--4814
		x"d3",	--4815
		x"3c",	--4816
		x"d3",	--4817
		x"4e",	--4818
		x"00",	--4819
		x"40",	--4820
		x"ea",	--4821
		x"d0",	--4822
		x"00",	--4823
		x"00",	--4824
		x"40",	--4825
		x"ea",	--4826
		x"40",	--4827
		x"00",	--4828
		x"00",	--4829
		x"40",	--4830
		x"ea",	--4831
		x"90",	--4832
		x"00",	--4833
		x"00",	--4834
		x"20",	--4835
		x"40",	--4836
		x"ea",	--4837
		x"40",	--4838
		x"00",	--4839
		x"00",	--4840
		x"40",	--4841
		x"ea",	--4842
		x"93",	--4843
		x"00",	--4844
		x"24",	--4845
		x"40",	--4846
		x"ea",	--4847
		x"43",	--4848
		x"00",	--4849
		x"40",	--4850
		x"ea",	--4851
		x"45",	--4852
		x"53",	--4853
		x"45",	--4854
		x"93",	--4855
		x"38",	--4856
		x"4a",	--4857
		x"00",	--4858
		x"3c",	--4859
		x"93",	--4860
		x"00",	--4861
		x"24",	--4862
		x"40",	--4863
		x"ea",	--4864
		x"d0",	--4865
		x"00",	--4866
		x"00",	--4867
		x"e3",	--4868
		x"4a",	--4869
		x"00",	--4870
		x"53",	--4871
		x"00",	--4872
		x"4e",	--4873
		x"3c",	--4874
		x"93",	--4875
		x"00",	--4876
		x"20",	--4877
		x"93",	--4878
		x"00",	--4879
		x"20",	--4880
		x"41",	--4881
		x"f0",	--4882
		x"00",	--4883
		x"43",	--4884
		x"24",	--4885
		x"43",	--4886
		x"4e",	--4887
		x"11",	--4888
		x"43",	--4889
		x"10",	--4890
		x"41",	--4891
		x"f0",	--4892
		x"00",	--4893
		x"de",	--4894
		x"4a",	--4895
		x"00",	--4896
		x"40",	--4897
		x"ea",	--4898
		x"41",	--4899
		x"00",	--4900
		x"5a",	--4901
		x"4a",	--4902
		x"5c",	--4903
		x"5c",	--4904
		x"5c",	--4905
		x"4a",	--4906
		x"00",	--4907
		x"50",	--4908
		x"ff",	--4909
		x"00",	--4910
		x"11",	--4911
		x"5e",	--4912
		x"00",	--4913
		x"43",	--4914
		x"00",	--4915
		x"40",	--4916
		x"ea",	--4917
		x"45",	--4918
		x"53",	--4919
		x"45",	--4920
		x"93",	--4921
		x"00",	--4922
		x"20",	--4923
		x"93",	--4924
		x"00",	--4925
		x"27",	--4926
		x"4e",	--4927
		x"00",	--4928
		x"43",	--4929
		x"00",	--4930
		x"41",	--4931
		x"52",	--4932
		x"3c",	--4933
		x"45",	--4934
		x"53",	--4935
		x"45",	--4936
		x"93",	--4937
		x"00",	--4938
		x"24",	--4939
		x"d2",	--4940
		x"00",	--4941
		x"41",	--4942
		x"00",	--4943
		x"4f",	--4944
		x"00",	--4945
		x"3c",	--4946
		x"93",	--4947
		x"00",	--4948
		x"24",	--4949
		x"41",	--4950
		x"00",	--4951
		x"00",	--4952
		x"93",	--4953
		x"20",	--4954
		x"40",	--4955
		x"f0",	--4956
		x"12",	--4957
		x"00",	--4958
		x"12",	--4959
		x"00",	--4960
		x"41",	--4961
		x"00",	--4962
		x"41",	--4963
		x"00",	--4964
		x"12",	--4965
		x"e2",	--4966
		x"52",	--4967
		x"5f",	--4968
		x"00",	--4969
		x"47",	--4970
		x"40",	--4971
		x"ea",	--4972
		x"45",	--4973
		x"53",	--4974
		x"45",	--4975
		x"49",	--4976
		x"00",	--4977
		x"43",	--4978
		x"93",	--4979
		x"20",	--4980
		x"43",	--4981
		x"5e",	--4982
		x"5e",	--4983
		x"5e",	--4984
		x"41",	--4985
		x"f0",	--4986
		x"ff",	--4987
		x"de",	--4988
		x"4a",	--4989
		x"00",	--4990
		x"47",	--4991
		x"40",	--4992
		x"00",	--4993
		x"00",	--4994
		x"3c",	--4995
		x"d3",	--4996
		x"00",	--4997
		x"3c",	--4998
		x"d2",	--4999
		x"00",	--5000
		x"40",	--5001
		x"00",	--5002
		x"00",	--5003
		x"3c",	--5004
		x"40",	--5005
		x"00",	--5006
		x"00",	--5007
		x"41",	--5008
		x"b3",	--5009
		x"24",	--5010
		x"45",	--5011
		x"52",	--5012
		x"45",	--5013
		x"45",	--5014
		x"00",	--5015
		x"45",	--5016
		x"00",	--5017
		x"45",	--5018
		x"00",	--5019
		x"48",	--5020
		x"00",	--5021
		x"47",	--5022
		x"00",	--5023
		x"46",	--5024
		x"00",	--5025
		x"4b",	--5026
		x"00",	--5027
		x"43",	--5028
		x"00",	--5029
		x"93",	--5030
		x"20",	--5031
		x"93",	--5032
		x"20",	--5033
		x"93",	--5034
		x"20",	--5035
		x"93",	--5036
		x"24",	--5037
		x"43",	--5038
		x"00",	--5039
		x"5b",	--5040
		x"43",	--5041
		x"6b",	--5042
		x"4b",	--5043
		x"00",	--5044
		x"4c",	--5045
		x"3c",	--5046
		x"f3",	--5047
		x"45",	--5048
		x"24",	--5049
		x"52",	--5050
		x"45",	--5051
		x"45",	--5052
		x"00",	--5053
		x"48",	--5054
		x"00",	--5055
		x"4b",	--5056
		x"00",	--5057
		x"43",	--5058
		x"00",	--5059
		x"93",	--5060
		x"20",	--5061
		x"3c",	--5062
		x"53",	--5063
		x"45",	--5064
		x"4b",	--5065
		x"00",	--5066
		x"43",	--5067
		x"00",	--5068
		x"93",	--5069
		x"24",	--5070
		x"43",	--5071
		x"00",	--5072
		x"5b",	--5073
		x"43",	--5074
		x"6b",	--5075
		x"4b",	--5076
		x"00",	--5077
		x"47",	--5078
		x"b2",	--5079
		x"00",	--5080
		x"24",	--5081
		x"93",	--5082
		x"00",	--5083
		x"20",	--5084
		x"41",	--5085
		x"90",	--5086
		x"00",	--5087
		x"00",	--5088
		x"20",	--5089
		x"d0",	--5090
		x"00",	--5091
		x"3c",	--5092
		x"92",	--5093
		x"00",	--5094
		x"20",	--5095
		x"d0",	--5096
		x"00",	--5097
		x"48",	--5098
		x"00",	--5099
		x"41",	--5100
		x"b2",	--5101
		x"24",	--5102
		x"93",	--5103
		x"00",	--5104
		x"24",	--5105
		x"40",	--5106
		x"00",	--5107
		x"00",	--5108
		x"b3",	--5109
		x"24",	--5110
		x"e3",	--5111
		x"00",	--5112
		x"e3",	--5113
		x"00",	--5114
		x"e3",	--5115
		x"00",	--5116
		x"e3",	--5117
		x"00",	--5118
		x"53",	--5119
		x"00",	--5120
		x"63",	--5121
		x"00",	--5122
		x"63",	--5123
		x"00",	--5124
		x"63",	--5125
		x"00",	--5126
		x"3c",	--5127
		x"b3",	--5128
		x"24",	--5129
		x"41",	--5130
		x"00",	--5131
		x"41",	--5132
		x"00",	--5133
		x"e3",	--5134
		x"e3",	--5135
		x"4a",	--5136
		x"4b",	--5137
		x"53",	--5138
		x"63",	--5139
		x"4e",	--5140
		x"00",	--5141
		x"4f",	--5142
		x"00",	--5143
		x"3c",	--5144
		x"41",	--5145
		x"00",	--5146
		x"e3",	--5147
		x"53",	--5148
		x"4a",	--5149
		x"00",	--5150
		x"43",	--5151
		x"00",	--5152
		x"b3",	--5153
		x"24",	--5154
		x"41",	--5155
		x"00",	--5156
		x"41",	--5157
		x"00",	--5158
		x"00",	--5159
		x"41",	--5160
		x"00",	--5161
		x"41",	--5162
		x"00",	--5163
		x"41",	--5164
		x"50",	--5165
		x"00",	--5166
		x"46",	--5167
		x"41",	--5168
		x"00",	--5169
		x"00",	--5170
		x"41",	--5171
		x"00",	--5172
		x"10",	--5173
		x"11",	--5174
		x"10",	--5175
		x"11",	--5176
		x"4b",	--5177
		x"00",	--5178
		x"4b",	--5179
		x"00",	--5180
		x"4b",	--5181
		x"00",	--5182
		x"12",	--5183
		x"00",	--5184
		x"12",	--5185
		x"00",	--5186
		x"12",	--5187
		x"00",	--5188
		x"12",	--5189
		x"00",	--5190
		x"49",	--5191
		x"41",	--5192
		x"00",	--5193
		x"48",	--5194
		x"44",	--5195
		x"12",	--5196
		x"ec",	--5197
		x"52",	--5198
		x"4c",	--5199
		x"90",	--5200
		x"00",	--5201
		x"34",	--5202
		x"50",	--5203
		x"00",	--5204
		x"4b",	--5205
		x"00",	--5206
		x"3c",	--5207
		x"4c",	--5208
		x"b3",	--5209
		x"00",	--5210
		x"24",	--5211
		x"40",	--5212
		x"00",	--5213
		x"3c",	--5214
		x"40",	--5215
		x"00",	--5216
		x"5b",	--5217
		x"4a",	--5218
		x"00",	--5219
		x"47",	--5220
		x"53",	--5221
		x"12",	--5222
		x"00",	--5223
		x"12",	--5224
		x"00",	--5225
		x"12",	--5226
		x"00",	--5227
		x"12",	--5228
		x"00",	--5229
		x"49",	--5230
		x"41",	--5231
		x"00",	--5232
		x"48",	--5233
		x"44",	--5234
		x"12",	--5235
		x"ec",	--5236
		x"52",	--5237
		x"4c",	--5238
		x"4d",	--5239
		x"00",	--5240
		x"4e",	--5241
		x"4f",	--5242
		x"53",	--5243
		x"93",	--5244
		x"23",	--5245
		x"93",	--5246
		x"23",	--5247
		x"93",	--5248
		x"23",	--5249
		x"93",	--5250
		x"23",	--5251
		x"43",	--5252
		x"00",	--5253
		x"43",	--5254
		x"00",	--5255
		x"43",	--5256
		x"00",	--5257
		x"43",	--5258
		x"00",	--5259
		x"3c",	--5260
		x"b3",	--5261
		x"24",	--5262
		x"41",	--5263
		x"00",	--5264
		x"41",	--5265
		x"00",	--5266
		x"41",	--5267
		x"50",	--5268
		x"00",	--5269
		x"41",	--5270
		x"00",	--5271
		x"10",	--5272
		x"11",	--5273
		x"10",	--5274
		x"11",	--5275
		x"41",	--5276
		x"00",	--5277
		x"49",	--5278
		x"44",	--5279
		x"47",	--5280
		x"12",	--5281
		x"eb",	--5282
		x"4e",	--5283
		x"90",	--5284
		x"00",	--5285
		x"34",	--5286
		x"50",	--5287
		x"00",	--5288
		x"4b",	--5289
		x"00",	--5290
		x"3c",	--5291
		x"4e",	--5292
		x"b3",	--5293
		x"00",	--5294
		x"24",	--5295
		x"40",	--5296
		x"00",	--5297
		x"3c",	--5298
		x"40",	--5299
		x"00",	--5300
		x"5b",	--5301
		x"4a",	--5302
		x"00",	--5303
		x"48",	--5304
		x"53",	--5305
		x"41",	--5306
		x"00",	--5307
		x"49",	--5308
		x"44",	--5309
		x"47",	--5310
		x"12",	--5311
		x"eb",	--5312
		x"4e",	--5313
		x"4f",	--5314
		x"53",	--5315
		x"93",	--5316
		x"23",	--5317
		x"93",	--5318
		x"23",	--5319
		x"43",	--5320
		x"00",	--5321
		x"43",	--5322
		x"00",	--5323
		x"3c",	--5324
		x"41",	--5325
		x"00",	--5326
		x"41",	--5327
		x"50",	--5328
		x"00",	--5329
		x"41",	--5330
		x"00",	--5331
		x"47",	--5332
		x"12",	--5333
		x"eb",	--5334
		x"4f",	--5335
		x"90",	--5336
		x"00",	--5337
		x"34",	--5338
		x"50",	--5339
		x"00",	--5340
		x"4d",	--5341
		x"00",	--5342
		x"3c",	--5343
		x"4f",	--5344
		x"b3",	--5345
		x"00",	--5346
		x"24",	--5347
		x"40",	--5348
		x"00",	--5349
		x"3c",	--5350
		x"40",	--5351
		x"00",	--5352
		x"5d",	--5353
		x"4c",	--5354
		x"00",	--5355
		x"48",	--5356
		x"53",	--5357
		x"41",	--5358
		x"00",	--5359
		x"47",	--5360
		x"12",	--5361
		x"eb",	--5362
		x"4f",	--5363
		x"53",	--5364
		x"93",	--5365
		x"23",	--5366
		x"43",	--5367
		x"00",	--5368
		x"90",	--5369
		x"00",	--5370
		x"00",	--5371
		x"24",	--5372
		x"43",	--5373
		x"00",	--5374
		x"93",	--5375
		x"00",	--5376
		x"24",	--5377
		x"41",	--5378
		x"50",	--5379
		x"00",	--5380
		x"4f",	--5381
		x"00",	--5382
		x"41",	--5383
		x"00",	--5384
		x"10",	--5385
		x"11",	--5386
		x"10",	--5387
		x"11",	--5388
		x"4a",	--5389
		x"00",	--5390
		x"46",	--5391
		x"00",	--5392
		x"46",	--5393
		x"10",	--5394
		x"11",	--5395
		x"10",	--5396
		x"11",	--5397
		x"4a",	--5398
		x"00",	--5399
		x"41",	--5400
		x"00",	--5401
		x"41",	--5402
		x"00",	--5403
		x"81",	--5404
		x"00",	--5405
		x"71",	--5406
		x"00",	--5407
		x"83",	--5408
		x"91",	--5409
		x"00",	--5410
		x"2c",	--5411
		x"d3",	--5412
		x"00",	--5413
		x"41",	--5414
		x"00",	--5415
		x"8c",	--5416
		x"4e",	--5417
		x"00",	--5418
		x"3c",	--5419
		x"93",	--5420
		x"00",	--5421
		x"24",	--5422
		x"41",	--5423
		x"00",	--5424
		x"00",	--5425
		x"12",	--5426
		x"00",	--5427
		x"12",	--5428
		x"00",	--5429
		x"41",	--5430
		x"00",	--5431
		x"46",	--5432
		x"53",	--5433
		x"41",	--5434
		x"00",	--5435
		x"12",	--5436
		x"e2",	--5437
		x"52",	--5438
		x"5f",	--5439
		x"00",	--5440
		x"3c",	--5441
		x"49",	--5442
		x"11",	--5443
		x"12",	--5444
		x"00",	--5445
		x"49",	--5446
		x"58",	--5447
		x"91",	--5448
		x"00",	--5449
		x"2b",	--5450
		x"49",	--5451
		x"00",	--5452
		x"4e",	--5453
		x"00",	--5454
		x"43",	--5455
		x"3c",	--5456
		x"41",	--5457
		x"00",	--5458
		x"00",	--5459
		x"43",	--5460
		x"00",	--5461
		x"43",	--5462
		x"00",	--5463
		x"3c",	--5464
		x"4e",	--5465
		x"43",	--5466
		x"00",	--5467
		x"43",	--5468
		x"00",	--5469
		x"43",	--5470
		x"41",	--5471
		x"00",	--5472
		x"46",	--5473
		x"93",	--5474
		x"24",	--5475
		x"40",	--5476
		x"e4",	--5477
		x"41",	--5478
		x"00",	--5479
		x"50",	--5480
		x"00",	--5481
		x"41",	--5482
		x"41",	--5483
		x"41",	--5484
		x"41",	--5485
		x"41",	--5486
		x"41",	--5487
		x"41",	--5488
		x"41",	--5489
		x"41",	--5490
		x"43",	--5491
		x"93",	--5492
		x"34",	--5493
		x"40",	--5494
		x"00",	--5495
		x"e3",	--5496
		x"53",	--5497
		x"93",	--5498
		x"34",	--5499
		x"e3",	--5500
		x"e3",	--5501
		x"53",	--5502
		x"12",	--5503
		x"12",	--5504
		x"eb",	--5505
		x"41",	--5506
		x"b3",	--5507
		x"24",	--5508
		x"e3",	--5509
		x"53",	--5510
		x"b3",	--5511
		x"24",	--5512
		x"e3",	--5513
		x"53",	--5514
		x"41",	--5515
		x"12",	--5516
		x"ea",	--5517
		x"4e",	--5518
		x"41",	--5519
		x"12",	--5520
		x"12",	--5521
		x"12",	--5522
		x"40",	--5523
		x"00",	--5524
		x"4c",	--5525
		x"4d",	--5526
		x"43",	--5527
		x"43",	--5528
		x"5e",	--5529
		x"6f",	--5530
		x"6c",	--5531
		x"6d",	--5532
		x"9b",	--5533
		x"28",	--5534
		x"20",	--5535
		x"9a",	--5536
		x"28",	--5537
		x"8a",	--5538
		x"7b",	--5539
		x"d3",	--5540
		x"83",	--5541
		x"23",	--5542
		x"41",	--5543
		x"41",	--5544
		x"41",	--5545
		x"41",	--5546
		x"12",	--5547
		x"eb",	--5548
		x"4c",	--5549
		x"4d",	--5550
		x"41",	--5551
		x"12",	--5552
		x"43",	--5553
		x"93",	--5554
		x"34",	--5555
		x"40",	--5556
		x"00",	--5557
		x"e3",	--5558
		x"e3",	--5559
		x"53",	--5560
		x"63",	--5561
		x"93",	--5562
		x"34",	--5563
		x"e3",	--5564
		x"e3",	--5565
		x"e3",	--5566
		x"53",	--5567
		x"63",	--5568
		x"12",	--5569
		x"eb",	--5570
		x"b3",	--5571
		x"24",	--5572
		x"e3",	--5573
		x"e3",	--5574
		x"53",	--5575
		x"63",	--5576
		x"b3",	--5577
		x"24",	--5578
		x"e3",	--5579
		x"e3",	--5580
		x"53",	--5581
		x"63",	--5582
		x"41",	--5583
		x"41",	--5584
		x"12",	--5585
		x"eb",	--5586
		x"4c",	--5587
		x"4d",	--5588
		x"41",	--5589
		x"40",	--5590
		x"00",	--5591
		x"4e",	--5592
		x"43",	--5593
		x"5f",	--5594
		x"6e",	--5595
		x"9d",	--5596
		x"28",	--5597
		x"8d",	--5598
		x"d3",	--5599
		x"83",	--5600
		x"23",	--5601
		x"41",	--5602
		x"12",	--5603
		x"eb",	--5604
		x"4e",	--5605
		x"41",	--5606
		x"12",	--5607
		x"12",	--5608
		x"12",	--5609
		x"12",	--5610
		x"12",	--5611
		x"00",	--5612
		x"48",	--5613
		x"49",	--5614
		x"4a",	--5615
		x"4b",	--5616
		x"43",	--5617
		x"43",	--5618
		x"43",	--5619
		x"43",	--5620
		x"5c",	--5621
		x"6d",	--5622
		x"6e",	--5623
		x"6f",	--5624
		x"68",	--5625
		x"69",	--5626
		x"6a",	--5627
		x"6b",	--5628
		x"97",	--5629
		x"28",	--5630
		x"20",	--5631
		x"96",	--5632
		x"28",	--5633
		x"20",	--5634
		x"95",	--5635
		x"28",	--5636
		x"20",	--5637
		x"94",	--5638
		x"28",	--5639
		x"84",	--5640
		x"75",	--5641
		x"76",	--5642
		x"77",	--5643
		x"d3",	--5644
		x"83",	--5645
		x"00",	--5646
		x"23",	--5647
		x"53",	--5648
		x"41",	--5649
		x"41",	--5650
		x"41",	--5651
		x"41",	--5652
		x"41",	--5653
		x"12",	--5654
		x"12",	--5655
		x"12",	--5656
		x"12",	--5657
		x"41",	--5658
		x"00",	--5659
		x"41",	--5660
		x"00",	--5661
		x"41",	--5662
		x"00",	--5663
		x"41",	--5664
		x"00",	--5665
		x"12",	--5666
		x"eb",	--5667
		x"41",	--5668
		x"41",	--5669
		x"41",	--5670
		x"41",	--5671
		x"41",	--5672
		x"12",	--5673
		x"12",	--5674
		x"12",	--5675
		x"12",	--5676
		x"41",	--5677
		x"00",	--5678
		x"41",	--5679
		x"00",	--5680
		x"41",	--5681
		x"00",	--5682
		x"41",	--5683
		x"00",	--5684
		x"12",	--5685
		x"eb",	--5686
		x"48",	--5687
		x"49",	--5688
		x"4a",	--5689
		x"4b",	--5690
		x"41",	--5691
		x"41",	--5692
		x"41",	--5693
		x"41",	--5694
		x"41",	--5695
		x"12",	--5696
		x"12",	--5697
		x"12",	--5698
		x"12",	--5699
		x"12",	--5700
		x"41",	--5701
		x"00",	--5702
		x"41",	--5703
		x"00",	--5704
		x"41",	--5705
		x"00",	--5706
		x"41",	--5707
		x"00",	--5708
		x"12",	--5709
		x"eb",	--5710
		x"41",	--5711
		x"00",	--5712
		x"48",	--5713
		x"00",	--5714
		x"49",	--5715
		x"00",	--5716
		x"4a",	--5717
		x"00",	--5718
		x"4b",	--5719
		x"00",	--5720
		x"41",	--5721
		x"41",	--5722
		x"41",	--5723
		x"41",	--5724
		x"41",	--5725
		x"41",	--5726
		x"13",	--5727
		x"d0",	--5728
		x"00",	--5729
		x"3f",	--5730
		x"74",	--5731
		x"70",	--5732
		x"0a",	--5733
		x"63",	--5734
		x"72",	--5735
		x"65",	--5736
		x"74",	--5737
		x"75",	--5738
		x"61",	--5739
		x"65",	--5740
		x"0d",	--5741
		x"00",	--5742
		x"25",	--5743
		x"20",	--5744
		x"45",	--5745
		x"54",	--5746
		x"52",	--5747
		x"47",	--5748
		x"54",	--5749
		x"3c",	--5750
		x"49",	--5751
		x"45",	--5752
		x"55",	--5753
		x"3e",	--5754
		x"0a",	--5755
		x"25",	--5756
		x"20",	--5757
		x"64",	--5758
		x"0a",	--5759
		x"4e",	--5760
		x"74",	--5761
		x"69",	--5762
		x"70",	--5763
		x"65",	--5764
		x"65",	--5765
		x"74",	--5766
		x"64",	--5767
		x"59",	--5768
		x"74",	--5769
		x"0a",	--5770
		x"57",	--5771
		x"69",	--5772
		x"69",	--5773
		x"67",	--5774
		x"66",	--5775
		x"72",	--5776
		x"61",	--5777
		x"6e",	--5778
		x"77",	--5779
		x"2e",	--5780
		x"69",	--5781
		x"20",	--5782
		x"69",	--5783
		x"65",	--5784
		x"0a",	--5785
		x"57",	--5786
		x"20",	--5787
		x"68",	--5788
		x"75",	--5789
		x"64",	--5790
		x"6e",	--5791
		x"74",	--5792
		x"73",	--5793
		x"65",	--5794
		x"74",	--5795
		x"61",	--5796
		x"0d",	--5797
		x"00",	--5798
		x"74",	--5799
		x"70",	--5800
		x"0a",	--5801
		x"65",	--5802
		x"72",	--5803
		x"72",	--5804
		x"20",	--5805
		x"69",	--5806
		x"73",	--5807
		x"6e",	--5808
		x"20",	--5809
		x"72",	--5810
		x"75",	--5811
		x"65",	--5812
		x"74",	--5813
		x"0a",	--5814
		x"63",	--5815
		x"72",	--5816
		x"65",	--5817
		x"74",	--5818
		x"75",	--5819
		x"61",	--5820
		x"65",	--5821
		x"0d",	--5822
		x"00",	--5823
		x"25",	--5824
		x"20",	--5825
		x"45",	--5826
		x"54",	--5827
		x"52",	--5828
		x"47",	--5829
		x"54",	--5830
		x"3c",	--5831
		x"49",	--5832
		x"45",	--5833
		x"55",	--5834
		x"3e",	--5835
		x"0a",	--5836
		x"25",	--5837
		x"20",	--5838
		x"64",	--5839
		x"0a",	--5840
		x"25",	--5841
		x"64",	--5842
		x"25",	--5843
		x"64",	--5844
		x"25",	--5845
		x"0d",	--5846
		x"00",	--5847
		x"64",	--5848
		x"25",	--5849
		x"0d",	--5850
		x"00",	--5851
		x"c9",	--5852
		x"c9",	--5853
		x"c9",	--5854
		x"c9",	--5855
		x"c9",	--5856
		x"c9",	--5857
		x"c9",	--5858
		x"c9",	--5859
		x"0a",	--5860
		x"3d",	--5861
		x"3d",	--5862
		x"3d",	--5863
		x"4d",	--5864
		x"72",	--5865
		x"65",	--5866
		x"20",	--5867
		x"43",	--5868
		x"20",	--5869
		x"3d",	--5870
		x"3d",	--5871
		x"3d",	--5872
		x"0a",	--5873
		x"69",	--5874
		x"74",	--5875
		x"72",	--5876
		x"63",	--5877
		x"69",	--5878
		x"65",	--5879
		x"6d",	--5880
		x"64",	--5881
		x"00",	--5882
		x"72",	--5883
		x"74",	--5884
		x"00",	--5885
		x"65",	--5886
		x"64",	--5887
		x"62",	--5888
		x"7a",	--5889
		x"65",	--5890
		x"00",	--5891
		x"77",	--5892
		x"00",	--5893
		x"6e",	--5894
		x"6f",	--5895
		x"65",	--5896
		x"00",	--5897
		x"70",	--5898
		x"65",	--5899
		x"20",	--5900
		x"6f",	--5901
		x"74",	--5902
		x"6f",	--5903
		x"6c",	--5904
		x"72",	--5905
		x"73",	--5906
		x"65",	--5907
		x"64",	--5908
		x"63",	--5909
		x"6e",	--5910
		x"69",	--5911
		x"75",	--5912
		x"61",	--5913
		x"69",	--5914
		x"6e",	--5915
		x"62",	--5916
		x"6f",	--5917
		x"6c",	--5918
		x"61",	--5919
		x"65",	--5920
		x"00",	--5921
		x"0a",	--5922
		x"08",	--5923
		x"08",	--5924
		x"25",	--5925
		x"00",	--5926
		x"50",	--5927
		x"0a",	--5928
		x"44",	--5929
		x"57",	--5930
		x"0d",	--5931
		x"00",	--5932
		x"49",	--5933
		x"48",	--5934
		x"0d",	--5935
		x"00",	--5936
		x"45",	--5937
		x"54",	--5938
		x"0a",	--5939
		x"00",	--5940
		x"72",	--5941
		x"74",	--5942
		x"0a",	--5943
		x"00",	--5944
		x"72",	--5945
		x"6f",	--5946
		x"3a",	--5947
		x"6d",	--5948
		x"73",	--5949
		x"69",	--5950
		x"67",	--5951
		x"61",	--5952
		x"67",	--5953
		x"6d",	--5954
		x"6e",	--5955
		x"0d",	--5956
		x"00",	--5957
		x"6f",	--5958
		x"72",	--5959
		x"63",	--5960
		x"20",	--5961
		x"73",	--5962
		x"67",	--5963
		x"3a",	--5964
		x"0a",	--5965
		x"09",	--5966
		x"73",	--5967
		x"52",	--5968
		x"47",	--5969
		x"53",	--5970
		x"45",	--5971
		x"20",	--5972
		x"41",	--5973
		x"55",	--5974
		x"0d",	--5975
		x"00",	--5976
		x"3d",	--5977
		x"64",	--5978
		x"76",	--5979
		x"25",	--5980
		x"0d",	--5981
		x"00",	--5982
		x"25",	--5983
		x"20",	--5984
		x"45",	--5985
		x"49",	--5986
		x"54",	--5987
		x"52",	--5988
		x"0a",	--5989
		x"72",	--5990
		x"61",	--5991
		x"0a",	--5992
		x"00",	--5993
		x"63",	--5994
		x"69",	--5995
		x"20",	--5996
		x"6f",	--5997
		x"20",	--5998
		x"20",	--5999
		x"75",	--6000
		x"62",	--6001
		x"72",	--6002
		x"0a",	--6003
		x"25",	--6004
		x"20",	--6005
		x"73",	--6006
		x"0a",	--6007
		x"25",	--6008
		x"3a",	--6009
		x"6e",	--6010
		x"20",	--6011
		x"75",	--6012
		x"68",	--6013
		x"63",	--6014
		x"6d",	--6015
		x"61",	--6016
		x"64",	--6017
		x"0a",	--6018
		x"00",	--6019
		x"d3",	--6020
		x"d2",	--6021
		x"d2",	--6022
		x"d2",	--6023
		x"d2",	--6024
		x"d2",	--6025
		x"d2",	--6026
		x"d2",	--6027
		x"d2",	--6028
		x"d2",	--6029
		x"d2",	--6030
		x"d2",	--6031
		x"d2",	--6032
		x"d2",	--6033
		x"d2",	--6034
		x"d2",	--6035
		x"d2",	--6036
		x"d2",	--6037
		x"d2",	--6038
		x"d2",	--6039
		x"d2",	--6040
		x"d2",	--6041
		x"d2",	--6042
		x"d2",	--6043
		x"d2",	--6044
		x"d2",	--6045
		x"d2",	--6046
		x"d2",	--6047
		x"d2",	--6048
		x"d3",	--6049
		x"d2",	--6050
		x"d2",	--6051
		x"d2",	--6052
		x"d2",	--6053
		x"d2",	--6054
		x"d2",	--6055
		x"d2",	--6056
		x"d2",	--6057
		x"d2",	--6058
		x"d2",	--6059
		x"d2",	--6060
		x"d2",	--6061
		x"d2",	--6062
		x"d2",	--6063
		x"d2",	--6064
		x"d2",	--6065
		x"d2",	--6066
		x"d2",	--6067
		x"d2",	--6068
		x"d2",	--6069
		x"d2",	--6070
		x"d2",	--6071
		x"d2",	--6072
		x"d2",	--6073
		x"d2",	--6074
		x"d2",	--6075
		x"d2",	--6076
		x"d2",	--6077
		x"d2",	--6078
		x"d2",	--6079
		x"d2",	--6080
		x"d3",	--6081
		x"d3",	--6082
		x"d2",	--6083
		x"d2",	--6084
		x"d2",	--6085
		x"d2",	--6086
		x"d2",	--6087
		x"d2",	--6088
		x"d2",	--6089
		x"d2",	--6090
		x"d2",	--6091
		x"d2",	--6092
		x"d2",	--6093
		x"d2",	--6094
		x"d2",	--6095
		x"d2",	--6096
		x"d2",	--6097
		x"d2",	--6098
		x"d2",	--6099
		x"d2",	--6100
		x"d2",	--6101
		x"d2",	--6102
		x"d2",	--6103
		x"31",	--6104
		x"33",	--6105
		x"35",	--6106
		x"37",	--6107
		x"39",	--6108
		x"62",	--6109
		x"64",	--6110
		x"66",	--6111
		x"00",	--6112
		x"00",	--6113
		x"00",	--6114
		x"00",	--6115
		x"00",	--6116
		x"01",	--6117
		x"02",	--6118
		x"03",	--6119
		x"03",	--6120
		x"04",	--6121
		x"04",	--6122
		x"04",	--6123
		x"04",	--6124
		x"05",	--6125
		x"05",	--6126
		x"05",	--6127
		x"05",	--6128
		x"05",	--6129
		x"05",	--6130
		x"05",	--6131
		x"05",	--6132
		x"06",	--6133
		x"06",	--6134
		x"06",	--6135
		x"06",	--6136
		x"06",	--6137
		x"06",	--6138
		x"06",	--6139
		x"06",	--6140
		x"06",	--6141
		x"06",	--6142
		x"06",	--6143
		x"06",	--6144
		x"06",	--6145
		x"06",	--6146
		x"06",	--6147
		x"06",	--6148
		x"07",	--6149
		x"07",	--6150
		x"07",	--6151
		x"07",	--6152
		x"07",	--6153
		x"07",	--6154
		x"07",	--6155
		x"07",	--6156
		x"07",	--6157
		x"07",	--6158
		x"07",	--6159
		x"07",	--6160
		x"07",	--6161
		x"07",	--6162
		x"07",	--6163
		x"07",	--6164
		x"07",	--6165
		x"07",	--6166
		x"07",	--6167
		x"07",	--6168
		x"07",	--6169
		x"07",	--6170
		x"07",	--6171
		x"07",	--6172
		x"07",	--6173
		x"07",	--6174
		x"07",	--6175
		x"07",	--6176
		x"07",	--6177
		x"07",	--6178
		x"07",	--6179
		x"07",	--6180
		x"08",	--6181
		x"08",	--6182
		x"08",	--6183
		x"08",	--6184
		x"08",	--6185
		x"08",	--6186
		x"08",	--6187
		x"08",	--6188
		x"08",	--6189
		x"08",	--6190
		x"08",	--6191
		x"08",	--6192
		x"08",	--6193
		x"08",	--6194
		x"08",	--6195
		x"08",	--6196
		x"08",	--6197
		x"08",	--6198
		x"08",	--6199
		x"08",	--6200
		x"08",	--6201
		x"08",	--6202
		x"08",	--6203
		x"08",	--6204
		x"08",	--6205
		x"08",	--6206
		x"08",	--6207
		x"08",	--6208
		x"08",	--6209
		x"08",	--6210
		x"08",	--6211
		x"08",	--6212
		x"08",	--6213
		x"08",	--6214
		x"08",	--6215
		x"08",	--6216
		x"08",	--6217
		x"08",	--6218
		x"08",	--6219
		x"08",	--6220
		x"08",	--6221
		x"08",	--6222
		x"08",	--6223
		x"08",	--6224
		x"08",	--6225
		x"08",	--6226
		x"08",	--6227
		x"08",	--6228
		x"08",	--6229
		x"08",	--6230
		x"08",	--6231
		x"08",	--6232
		x"08",	--6233
		x"08",	--6234
		x"08",	--6235
		x"08",	--6236
		x"08",	--6237
		x"08",	--6238
		x"08",	--6239
		x"08",	--6240
		x"08",	--6241
		x"08",	--6242
		x"08",	--6243
		x"08",	--6244
		x"6e",	--6245
		x"6c",	--6246
		x"29",	--6247
		x"00",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"65",	--6252
		x"70",	--6253
		x"00",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"c3",	--8176
		x"c3",	--8177
		x"c3",	--8178
		x"c3",	--8179
		x"c3",	--8180
		x"c3",	--8181
		x"c3",	--8182
		x"d3",	--8183
		x"cf",	--8184
		x"c3",	--8185
		x"c3",	--8186
		x"c3",	--8187
		x"c3",	--8188
		x"c3",	--8189
		x"c3",	--8190
		x"c0");	--8191

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
