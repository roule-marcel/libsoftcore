library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package log2_pkg is
	function log2ceil (n : natural) return natural;
end package log2_pkg;
