library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"5c",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"08",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"5c",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"d0",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"54",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"5c",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"08",	--29
		x"f9",	--30
		x"31",	--31
		x"be",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"80",	--41
		x"0f",	--42
		x"b0",	--43
		x"7a",	--44
		x"b0",	--45
		x"74",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"26",	--50
		x"b0",	--51
		x"3e",	--52
		x"21",	--53
		x"3d",	--54
		x"43",	--55
		x"3e",	--56
		x"ac",	--57
		x"7f",	--58
		x"77",	--59
		x"b0",	--60
		x"a4",	--61
		x"3d",	--62
		x"49",	--63
		x"3e",	--64
		x"20",	--65
		x"7f",	--66
		x"72",	--67
		x"b0",	--68
		x"a4",	--69
		x"3d",	--70
		x"4e",	--71
		x"3e",	--72
		x"fc",	--73
		x"7f",	--74
		x"70",	--75
		x"b0",	--76
		x"a4",	--77
		x"3d",	--78
		x"52",	--79
		x"3e",	--80
		x"cc",	--81
		x"7f",	--82
		x"65",	--83
		x"b0",	--84
		x"a4",	--85
		x"3d",	--86
		x"5a",	--87
		x"3e",	--88
		x"c6",	--89
		x"7f",	--90
		x"62",	--91
		x"b0",	--92
		x"a4",	--93
		x"0e",	--94
		x"0f",	--95
		x"b0",	--96
		x"3a",	--97
		x"2c",	--98
		x"3d",	--99
		x"20",	--100
		x"3e",	--101
		x"80",	--102
		x"0f",	--103
		x"3f",	--104
		x"0e",	--105
		x"b0",	--106
		x"4a",	--107
		x"0f",	--108
		x"3f",	--109
		x"0e",	--110
		x"b0",	--111
		x"92",	--112
		x"2c",	--113
		x"3d",	--114
		x"20",	--115
		x"3e",	--116
		x"88",	--117
		x"0f",	--118
		x"2f",	--119
		x"b0",	--120
		x"4a",	--121
		x"0f",	--122
		x"2f",	--123
		x"b0",	--124
		x"92",	--125
		x"0e",	--126
		x"2e",	--127
		x"0f",	--128
		x"3f",	--129
		x"0e",	--130
		x"b0",	--131
		x"f2",	--132
		x"3e",	--133
		x"98",	--134
		x"0f",	--135
		x"2f",	--136
		x"b0",	--137
		x"54",	--138
		x"3e",	--139
		x"9c",	--140
		x"0f",	--141
		x"b0",	--142
		x"54",	--143
		x"0e",	--144
		x"0f",	--145
		x"2f",	--146
		x"b0",	--147
		x"c2",	--148
		x"b0",	--149
		x"70",	--150
		x"0e",	--151
		x"3f",	--152
		x"38",	--153
		x"b0",	--154
		x"80",	--155
		x"1e",	--156
		x"b0",	--157
		x"be",	--158
		x"f2",	--159
		x"80",	--160
		x"19",	--161
		x"32",	--162
		x"0b",	--163
		x"b0",	--164
		x"88",	--165
		x"0f",	--166
		x"fc",	--167
		x"b0",	--168
		x"b0",	--169
		x"7f",	--170
		x"15",	--171
		x"7f",	--172
		x"0d",	--173
		x"1b",	--174
		x"30",	--175
		x"65",	--176
		x"b0",	--177
		x"3e",	--178
		x"21",	--179
		x"3f",	--180
		x"18",	--181
		x"0f",	--182
		x"0b",	--183
		x"cb",	--184
		x"00",	--185
		x"0e",	--186
		x"5f",	--187
		x"18",	--188
		x"b0",	--189
		x"d8",	--190
		x"0b",	--191
		x"e3",	--192
		x"0b",	--193
		x"e1",	--194
		x"3b",	--195
		x"30",	--196
		x"68",	--197
		x"b0",	--198
		x"3e",	--199
		x"21",	--200
		x"da",	--201
		x"3b",	--202
		x"28",	--203
		x"d7",	--204
		x"4e",	--205
		x"8e",	--206
		x"0e",	--207
		x"30",	--208
		x"6c",	--209
		x"81",	--210
		x"44",	--211
		x"b0",	--212
		x"3e",	--213
		x"21",	--214
		x"3e",	--215
		x"18",	--216
		x"0e",	--217
		x"0e",	--218
		x"1f",	--219
		x"40",	--220
		x"ce",	--221
		x"00",	--222
		x"1b",	--223
		x"c3",	--224
		x"30",	--225
		x"84",	--226
		x"b2",	--227
		x"00",	--228
		x"92",	--229
		x"a2",	--230
		x"94",	--231
		x"b2",	--232
		x"6d",	--233
		x"96",	--234
		x"30",	--235
		x"8c",	--236
		x"b0",	--237
		x"3e",	--238
		x"92",	--239
		x"90",	--240
		x"b1",	--241
		x"aa",	--242
		x"00",	--243
		x"b0",	--244
		x"3e",	--245
		x"21",	--246
		x"0f",	--247
		x"30",	--248
		x"82",	--249
		x"16",	--250
		x"82",	--251
		x"14",	--252
		x"30",	--253
		x"0b",	--254
		x"0a",	--255
		x"21",	--256
		x"0b",	--257
		x"2f",	--258
		x"38",	--259
		x"37",	--260
		x"0e",	--261
		x"1f",	--262
		x"02",	--263
		x"b0",	--264
		x"7c",	--265
		x"0a",	--266
		x"0e",	--267
		x"1f",	--268
		x"04",	--269
		x"b0",	--270
		x"7c",	--271
		x"0b",	--272
		x"0f",	--273
		x"0a",	--274
		x"30",	--275
		x"ff",	--276
		x"b0",	--277
		x"3e",	--278
		x"31",	--279
		x"06",	--280
		x"0e",	--281
		x"0f",	--282
		x"b0",	--283
		x"a2",	--284
		x"0c",	--285
		x"3d",	--286
		x"c8",	--287
		x"b0",	--288
		x"72",	--289
		x"0d",	--290
		x"0e",	--291
		x"1f",	--292
		x"16",	--293
		x"b0",	--294
		x"e6",	--295
		x"0e",	--296
		x"0f",	--297
		x"b0",	--298
		x"a2",	--299
		x"0c",	--300
		x"3d",	--301
		x"c8",	--302
		x"b0",	--303
		x"72",	--304
		x"0d",	--305
		x"0e",	--306
		x"1f",	--307
		x"14",	--308
		x"b0",	--309
		x"e6",	--310
		x"0f",	--311
		x"21",	--312
		x"3a",	--313
		x"3b",	--314
		x"30",	--315
		x"30",	--316
		x"c3",	--317
		x"b0",	--318
		x"3e",	--319
		x"b1",	--320
		x"dd",	--321
		x"00",	--322
		x"b0",	--323
		x"3e",	--324
		x"a1",	--325
		x"00",	--326
		x"30",	--327
		x"ee",	--328
		x"b0",	--329
		x"3e",	--330
		x"21",	--331
		x"3f",	--332
		x"ea",	--333
		x"1f",	--334
		x"1a",	--335
		x"2e",	--336
		x"1f",	--337
		x"18",	--338
		x"2f",	--339
		x"2e",	--340
		x"1e",	--341
		x"02",	--342
		x"2f",	--343
		x"1f",	--344
		x"02",	--345
		x"30",	--346
		x"07",	--347
		x"b0",	--348
		x"3e",	--349
		x"31",	--350
		x"0a",	--351
		x"30",	--352
		x"82",	--353
		x"18",	--354
		x"82",	--355
		x"1a",	--356
		x"30",	--357
		x"0b",	--358
		x"21",	--359
		x"0b",	--360
		x"81",	--361
		x"00",	--362
		x"1f",	--363
		x"13",	--364
		x"b2",	--365
		x"00",	--366
		x"24",	--367
		x"92",	--368
		x"08",	--369
		x"0e",	--370
		x"1f",	--371
		x"02",	--372
		x"b0",	--373
		x"7c",	--374
		x"0e",	--375
		x"1f",	--376
		x"00",	--377
		x"b0",	--378
		x"be",	--379
		x"0f",	--380
		x"21",	--381
		x"3b",	--382
		x"30",	--383
		x"82",	--384
		x"08",	--385
		x"0a",	--386
		x"82",	--387
		x"08",	--388
		x"1f",	--389
		x"00",	--390
		x"b0",	--391
		x"dc",	--392
		x"0f",	--393
		x"21",	--394
		x"3b",	--395
		x"30",	--396
		x"0f",	--397
		x"b0",	--398
		x"9c",	--399
		x"0f",	--400
		x"21",	--401
		x"3b",	--402
		x"30",	--403
		x"0e",	--404
		x"3f",	--405
		x"9c",	--406
		x"b0",	--407
		x"80",	--408
		x"82",	--409
		x"00",	--410
		x"d4",	--411
		x"1e",	--412
		x"0a",	--413
		x"3e",	--414
		x"06",	--415
		x"0f",	--416
		x"0f",	--417
		x"10",	--418
		x"16",	--419
		x"c2",	--420
		x"19",	--421
		x"3e",	--422
		x"07",	--423
		x"03",	--424
		x"82",	--425
		x"0a",	--426
		x"30",	--427
		x"1e",	--428
		x"82",	--429
		x"0a",	--430
		x"30",	--431
		x"f2",	--432
		x"0e",	--433
		x"19",	--434
		x"f2",	--435
		x"f2",	--436
		x"0a",	--437
		x"19",	--438
		x"ee",	--439
		x"e2",	--440
		x"19",	--441
		x"eb",	--442
		x"f2",	--443
		x"0d",	--444
		x"19",	--445
		x"e7",	--446
		x"f2",	--447
		x"09",	--448
		x"19",	--449
		x"e3",	--450
		x"f2",	--451
		x"03",	--452
		x"19",	--453
		x"df",	--454
		x"f2",	--455
		x"07",	--456
		x"19",	--457
		x"db",	--458
		x"5e",	--459
		x"19",	--460
		x"4e",	--461
		x"0f",	--462
		x"03",	--463
		x"c2",	--464
		x"19",	--465
		x"30",	--466
		x"c2",	--467
		x"19",	--468
		x"30",	--469
		x"0b",	--470
		x"0a",	--471
		x"21",	--472
		x"0a",	--473
		x"0b",	--474
		x"30",	--475
		x"70",	--476
		x"b0",	--477
		x"3e",	--478
		x"21",	--479
		x"3a",	--480
		x"03",	--481
		x"1b",	--482
		x"0e",	--483
		x"1f",	--484
		x"02",	--485
		x"b0",	--486
		x"7c",	--487
		x"0a",	--488
		x"0e",	--489
		x"1f",	--490
		x"04",	--491
		x"b0",	--492
		x"7c",	--493
		x"0b",	--494
		x"0f",	--495
		x"0a",	--496
		x"30",	--497
		x"b8",	--498
		x"b0",	--499
		x"3e",	--500
		x"31",	--501
		x"06",	--502
		x"8a",	--503
		x"00",	--504
		x"0f",	--505
		x"21",	--506
		x"3a",	--507
		x"3b",	--508
		x"30",	--509
		x"30",	--510
		x"78",	--511
		x"b0",	--512
		x"3e",	--513
		x"b1",	--514
		x"92",	--515
		x"00",	--516
		x"b0",	--517
		x"3e",	--518
		x"a1",	--519
		x"00",	--520
		x"30",	--521
		x"a3",	--522
		x"b0",	--523
		x"3e",	--524
		x"21",	--525
		x"3f",	--526
		x"ea",	--527
		x"0b",	--528
		x"21",	--529
		x"0b",	--530
		x"1f",	--531
		x"17",	--532
		x"16",	--533
		x"30",	--534
		x"d3",	--535
		x"b0",	--536
		x"3e",	--537
		x"21",	--538
		x"0e",	--539
		x"1f",	--540
		x"02",	--541
		x"b0",	--542
		x"7c",	--543
		x"2f",	--544
		x"0f",	--545
		x"30",	--546
		x"b8",	--547
		x"b0",	--548
		x"3e",	--549
		x"31",	--550
		x"06",	--551
		x"0f",	--552
		x"21",	--553
		x"3b",	--554
		x"30",	--555
		x"30",	--556
		x"78",	--557
		x"b0",	--558
		x"3e",	--559
		x"b1",	--560
		x"92",	--561
		x"00",	--562
		x"b0",	--563
		x"3e",	--564
		x"a1",	--565
		x"00",	--566
		x"30",	--567
		x"c4",	--568
		x"b0",	--569
		x"3e",	--570
		x"21",	--571
		x"3f",	--572
		x"eb",	--573
		x"0b",	--574
		x"0a",	--575
		x"8e",	--576
		x"00",	--577
		x"6d",	--578
		x"4d",	--579
		x"5e",	--580
		x"1f",	--581
		x"0a",	--582
		x"0c",	--583
		x"0f",	--584
		x"7b",	--585
		x"0a",	--586
		x"2b",	--587
		x"0c",	--588
		x"0c",	--589
		x"0c",	--590
		x"0c",	--591
		x"8d",	--592
		x"0c",	--593
		x"3c",	--594
		x"d0",	--595
		x"1a",	--596
		x"7d",	--597
		x"4d",	--598
		x"17",	--599
		x"7d",	--600
		x"78",	--601
		x"1a",	--602
		x"4b",	--603
		x"7b",	--604
		x"d0",	--605
		x"0a",	--606
		x"e9",	--607
		x"7b",	--608
		x"0a",	--609
		x"34",	--610
		x"0c",	--611
		x"0b",	--612
		x"0b",	--613
		x"0b",	--614
		x"0c",	--615
		x"8d",	--616
		x"0c",	--617
		x"3c",	--618
		x"d0",	--619
		x"7d",	--620
		x"4d",	--621
		x"e9",	--622
		x"9e",	--623
		x"00",	--624
		x"0f",	--625
		x"3a",	--626
		x"3b",	--627
		x"30",	--628
		x"1a",	--629
		x"de",	--630
		x"4b",	--631
		x"7b",	--632
		x"9f",	--633
		x"7b",	--634
		x"06",	--635
		x"0a",	--636
		x"0c",	--637
		x"0c",	--638
		x"0c",	--639
		x"0c",	--640
		x"8d",	--641
		x"0c",	--642
		x"3c",	--643
		x"a9",	--644
		x"1a",	--645
		x"ce",	--646
		x"4b",	--647
		x"7b",	--648
		x"bf",	--649
		x"7b",	--650
		x"06",	--651
		x"0a",	--652
		x"0c",	--653
		x"0c",	--654
		x"0c",	--655
		x"0c",	--656
		x"8d",	--657
		x"0c",	--658
		x"3c",	--659
		x"c9",	--660
		x"1a",	--661
		x"be",	--662
		x"8d",	--663
		x"0d",	--664
		x"30",	--665
		x"da",	--666
		x"b0",	--667
		x"3e",	--668
		x"21",	--669
		x"0c",	--670
		x"0f",	--671
		x"3a",	--672
		x"3b",	--673
		x"30",	--674
		x"0c",	--675
		x"ca",	--676
		x"0b",	--677
		x"0a",	--678
		x"0b",	--679
		x"0a",	--680
		x"8f",	--681
		x"00",	--682
		x"8f",	--683
		x"02",	--684
		x"8f",	--685
		x"04",	--686
		x"0c",	--687
		x"0d",	--688
		x"3e",	--689
		x"00",	--690
		x"3f",	--691
		x"6e",	--692
		x"b0",	--693
		x"d6",	--694
		x"8b",	--695
		x"02",	--696
		x"02",	--697
		x"32",	--698
		x"03",	--699
		x"82",	--700
		x"32",	--701
		x"b2",	--702
		x"18",	--703
		x"38",	--704
		x"9b",	--705
		x"3a",	--706
		x"06",	--707
		x"32",	--708
		x"0f",	--709
		x"3a",	--710
		x"3b",	--711
		x"30",	--712
		x"0b",	--713
		x"09",	--714
		x"08",	--715
		x"8f",	--716
		x"06",	--717
		x"bf",	--718
		x"00",	--719
		x"08",	--720
		x"2b",	--721
		x"1e",	--722
		x"02",	--723
		x"0f",	--724
		x"b0",	--725
		x"a2",	--726
		x"0c",	--727
		x"3d",	--728
		x"00",	--729
		x"b0",	--730
		x"4e",	--731
		x"08",	--732
		x"09",	--733
		x"1e",	--734
		x"06",	--735
		x"0f",	--736
		x"b0",	--737
		x"a2",	--738
		x"0c",	--739
		x"0d",	--740
		x"0e",	--741
		x"0f",	--742
		x"b0",	--743
		x"fe",	--744
		x"b0",	--745
		x"de",	--746
		x"8b",	--747
		x"04",	--748
		x"9b",	--749
		x"00",	--750
		x"38",	--751
		x"39",	--752
		x"3b",	--753
		x"30",	--754
		x"0b",	--755
		x"0a",	--756
		x"09",	--757
		x"0a",	--758
		x"0b",	--759
		x"8f",	--760
		x"06",	--761
		x"8f",	--762
		x"08",	--763
		x"29",	--764
		x"1e",	--765
		x"02",	--766
		x"0f",	--767
		x"b0",	--768
		x"a2",	--769
		x"0c",	--770
		x"0d",	--771
		x"0e",	--772
		x"0f",	--773
		x"b0",	--774
		x"4e",	--775
		x"0a",	--776
		x"0b",	--777
		x"1e",	--778
		x"06",	--779
		x"0f",	--780
		x"b0",	--781
		x"a2",	--782
		x"0c",	--783
		x"0d",	--784
		x"0e",	--785
		x"0f",	--786
		x"b0",	--787
		x"fe",	--788
		x"b0",	--789
		x"de",	--790
		x"89",	--791
		x"04",	--792
		x"39",	--793
		x"3a",	--794
		x"3b",	--795
		x"30",	--796
		x"0b",	--797
		x"0a",	--798
		x"92",	--799
		x"0c",	--800
		x"14",	--801
		x"3b",	--802
		x"20",	--803
		x"0a",	--804
		x"2b",	--805
		x"5f",	--806
		x"fc",	--807
		x"8f",	--808
		x"0f",	--809
		x"30",	--810
		x"ef",	--811
		x"b0",	--812
		x"3e",	--813
		x"31",	--814
		x"06",	--815
		x"1a",	--816
		x"3b",	--817
		x"06",	--818
		x"1a",	--819
		x"0c",	--820
		x"ef",	--821
		x"0f",	--822
		x"3a",	--823
		x"3b",	--824
		x"30",	--825
		x"1e",	--826
		x"0c",	--827
		x"3e",	--828
		x"20",	--829
		x"12",	--830
		x"0f",	--831
		x"0f",	--832
		x"0f",	--833
		x"0f",	--834
		x"3f",	--835
		x"1c",	--836
		x"ff",	--837
		x"68",	--838
		x"00",	--839
		x"bf",	--840
		x"3a",	--841
		x"02",	--842
		x"bf",	--843
		x"02",	--844
		x"04",	--845
		x"1e",	--846
		x"82",	--847
		x"0c",	--848
		x"30",	--849
		x"0b",	--850
		x"1b",	--851
		x"0c",	--852
		x"3b",	--853
		x"20",	--854
		x"12",	--855
		x"0c",	--856
		x"0c",	--857
		x"0c",	--858
		x"0c",	--859
		x"3c",	--860
		x"1c",	--861
		x"cc",	--862
		x"00",	--863
		x"8c",	--864
		x"02",	--865
		x"8c",	--866
		x"04",	--867
		x"1b",	--868
		x"82",	--869
		x"0c",	--870
		x"0f",	--871
		x"3b",	--872
		x"30",	--873
		x"3f",	--874
		x"fc",	--875
		x"0b",	--876
		x"31",	--877
		x"f0",	--878
		x"1b",	--879
		x"0c",	--880
		x"1b",	--881
		x"0f",	--882
		x"5f",	--883
		x"1c",	--884
		x"16",	--885
		x"3d",	--886
		x"22",	--887
		x"0c",	--888
		x"05",	--889
		x"3d",	--890
		x"06",	--891
		x"cd",	--892
		x"fa",	--893
		x"0e",	--894
		x"1c",	--895
		x"0c",	--896
		x"f8",	--897
		x"30",	--898
		x"f7",	--899
		x"b0",	--900
		x"3e",	--901
		x"21",	--902
		x"3f",	--903
		x"31",	--904
		x"10",	--905
		x"3b",	--906
		x"30",	--907
		x"0c",	--908
		x"81",	--909
		x"00",	--910
		x"6d",	--911
		x"4d",	--912
		x"24",	--913
		x"1e",	--914
		x"1f",	--915
		x"06",	--916
		x"6d",	--917
		x"4d",	--918
		x"11",	--919
		x"1e",	--920
		x"3f",	--921
		x"0e",	--922
		x"7d",	--923
		x"20",	--924
		x"f7",	--925
		x"ce",	--926
		x"ff",	--927
		x"0d",	--928
		x"0d",	--929
		x"0d",	--930
		x"8d",	--931
		x"00",	--932
		x"1f",	--933
		x"6d",	--934
		x"4d",	--935
		x"ef",	--936
		x"0e",	--937
		x"0e",	--938
		x"0c",	--939
		x"0c",	--940
		x"3c",	--941
		x"1c",	--942
		x"0e",	--943
		x"9c",	--944
		x"02",	--945
		x"31",	--946
		x"10",	--947
		x"3b",	--948
		x"30",	--949
		x"1f",	--950
		x"f1",	--951
		x"b2",	--952
		x"d2",	--953
		x"60",	--954
		x"b2",	--955
		x"b8",	--956
		x"72",	--957
		x"0f",	--958
		x"30",	--959
		x"0b",	--960
		x"0b",	--961
		x"1f",	--962
		x"0e",	--963
		x"3f",	--964
		x"20",	--965
		x"16",	--966
		x"0c",	--967
		x"0c",	--968
		x"0d",	--969
		x"0d",	--970
		x"0d",	--971
		x"0d",	--972
		x"3d",	--973
		x"dc",	--974
		x"8d",	--975
		x"00",	--976
		x"8d",	--977
		x"02",	--978
		x"8d",	--979
		x"06",	--980
		x"8d",	--981
		x"08",	--982
		x"0e",	--983
		x"1e",	--984
		x"82",	--985
		x"0e",	--986
		x"3b",	--987
		x"30",	--988
		x"3f",	--989
		x"fc",	--990
		x"0f",	--991
		x"0d",	--992
		x"0d",	--993
		x"0d",	--994
		x"0d",	--995
		x"3d",	--996
		x"dc",	--997
		x"8d",	--998
		x"02",	--999
		x"8d",	--1000
		x"04",	--1001
		x"9d",	--1002
		x"00",	--1003
		x"0f",	--1004
		x"30",	--1005
		x"0f",	--1006
		x"0e",	--1007
		x"0e",	--1008
		x"0e",	--1009
		x"0e",	--1010
		x"8e",	--1011
		x"dc",	--1012
		x"0f",	--1013
		x"30",	--1014
		x"0f",	--1015
		x"0e",	--1016
		x"0d",	--1017
		x"0c",	--1018
		x"0b",	--1019
		x"0a",	--1020
		x"92",	--1021
		x"0e",	--1022
		x"20",	--1023
		x"3b",	--1024
		x"de",	--1025
		x"0a",	--1026
		x"09",	--1027
		x"1f",	--1028
		x"8b",	--1029
		x"00",	--1030
		x"1a",	--1031
		x"3b",	--1032
		x"0a",	--1033
		x"1a",	--1034
		x"0e",	--1035
		x"13",	--1036
		x"8b",	--1037
		x"fe",	--1038
		x"f7",	--1039
		x"2f",	--1040
		x"1f",	--1041
		x"02",	--1042
		x"f0",	--1043
		x"8b",	--1044
		x"00",	--1045
		x"1f",	--1046
		x"06",	--1047
		x"9b",	--1048
		x"04",	--1049
		x"1a",	--1050
		x"3b",	--1051
		x"0a",	--1052
		x"1a",	--1053
		x"0e",	--1054
		x"ed",	--1055
		x"b2",	--1056
		x"fe",	--1057
		x"60",	--1058
		x"3a",	--1059
		x"3b",	--1060
		x"3c",	--1061
		x"3d",	--1062
		x"3e",	--1063
		x"3f",	--1064
		x"00",	--1065
		x"8f",	--1066
		x"00",	--1067
		x"0f",	--1068
		x"30",	--1069
		x"2f",	--1070
		x"2f",	--1071
		x"30",	--1072
		x"5e",	--1073
		x"81",	--1074
		x"3e",	--1075
		x"fc",	--1076
		x"c2",	--1077
		x"84",	--1078
		x"0f",	--1079
		x"30",	--1080
		x"3f",	--1081
		x"0f",	--1082
		x"5f",	--1083
		x"b6",	--1084
		x"8f",	--1085
		x"b0",	--1086
		x"62",	--1087
		x"30",	--1088
		x"0b",	--1089
		x"0b",	--1090
		x"0e",	--1091
		x"0e",	--1092
		x"0e",	--1093
		x"0e",	--1094
		x"0e",	--1095
		x"0f",	--1096
		x"b0",	--1097
		x"72",	--1098
		x"0f",	--1099
		x"b0",	--1100
		x"72",	--1101
		x"3b",	--1102
		x"30",	--1103
		x"0b",	--1104
		x"0a",	--1105
		x"0a",	--1106
		x"3b",	--1107
		x"07",	--1108
		x"0e",	--1109
		x"4d",	--1110
		x"7d",	--1111
		x"0f",	--1112
		x"03",	--1113
		x"0e",	--1114
		x"7d",	--1115
		x"fd",	--1116
		x"1e",	--1117
		x"0a",	--1118
		x"3f",	--1119
		x"31",	--1120
		x"b0",	--1121
		x"62",	--1122
		x"3b",	--1123
		x"3b",	--1124
		x"ef",	--1125
		x"3a",	--1126
		x"3b",	--1127
		x"30",	--1128
		x"3f",	--1129
		x"30",	--1130
		x"f5",	--1131
		x"0b",	--1132
		x"0b",	--1133
		x"0e",	--1134
		x"8e",	--1135
		x"8e",	--1136
		x"0f",	--1137
		x"b0",	--1138
		x"82",	--1139
		x"0f",	--1140
		x"b0",	--1141
		x"82",	--1142
		x"3b",	--1143
		x"30",	--1144
		x"0b",	--1145
		x"0a",	--1146
		x"0a",	--1147
		x"0b",	--1148
		x"0d",	--1149
		x"8d",	--1150
		x"8d",	--1151
		x"0f",	--1152
		x"b0",	--1153
		x"82",	--1154
		x"0f",	--1155
		x"b0",	--1156
		x"82",	--1157
		x"0c",	--1158
		x"0d",	--1159
		x"8d",	--1160
		x"8c",	--1161
		x"4d",	--1162
		x"0d",	--1163
		x"0f",	--1164
		x"b0",	--1165
		x"82",	--1166
		x"0f",	--1167
		x"b0",	--1168
		x"82",	--1169
		x"3a",	--1170
		x"3b",	--1171
		x"30",	--1172
		x"0b",	--1173
		x"0a",	--1174
		x"09",	--1175
		x"0a",	--1176
		x"0e",	--1177
		x"19",	--1178
		x"09",	--1179
		x"39",	--1180
		x"0b",	--1181
		x"0d",	--1182
		x"0d",	--1183
		x"6f",	--1184
		x"8f",	--1185
		x"b0",	--1186
		x"82",	--1187
		x"0b",	--1188
		x"0e",	--1189
		x"1b",	--1190
		x"3b",	--1191
		x"07",	--1192
		x"05",	--1193
		x"3f",	--1194
		x"20",	--1195
		x"b0",	--1196
		x"62",	--1197
		x"ef",	--1198
		x"3f",	--1199
		x"3a",	--1200
		x"b0",	--1201
		x"62",	--1202
		x"ea",	--1203
		x"39",	--1204
		x"3a",	--1205
		x"3b",	--1206
		x"30",	--1207
		x"0b",	--1208
		x"0a",	--1209
		x"09",	--1210
		x"0a",	--1211
		x"0e",	--1212
		x"17",	--1213
		x"09",	--1214
		x"39",	--1215
		x"0b",	--1216
		x"6f",	--1217
		x"8f",	--1218
		x"b0",	--1219
		x"72",	--1220
		x"0b",	--1221
		x"0e",	--1222
		x"1b",	--1223
		x"3b",	--1224
		x"07",	--1225
		x"f6",	--1226
		x"3f",	--1227
		x"20",	--1228
		x"b0",	--1229
		x"62",	--1230
		x"6f",	--1231
		x"8f",	--1232
		x"b0",	--1233
		x"72",	--1234
		x"0b",	--1235
		x"f2",	--1236
		x"39",	--1237
		x"3a",	--1238
		x"3b",	--1239
		x"30",	--1240
		x"0b",	--1241
		x"0a",	--1242
		x"09",	--1243
		x"31",	--1244
		x"ec",	--1245
		x"0b",	--1246
		x"0f",	--1247
		x"34",	--1248
		x"3b",	--1249
		x"0a",	--1250
		x"38",	--1251
		x"09",	--1252
		x"0a",	--1253
		x"0a",	--1254
		x"3e",	--1255
		x"0a",	--1256
		x"0f",	--1257
		x"b0",	--1258
		x"ce",	--1259
		x"7f",	--1260
		x"30",	--1261
		x"ca",	--1262
		x"00",	--1263
		x"19",	--1264
		x"3e",	--1265
		x"0a",	--1266
		x"0f",	--1267
		x"b0",	--1268
		x"9c",	--1269
		x"0b",	--1270
		x"3f",	--1271
		x"0a",	--1272
		x"eb",	--1273
		x"0a",	--1274
		x"1a",	--1275
		x"09",	--1276
		x"3e",	--1277
		x"0a",	--1278
		x"0f",	--1279
		x"b0",	--1280
		x"ce",	--1281
		x"7f",	--1282
		x"30",	--1283
		x"c9",	--1284
		x"00",	--1285
		x"3a",	--1286
		x"0f",	--1287
		x"0f",	--1288
		x"6f",	--1289
		x"8f",	--1290
		x"b0",	--1291
		x"62",	--1292
		x"0a",	--1293
		x"f7",	--1294
		x"31",	--1295
		x"14",	--1296
		x"39",	--1297
		x"3a",	--1298
		x"3b",	--1299
		x"30",	--1300
		x"3f",	--1301
		x"2d",	--1302
		x"b0",	--1303
		x"62",	--1304
		x"3b",	--1305
		x"1b",	--1306
		x"c5",	--1307
		x"1a",	--1308
		x"09",	--1309
		x"dd",	--1310
		x"0b",	--1311
		x"0a",	--1312
		x"09",	--1313
		x"0b",	--1314
		x"3b",	--1315
		x"39",	--1316
		x"6f",	--1317
		x"4f",	--1318
		x"0b",	--1319
		x"1a",	--1320
		x"8f",	--1321
		x"b0",	--1322
		x"62",	--1323
		x"0a",	--1324
		x"09",	--1325
		x"19",	--1326
		x"5f",	--1327
		x"01",	--1328
		x"4f",	--1329
		x"10",	--1330
		x"7f",	--1331
		x"25",	--1332
		x"f3",	--1333
		x"0a",	--1334
		x"1a",	--1335
		x"5f",	--1336
		x"01",	--1337
		x"7f",	--1338
		x"db",	--1339
		x"7f",	--1340
		x"54",	--1341
		x"ee",	--1342
		x"4f",	--1343
		x"0f",	--1344
		x"10",	--1345
		x"0e",	--1346
		x"39",	--1347
		x"3a",	--1348
		x"3b",	--1349
		x"30",	--1350
		x"09",	--1351
		x"29",	--1352
		x"1e",	--1353
		x"02",	--1354
		x"2f",	--1355
		x"b0",	--1356
		x"2a",	--1357
		x"0b",	--1358
		x"dd",	--1359
		x"09",	--1360
		x"29",	--1361
		x"2f",	--1362
		x"b0",	--1363
		x"d8",	--1364
		x"0b",	--1365
		x"d6",	--1366
		x"0f",	--1367
		x"2b",	--1368
		x"29",	--1369
		x"6f",	--1370
		x"4f",	--1371
		x"d0",	--1372
		x"19",	--1373
		x"8f",	--1374
		x"b0",	--1375
		x"62",	--1376
		x"7f",	--1377
		x"4f",	--1378
		x"fa",	--1379
		x"c8",	--1380
		x"09",	--1381
		x"29",	--1382
		x"1e",	--1383
		x"02",	--1384
		x"2f",	--1385
		x"b0",	--1386
		x"70",	--1387
		x"0b",	--1388
		x"bf",	--1389
		x"09",	--1390
		x"29",	--1391
		x"2e",	--1392
		x"0f",	--1393
		x"8f",	--1394
		x"8f",	--1395
		x"8f",	--1396
		x"8f",	--1397
		x"b0",	--1398
		x"f2",	--1399
		x"0b",	--1400
		x"b3",	--1401
		x"09",	--1402
		x"29",	--1403
		x"2f",	--1404
		x"b0",	--1405
		x"b2",	--1406
		x"0b",	--1407
		x"ac",	--1408
		x"09",	--1409
		x"29",	--1410
		x"2f",	--1411
		x"b0",	--1412
		x"62",	--1413
		x"0b",	--1414
		x"a5",	--1415
		x"09",	--1416
		x"29",	--1417
		x"2f",	--1418
		x"b0",	--1419
		x"82",	--1420
		x"0b",	--1421
		x"9e",	--1422
		x"09",	--1423
		x"29",	--1424
		x"2f",	--1425
		x"b0",	--1426
		x"a0",	--1427
		x"0b",	--1428
		x"97",	--1429
		x"3f",	--1430
		x"25",	--1431
		x"b0",	--1432
		x"62",	--1433
		x"92",	--1434
		x"0f",	--1435
		x"0e",	--1436
		x"1f",	--1437
		x"10",	--1438
		x"df",	--1439
		x"85",	--1440
		x"1c",	--1441
		x"1f",	--1442
		x"10",	--1443
		x"3f",	--1444
		x"3f",	--1445
		x"13",	--1446
		x"92",	--1447
		x"10",	--1448
		x"1e",	--1449
		x"10",	--1450
		x"1f",	--1451
		x"12",	--1452
		x"0e",	--1453
		x"02",	--1454
		x"92",	--1455
		x"12",	--1456
		x"f2",	--1457
		x"10",	--1458
		x"81",	--1459
		x"3e",	--1460
		x"3f",	--1461
		x"b1",	--1462
		x"f0",	--1463
		x"00",	--1464
		x"00",	--1465
		x"82",	--1466
		x"10",	--1467
		x"ec",	--1468
		x"b2",	--1469
		x"c3",	--1470
		x"82",	--1471
		x"f2",	--1472
		x"11",	--1473
		x"80",	--1474
		x"30",	--1475
		x"1e",	--1476
		x"10",	--1477
		x"1f",	--1478
		x"12",	--1479
		x"0e",	--1480
		x"05",	--1481
		x"1f",	--1482
		x"10",	--1483
		x"1f",	--1484
		x"12",	--1485
		x"30",	--1486
		x"1d",	--1487
		x"10",	--1488
		x"1e",	--1489
		x"12",	--1490
		x"3f",	--1491
		x"40",	--1492
		x"0f",	--1493
		x"0f",	--1494
		x"30",	--1495
		x"1f",	--1496
		x"12",	--1497
		x"5f",	--1498
		x"1c",	--1499
		x"1d",	--1500
		x"12",	--1501
		x"1e",	--1502
		x"10",	--1503
		x"0d",	--1504
		x"0b",	--1505
		x"1e",	--1506
		x"12",	--1507
		x"3e",	--1508
		x"3f",	--1509
		x"03",	--1510
		x"82",	--1511
		x"12",	--1512
		x"30",	--1513
		x"92",	--1514
		x"12",	--1515
		x"30",	--1516
		x"4f",	--1517
		x"30",	--1518
		x"0b",	--1519
		x"0a",	--1520
		x"0a",	--1521
		x"0b",	--1522
		x"0c",	--1523
		x"3d",	--1524
		x"00",	--1525
		x"b0",	--1526
		x"c2",	--1527
		x"0f",	--1528
		x"07",	--1529
		x"0e",	--1530
		x"0f",	--1531
		x"b0",	--1532
		x"12",	--1533
		x"3a",	--1534
		x"3b",	--1535
		x"30",	--1536
		x"0c",	--1537
		x"3d",	--1538
		x"00",	--1539
		x"0e",	--1540
		x"0f",	--1541
		x"b0",	--1542
		x"fe",	--1543
		x"b0",	--1544
		x"12",	--1545
		x"0e",	--1546
		x"3f",	--1547
		x"00",	--1548
		x"3a",	--1549
		x"3b",	--1550
		x"30",	--1551
		x"0b",	--1552
		x"0a",	--1553
		x"09",	--1554
		x"08",	--1555
		x"07",	--1556
		x"06",	--1557
		x"05",	--1558
		x"04",	--1559
		x"31",	--1560
		x"fa",	--1561
		x"08",	--1562
		x"6b",	--1563
		x"6b",	--1564
		x"67",	--1565
		x"6c",	--1566
		x"6c",	--1567
		x"e9",	--1568
		x"6b",	--1569
		x"02",	--1570
		x"30",	--1571
		x"a0",	--1572
		x"6c",	--1573
		x"e3",	--1574
		x"6c",	--1575
		x"bb",	--1576
		x"6b",	--1577
		x"df",	--1578
		x"91",	--1579
		x"02",	--1580
		x"00",	--1581
		x"1b",	--1582
		x"02",	--1583
		x"14",	--1584
		x"04",	--1585
		x"15",	--1586
		x"06",	--1587
		x"16",	--1588
		x"04",	--1589
		x"17",	--1590
		x"06",	--1591
		x"2c",	--1592
		x"0c",	--1593
		x"09",	--1594
		x"0c",	--1595
		x"bf",	--1596
		x"39",	--1597
		x"20",	--1598
		x"50",	--1599
		x"1c",	--1600
		x"d7",	--1601
		x"81",	--1602
		x"02",	--1603
		x"81",	--1604
		x"04",	--1605
		x"4c",	--1606
		x"7c",	--1607
		x"1f",	--1608
		x"0b",	--1609
		x"0a",	--1610
		x"0b",	--1611
		x"12",	--1612
		x"0b",	--1613
		x"0a",	--1614
		x"7c",	--1615
		x"fb",	--1616
		x"81",	--1617
		x"02",	--1618
		x"81",	--1619
		x"04",	--1620
		x"1c",	--1621
		x"0d",	--1622
		x"79",	--1623
		x"1f",	--1624
		x"04",	--1625
		x"0c",	--1626
		x"0d",	--1627
		x"79",	--1628
		x"fc",	--1629
		x"3c",	--1630
		x"3d",	--1631
		x"0c",	--1632
		x"0d",	--1633
		x"1a",	--1634
		x"0b",	--1635
		x"0c",	--1636
		x"02",	--1637
		x"0d",	--1638
		x"e5",	--1639
		x"16",	--1640
		x"02",	--1641
		x"17",	--1642
		x"04",	--1643
		x"06",	--1644
		x"07",	--1645
		x"5f",	--1646
		x"01",	--1647
		x"5f",	--1648
		x"01",	--1649
		x"28",	--1650
		x"c8",	--1651
		x"01",	--1652
		x"a8",	--1653
		x"02",	--1654
		x"0e",	--1655
		x"0f",	--1656
		x"0e",	--1657
		x"0f",	--1658
		x"88",	--1659
		x"04",	--1660
		x"88",	--1661
		x"06",	--1662
		x"f8",	--1663
		x"03",	--1664
		x"00",	--1665
		x"0f",	--1666
		x"4d",	--1667
		x"0f",	--1668
		x"31",	--1669
		x"06",	--1670
		x"34",	--1671
		x"35",	--1672
		x"36",	--1673
		x"37",	--1674
		x"38",	--1675
		x"39",	--1676
		x"3a",	--1677
		x"3b",	--1678
		x"30",	--1679
		x"2b",	--1680
		x"67",	--1681
		x"81",	--1682
		x"00",	--1683
		x"04",	--1684
		x"05",	--1685
		x"5f",	--1686
		x"01",	--1687
		x"5f",	--1688
		x"01",	--1689
		x"d8",	--1690
		x"4f",	--1691
		x"68",	--1692
		x"0e",	--1693
		x"0f",	--1694
		x"0e",	--1695
		x"0f",	--1696
		x"0f",	--1697
		x"69",	--1698
		x"c8",	--1699
		x"01",	--1700
		x"a8",	--1701
		x"02",	--1702
		x"88",	--1703
		x"04",	--1704
		x"88",	--1705
		x"06",	--1706
		x"0c",	--1707
		x"0d",	--1708
		x"3c",	--1709
		x"3d",	--1710
		x"3d",	--1711
		x"ff",	--1712
		x"05",	--1713
		x"3d",	--1714
		x"00",	--1715
		x"17",	--1716
		x"3c",	--1717
		x"15",	--1718
		x"1b",	--1719
		x"02",	--1720
		x"3b",	--1721
		x"0e",	--1722
		x"0f",	--1723
		x"0a",	--1724
		x"3b",	--1725
		x"0c",	--1726
		x"0d",	--1727
		x"3c",	--1728
		x"3d",	--1729
		x"3d",	--1730
		x"ff",	--1731
		x"f5",	--1732
		x"3c",	--1733
		x"88",	--1734
		x"04",	--1735
		x"88",	--1736
		x"06",	--1737
		x"88",	--1738
		x"02",	--1739
		x"f8",	--1740
		x"03",	--1741
		x"00",	--1742
		x"0f",	--1743
		x"b3",	--1744
		x"0c",	--1745
		x"0d",	--1746
		x"1c",	--1747
		x"0d",	--1748
		x"12",	--1749
		x"0f",	--1750
		x"0e",	--1751
		x"0a",	--1752
		x"0b",	--1753
		x"0a",	--1754
		x"0b",	--1755
		x"88",	--1756
		x"04",	--1757
		x"88",	--1758
		x"06",	--1759
		x"98",	--1760
		x"02",	--1761
		x"0f",	--1762
		x"a1",	--1763
		x"6b",	--1764
		x"9f",	--1765
		x"ad",	--1766
		x"00",	--1767
		x"9d",	--1768
		x"02",	--1769
		x"02",	--1770
		x"9d",	--1771
		x"04",	--1772
		x"04",	--1773
		x"9d",	--1774
		x"06",	--1775
		x"06",	--1776
		x"5e",	--1777
		x"01",	--1778
		x"5e",	--1779
		x"01",	--1780
		x"cd",	--1781
		x"01",	--1782
		x"0f",	--1783
		x"8c",	--1784
		x"06",	--1785
		x"07",	--1786
		x"9a",	--1787
		x"39",	--1788
		x"19",	--1789
		x"39",	--1790
		x"20",	--1791
		x"8f",	--1792
		x"3e",	--1793
		x"3c",	--1794
		x"b6",	--1795
		x"c1",	--1796
		x"0e",	--1797
		x"0f",	--1798
		x"0e",	--1799
		x"0f",	--1800
		x"97",	--1801
		x"0f",	--1802
		x"79",	--1803
		x"d8",	--1804
		x"01",	--1805
		x"a8",	--1806
		x"02",	--1807
		x"3e",	--1808
		x"3f",	--1809
		x"1e",	--1810
		x"0f",	--1811
		x"88",	--1812
		x"04",	--1813
		x"88",	--1814
		x"06",	--1815
		x"92",	--1816
		x"0c",	--1817
		x"7b",	--1818
		x"81",	--1819
		x"00",	--1820
		x"81",	--1821
		x"02",	--1822
		x"81",	--1823
		x"04",	--1824
		x"4d",	--1825
		x"7d",	--1826
		x"1f",	--1827
		x"0c",	--1828
		x"4b",	--1829
		x"0c",	--1830
		x"0d",	--1831
		x"12",	--1832
		x"0d",	--1833
		x"0c",	--1834
		x"7b",	--1835
		x"fb",	--1836
		x"81",	--1837
		x"02",	--1838
		x"81",	--1839
		x"04",	--1840
		x"1c",	--1841
		x"0d",	--1842
		x"79",	--1843
		x"1f",	--1844
		x"04",	--1845
		x"0c",	--1846
		x"0d",	--1847
		x"79",	--1848
		x"fc",	--1849
		x"3c",	--1850
		x"3d",	--1851
		x"0c",	--1852
		x"0d",	--1853
		x"1a",	--1854
		x"0b",	--1855
		x"0c",	--1856
		x"04",	--1857
		x"0d",	--1858
		x"02",	--1859
		x"0a",	--1860
		x"0b",	--1861
		x"14",	--1862
		x"02",	--1863
		x"15",	--1864
		x"04",	--1865
		x"04",	--1866
		x"05",	--1867
		x"49",	--1868
		x"0a",	--1869
		x"0b",	--1870
		x"18",	--1871
		x"6c",	--1872
		x"33",	--1873
		x"df",	--1874
		x"01",	--1875
		x"01",	--1876
		x"2f",	--1877
		x"3f",	--1878
		x"c8",	--1879
		x"2c",	--1880
		x"31",	--1881
		x"e0",	--1882
		x"81",	--1883
		x"04",	--1884
		x"81",	--1885
		x"06",	--1886
		x"81",	--1887
		x"00",	--1888
		x"81",	--1889
		x"02",	--1890
		x"0e",	--1891
		x"3e",	--1892
		x"18",	--1893
		x"0f",	--1894
		x"2f",	--1895
		x"b0",	--1896
		x"d4",	--1897
		x"0e",	--1898
		x"3e",	--1899
		x"10",	--1900
		x"0f",	--1901
		x"b0",	--1902
		x"d4",	--1903
		x"0d",	--1904
		x"3d",	--1905
		x"0e",	--1906
		x"3e",	--1907
		x"10",	--1908
		x"0f",	--1909
		x"3f",	--1910
		x"18",	--1911
		x"b0",	--1912
		x"20",	--1913
		x"b0",	--1914
		x"f6",	--1915
		x"31",	--1916
		x"20",	--1917
		x"30",	--1918
		x"31",	--1919
		x"e0",	--1920
		x"81",	--1921
		x"04",	--1922
		x"81",	--1923
		x"06",	--1924
		x"81",	--1925
		x"00",	--1926
		x"81",	--1927
		x"02",	--1928
		x"0e",	--1929
		x"3e",	--1930
		x"18",	--1931
		x"0f",	--1932
		x"2f",	--1933
		x"b0",	--1934
		x"d4",	--1935
		x"0e",	--1936
		x"3e",	--1937
		x"10",	--1938
		x"0f",	--1939
		x"b0",	--1940
		x"d4",	--1941
		x"d1",	--1942
		x"11",	--1943
		x"0d",	--1944
		x"3d",	--1945
		x"0e",	--1946
		x"3e",	--1947
		x"10",	--1948
		x"0f",	--1949
		x"3f",	--1950
		x"18",	--1951
		x"b0",	--1952
		x"20",	--1953
		x"b0",	--1954
		x"f6",	--1955
		x"31",	--1956
		x"20",	--1957
		x"30",	--1958
		x"0b",	--1959
		x"0a",	--1960
		x"09",	--1961
		x"08",	--1962
		x"07",	--1963
		x"06",	--1964
		x"05",	--1965
		x"04",	--1966
		x"31",	--1967
		x"dc",	--1968
		x"81",	--1969
		x"04",	--1970
		x"81",	--1971
		x"06",	--1972
		x"81",	--1973
		x"00",	--1974
		x"81",	--1975
		x"02",	--1976
		x"0e",	--1977
		x"3e",	--1978
		x"18",	--1979
		x"0f",	--1980
		x"2f",	--1981
		x"b0",	--1982
		x"d4",	--1983
		x"0e",	--1984
		x"3e",	--1985
		x"10",	--1986
		x"0f",	--1987
		x"b0",	--1988
		x"d4",	--1989
		x"5f",	--1990
		x"18",	--1991
		x"6f",	--1992
		x"b6",	--1993
		x"5e",	--1994
		x"10",	--1995
		x"6e",	--1996
		x"d9",	--1997
		x"6f",	--1998
		x"ae",	--1999
		x"6e",	--2000
		x"e2",	--2001
		x"6f",	--2002
		x"ac",	--2003
		x"6e",	--2004
		x"d1",	--2005
		x"14",	--2006
		x"1c",	--2007
		x"15",	--2008
		x"1e",	--2009
		x"18",	--2010
		x"14",	--2011
		x"19",	--2012
		x"16",	--2013
		x"3c",	--2014
		x"20",	--2015
		x"0e",	--2016
		x"0f",	--2017
		x"06",	--2018
		x"07",	--2019
		x"81",	--2020
		x"20",	--2021
		x"81",	--2022
		x"22",	--2023
		x"0a",	--2024
		x"0b",	--2025
		x"81",	--2026
		x"20",	--2027
		x"08",	--2028
		x"08",	--2029
		x"09",	--2030
		x"12",	--2031
		x"05",	--2032
		x"04",	--2033
		x"b1",	--2034
		x"20",	--2035
		x"19",	--2036
		x"14",	--2037
		x"0d",	--2038
		x"0a",	--2039
		x"0b",	--2040
		x"0e",	--2041
		x"0f",	--2042
		x"1c",	--2043
		x"0d",	--2044
		x"0b",	--2045
		x"03",	--2046
		x"0b",	--2047
		x"0c",	--2048
		x"0d",	--2049
		x"0e",	--2050
		x"0f",	--2051
		x"06",	--2052
		x"07",	--2053
		x"09",	--2054
		x"e5",	--2055
		x"16",	--2056
		x"07",	--2057
		x"e2",	--2058
		x"0a",	--2059
		x"f5",	--2060
		x"f2",	--2061
		x"81",	--2062
		x"20",	--2063
		x"81",	--2064
		x"22",	--2065
		x"0c",	--2066
		x"1a",	--2067
		x"1a",	--2068
		x"1a",	--2069
		x"12",	--2070
		x"06",	--2071
		x"26",	--2072
		x"81",	--2073
		x"0a",	--2074
		x"5d",	--2075
		x"d1",	--2076
		x"11",	--2077
		x"19",	--2078
		x"83",	--2079
		x"c1",	--2080
		x"09",	--2081
		x"0c",	--2082
		x"3c",	--2083
		x"3f",	--2084
		x"00",	--2085
		x"18",	--2086
		x"1d",	--2087
		x"0a",	--2088
		x"3d",	--2089
		x"1a",	--2090
		x"20",	--2091
		x"1b",	--2092
		x"22",	--2093
		x"0c",	--2094
		x"0e",	--2095
		x"0f",	--2096
		x"0b",	--2097
		x"2a",	--2098
		x"0a",	--2099
		x"0b",	--2100
		x"3d",	--2101
		x"3f",	--2102
		x"00",	--2103
		x"f5",	--2104
		x"81",	--2105
		x"20",	--2106
		x"81",	--2107
		x"22",	--2108
		x"81",	--2109
		x"0a",	--2110
		x"0c",	--2111
		x"0d",	--2112
		x"3c",	--2113
		x"7f",	--2114
		x"0d",	--2115
		x"3c",	--2116
		x"40",	--2117
		x"44",	--2118
		x"81",	--2119
		x"0c",	--2120
		x"81",	--2121
		x"0e",	--2122
		x"f1",	--2123
		x"03",	--2124
		x"08",	--2125
		x"0f",	--2126
		x"3f",	--2127
		x"b0",	--2128
		x"f6",	--2129
		x"31",	--2130
		x"24",	--2131
		x"34",	--2132
		x"35",	--2133
		x"36",	--2134
		x"37",	--2135
		x"38",	--2136
		x"39",	--2137
		x"3a",	--2138
		x"3b",	--2139
		x"30",	--2140
		x"1e",	--2141
		x"0f",	--2142
		x"d3",	--2143
		x"3a",	--2144
		x"03",	--2145
		x"08",	--2146
		x"1e",	--2147
		x"10",	--2148
		x"1c",	--2149
		x"20",	--2150
		x"1d",	--2151
		x"22",	--2152
		x"12",	--2153
		x"0d",	--2154
		x"0c",	--2155
		x"06",	--2156
		x"07",	--2157
		x"06",	--2158
		x"37",	--2159
		x"00",	--2160
		x"81",	--2161
		x"20",	--2162
		x"81",	--2163
		x"22",	--2164
		x"12",	--2165
		x"0f",	--2166
		x"0e",	--2167
		x"1a",	--2168
		x"0f",	--2169
		x"e7",	--2170
		x"81",	--2171
		x"0a",	--2172
		x"a6",	--2173
		x"6e",	--2174
		x"36",	--2175
		x"5f",	--2176
		x"d1",	--2177
		x"11",	--2178
		x"19",	--2179
		x"20",	--2180
		x"c1",	--2181
		x"19",	--2182
		x"0f",	--2183
		x"3f",	--2184
		x"18",	--2185
		x"c5",	--2186
		x"0d",	--2187
		x"ba",	--2188
		x"0c",	--2189
		x"0d",	--2190
		x"3c",	--2191
		x"80",	--2192
		x"0d",	--2193
		x"0c",	--2194
		x"b3",	--2195
		x"0d",	--2196
		x"b1",	--2197
		x"81",	--2198
		x"20",	--2199
		x"03",	--2200
		x"81",	--2201
		x"22",	--2202
		x"ab",	--2203
		x"3e",	--2204
		x"40",	--2205
		x"0f",	--2206
		x"3e",	--2207
		x"80",	--2208
		x"3f",	--2209
		x"a4",	--2210
		x"4d",	--2211
		x"7b",	--2212
		x"4f",	--2213
		x"de",	--2214
		x"5f",	--2215
		x"d1",	--2216
		x"11",	--2217
		x"19",	--2218
		x"06",	--2219
		x"c1",	--2220
		x"11",	--2221
		x"0f",	--2222
		x"3f",	--2223
		x"10",	--2224
		x"9e",	--2225
		x"4f",	--2226
		x"f8",	--2227
		x"6f",	--2228
		x"f1",	--2229
		x"3f",	--2230
		x"c8",	--2231
		x"97",	--2232
		x"0b",	--2233
		x"0a",	--2234
		x"09",	--2235
		x"08",	--2236
		x"07",	--2237
		x"31",	--2238
		x"e8",	--2239
		x"81",	--2240
		x"04",	--2241
		x"81",	--2242
		x"06",	--2243
		x"81",	--2244
		x"00",	--2245
		x"81",	--2246
		x"02",	--2247
		x"0e",	--2248
		x"3e",	--2249
		x"10",	--2250
		x"0f",	--2251
		x"2f",	--2252
		x"b0",	--2253
		x"d4",	--2254
		x"0e",	--2255
		x"3e",	--2256
		x"0f",	--2257
		x"b0",	--2258
		x"d4",	--2259
		x"5f",	--2260
		x"10",	--2261
		x"6f",	--2262
		x"5d",	--2263
		x"5e",	--2264
		x"08",	--2265
		x"6e",	--2266
		x"82",	--2267
		x"d1",	--2268
		x"09",	--2269
		x"11",	--2270
		x"6f",	--2271
		x"58",	--2272
		x"6f",	--2273
		x"56",	--2274
		x"6e",	--2275
		x"6f",	--2276
		x"6e",	--2277
		x"4c",	--2278
		x"1d",	--2279
		x"12",	--2280
		x"1d",	--2281
		x"0a",	--2282
		x"81",	--2283
		x"12",	--2284
		x"1e",	--2285
		x"14",	--2286
		x"1f",	--2287
		x"16",	--2288
		x"18",	--2289
		x"0c",	--2290
		x"19",	--2291
		x"0e",	--2292
		x"0f",	--2293
		x"1e",	--2294
		x"0e",	--2295
		x"0f",	--2296
		x"3d",	--2297
		x"81",	--2298
		x"12",	--2299
		x"37",	--2300
		x"1f",	--2301
		x"0c",	--2302
		x"3d",	--2303
		x"00",	--2304
		x"0a",	--2305
		x"0b",	--2306
		x"0b",	--2307
		x"0a",	--2308
		x"0b",	--2309
		x"0e",	--2310
		x"0f",	--2311
		x"12",	--2312
		x"0d",	--2313
		x"0c",	--2314
		x"0e",	--2315
		x"0f",	--2316
		x"37",	--2317
		x"0b",	--2318
		x"0f",	--2319
		x"f7",	--2320
		x"f2",	--2321
		x"0e",	--2322
		x"f4",	--2323
		x"ef",	--2324
		x"09",	--2325
		x"e5",	--2326
		x"0e",	--2327
		x"e3",	--2328
		x"dd",	--2329
		x"0c",	--2330
		x"0d",	--2331
		x"3c",	--2332
		x"7f",	--2333
		x"0d",	--2334
		x"3c",	--2335
		x"40",	--2336
		x"1c",	--2337
		x"81",	--2338
		x"14",	--2339
		x"81",	--2340
		x"16",	--2341
		x"0f",	--2342
		x"3f",	--2343
		x"10",	--2344
		x"b0",	--2345
		x"f6",	--2346
		x"31",	--2347
		x"18",	--2348
		x"37",	--2349
		x"38",	--2350
		x"39",	--2351
		x"3a",	--2352
		x"3b",	--2353
		x"30",	--2354
		x"e1",	--2355
		x"10",	--2356
		x"0f",	--2357
		x"3f",	--2358
		x"10",	--2359
		x"f0",	--2360
		x"4f",	--2361
		x"fa",	--2362
		x"3f",	--2363
		x"c8",	--2364
		x"eb",	--2365
		x"0d",	--2366
		x"e2",	--2367
		x"0c",	--2368
		x"0d",	--2369
		x"3c",	--2370
		x"80",	--2371
		x"0d",	--2372
		x"0c",	--2373
		x"db",	--2374
		x"0d",	--2375
		x"d9",	--2376
		x"0e",	--2377
		x"02",	--2378
		x"0f",	--2379
		x"d5",	--2380
		x"3a",	--2381
		x"40",	--2382
		x"0b",	--2383
		x"3a",	--2384
		x"80",	--2385
		x"3b",	--2386
		x"ce",	--2387
		x"81",	--2388
		x"14",	--2389
		x"81",	--2390
		x"16",	--2391
		x"81",	--2392
		x"12",	--2393
		x"0f",	--2394
		x"3f",	--2395
		x"10",	--2396
		x"cb",	--2397
		x"0f",	--2398
		x"3f",	--2399
		x"c8",	--2400
		x"31",	--2401
		x"e8",	--2402
		x"81",	--2403
		x"04",	--2404
		x"81",	--2405
		x"06",	--2406
		x"81",	--2407
		x"00",	--2408
		x"81",	--2409
		x"02",	--2410
		x"0e",	--2411
		x"3e",	--2412
		x"10",	--2413
		x"0f",	--2414
		x"2f",	--2415
		x"b0",	--2416
		x"d4",	--2417
		x"0e",	--2418
		x"3e",	--2419
		x"0f",	--2420
		x"b0",	--2421
		x"d4",	--2422
		x"e1",	--2423
		x"10",	--2424
		x"0d",	--2425
		x"e1",	--2426
		x"08",	--2427
		x"0a",	--2428
		x"0e",	--2429
		x"3e",	--2430
		x"0f",	--2431
		x"3f",	--2432
		x"10",	--2433
		x"b0",	--2434
		x"f8",	--2435
		x"31",	--2436
		x"18",	--2437
		x"30",	--2438
		x"3f",	--2439
		x"fb",	--2440
		x"31",	--2441
		x"f4",	--2442
		x"81",	--2443
		x"00",	--2444
		x"81",	--2445
		x"02",	--2446
		x"0e",	--2447
		x"2e",	--2448
		x"0f",	--2449
		x"b0",	--2450
		x"d4",	--2451
		x"5f",	--2452
		x"04",	--2453
		x"6f",	--2454
		x"28",	--2455
		x"27",	--2456
		x"6f",	--2457
		x"07",	--2458
		x"1d",	--2459
		x"06",	--2460
		x"0d",	--2461
		x"21",	--2462
		x"3d",	--2463
		x"1f",	--2464
		x"09",	--2465
		x"c1",	--2466
		x"05",	--2467
		x"26",	--2468
		x"3e",	--2469
		x"3f",	--2470
		x"ff",	--2471
		x"31",	--2472
		x"0c",	--2473
		x"30",	--2474
		x"1e",	--2475
		x"08",	--2476
		x"1f",	--2477
		x"0a",	--2478
		x"3c",	--2479
		x"1e",	--2480
		x"4c",	--2481
		x"4d",	--2482
		x"7d",	--2483
		x"1f",	--2484
		x"0f",	--2485
		x"c1",	--2486
		x"05",	--2487
		x"ef",	--2488
		x"3e",	--2489
		x"3f",	--2490
		x"1e",	--2491
		x"0f",	--2492
		x"31",	--2493
		x"0c",	--2494
		x"30",	--2495
		x"0e",	--2496
		x"0f",	--2497
		x"31",	--2498
		x"0c",	--2499
		x"30",	--2500
		x"12",	--2501
		x"0f",	--2502
		x"0e",	--2503
		x"7d",	--2504
		x"fb",	--2505
		x"eb",	--2506
		x"0e",	--2507
		x"3f",	--2508
		x"00",	--2509
		x"31",	--2510
		x"0c",	--2511
		x"30",	--2512
		x"0b",	--2513
		x"0a",	--2514
		x"09",	--2515
		x"08",	--2516
		x"31",	--2517
		x"0a",	--2518
		x"0b",	--2519
		x"c1",	--2520
		x"01",	--2521
		x"0e",	--2522
		x"0d",	--2523
		x"0b",	--2524
		x"0b",	--2525
		x"e1",	--2526
		x"00",	--2527
		x"0f",	--2528
		x"b0",	--2529
		x"f6",	--2530
		x"31",	--2531
		x"38",	--2532
		x"39",	--2533
		x"3a",	--2534
		x"3b",	--2535
		x"30",	--2536
		x"f1",	--2537
		x"03",	--2538
		x"00",	--2539
		x"b1",	--2540
		x"1e",	--2541
		x"02",	--2542
		x"81",	--2543
		x"04",	--2544
		x"81",	--2545
		x"06",	--2546
		x"0e",	--2547
		x"0f",	--2548
		x"b0",	--2549
		x"84",	--2550
		x"3f",	--2551
		x"0f",	--2552
		x"18",	--2553
		x"e5",	--2554
		x"81",	--2555
		x"04",	--2556
		x"81",	--2557
		x"06",	--2558
		x"4e",	--2559
		x"7e",	--2560
		x"1f",	--2561
		x"06",	--2562
		x"3e",	--2563
		x"1e",	--2564
		x"0e",	--2565
		x"81",	--2566
		x"02",	--2567
		x"d7",	--2568
		x"91",	--2569
		x"04",	--2570
		x"04",	--2571
		x"91",	--2572
		x"06",	--2573
		x"06",	--2574
		x"7e",	--2575
		x"f8",	--2576
		x"f1",	--2577
		x"0e",	--2578
		x"3e",	--2579
		x"1e",	--2580
		x"1c",	--2581
		x"0d",	--2582
		x"48",	--2583
		x"78",	--2584
		x"1f",	--2585
		x"04",	--2586
		x"0c",	--2587
		x"0d",	--2588
		x"78",	--2589
		x"fc",	--2590
		x"3c",	--2591
		x"3d",	--2592
		x"0c",	--2593
		x"0d",	--2594
		x"18",	--2595
		x"09",	--2596
		x"0c",	--2597
		x"04",	--2598
		x"0d",	--2599
		x"02",	--2600
		x"08",	--2601
		x"09",	--2602
		x"7e",	--2603
		x"1f",	--2604
		x"0e",	--2605
		x"0d",	--2606
		x"0e",	--2607
		x"0d",	--2608
		x"0e",	--2609
		x"81",	--2610
		x"04",	--2611
		x"81",	--2612
		x"06",	--2613
		x"3e",	--2614
		x"1e",	--2615
		x"0e",	--2616
		x"81",	--2617
		x"02",	--2618
		x"a4",	--2619
		x"12",	--2620
		x"0b",	--2621
		x"0a",	--2622
		x"7e",	--2623
		x"fb",	--2624
		x"ec",	--2625
		x"0b",	--2626
		x"0a",	--2627
		x"09",	--2628
		x"1f",	--2629
		x"17",	--2630
		x"3e",	--2631
		x"00",	--2632
		x"2c",	--2633
		x"3a",	--2634
		x"18",	--2635
		x"0b",	--2636
		x"39",	--2637
		x"0c",	--2638
		x"0d",	--2639
		x"4f",	--2640
		x"4f",	--2641
		x"17",	--2642
		x"3c",	--2643
		x"d0",	--2644
		x"6e",	--2645
		x"0f",	--2646
		x"0a",	--2647
		x"0b",	--2648
		x"0f",	--2649
		x"39",	--2650
		x"3a",	--2651
		x"3b",	--2652
		x"30",	--2653
		x"3f",	--2654
		x"00",	--2655
		x"0f",	--2656
		x"3a",	--2657
		x"0b",	--2658
		x"39",	--2659
		x"18",	--2660
		x"0c",	--2661
		x"0d",	--2662
		x"4f",	--2663
		x"4f",	--2664
		x"e9",	--2665
		x"12",	--2666
		x"0d",	--2667
		x"0c",	--2668
		x"7f",	--2669
		x"fb",	--2670
		x"e3",	--2671
		x"3a",	--2672
		x"10",	--2673
		x"0b",	--2674
		x"39",	--2675
		x"10",	--2676
		x"ef",	--2677
		x"3a",	--2678
		x"20",	--2679
		x"0b",	--2680
		x"09",	--2681
		x"ea",	--2682
		x"0b",	--2683
		x"0a",	--2684
		x"09",	--2685
		x"08",	--2686
		x"07",	--2687
		x"0d",	--2688
		x"1e",	--2689
		x"04",	--2690
		x"1f",	--2691
		x"06",	--2692
		x"5a",	--2693
		x"01",	--2694
		x"6c",	--2695
		x"6c",	--2696
		x"70",	--2697
		x"6c",	--2698
		x"6a",	--2699
		x"6c",	--2700
		x"36",	--2701
		x"0e",	--2702
		x"32",	--2703
		x"1b",	--2704
		x"02",	--2705
		x"3b",	--2706
		x"82",	--2707
		x"6d",	--2708
		x"3b",	--2709
		x"80",	--2710
		x"5e",	--2711
		x"0c",	--2712
		x"0d",	--2713
		x"3c",	--2714
		x"7f",	--2715
		x"0d",	--2716
		x"3c",	--2717
		x"40",	--2718
		x"40",	--2719
		x"3e",	--2720
		x"3f",	--2721
		x"0f",	--2722
		x"0f",	--2723
		x"4a",	--2724
		x"0d",	--2725
		x"3d",	--2726
		x"7f",	--2727
		x"12",	--2728
		x"0f",	--2729
		x"0e",	--2730
		x"12",	--2731
		x"0f",	--2732
		x"0e",	--2733
		x"12",	--2734
		x"0f",	--2735
		x"0e",	--2736
		x"12",	--2737
		x"0f",	--2738
		x"0e",	--2739
		x"12",	--2740
		x"0f",	--2741
		x"0e",	--2742
		x"12",	--2743
		x"0f",	--2744
		x"0e",	--2745
		x"12",	--2746
		x"0f",	--2747
		x"0e",	--2748
		x"3e",	--2749
		x"3f",	--2750
		x"7f",	--2751
		x"4d",	--2752
		x"05",	--2753
		x"0f",	--2754
		x"cc",	--2755
		x"4d",	--2756
		x"0e",	--2757
		x"0f",	--2758
		x"4d",	--2759
		x"0d",	--2760
		x"0d",	--2761
		x"0d",	--2762
		x"0d",	--2763
		x"0d",	--2764
		x"0d",	--2765
		x"0d",	--2766
		x"0c",	--2767
		x"3c",	--2768
		x"7f",	--2769
		x"0c",	--2770
		x"4f",	--2771
		x"0f",	--2772
		x"0f",	--2773
		x"0f",	--2774
		x"0d",	--2775
		x"0d",	--2776
		x"0f",	--2777
		x"37",	--2778
		x"38",	--2779
		x"39",	--2780
		x"3a",	--2781
		x"3b",	--2782
		x"30",	--2783
		x"0d",	--2784
		x"be",	--2785
		x"0c",	--2786
		x"0d",	--2787
		x"3c",	--2788
		x"80",	--2789
		x"0d",	--2790
		x"0c",	--2791
		x"02",	--2792
		x"0d",	--2793
		x"b8",	--2794
		x"3e",	--2795
		x"40",	--2796
		x"0f",	--2797
		x"b4",	--2798
		x"12",	--2799
		x"0f",	--2800
		x"0e",	--2801
		x"0d",	--2802
		x"3d",	--2803
		x"80",	--2804
		x"b2",	--2805
		x"7d",	--2806
		x"0e",	--2807
		x"0f",	--2808
		x"cd",	--2809
		x"0e",	--2810
		x"3f",	--2811
		x"10",	--2812
		x"3e",	--2813
		x"3f",	--2814
		x"7f",	--2815
		x"7d",	--2816
		x"c5",	--2817
		x"37",	--2818
		x"82",	--2819
		x"07",	--2820
		x"37",	--2821
		x"1a",	--2822
		x"4f",	--2823
		x"0c",	--2824
		x"0d",	--2825
		x"4b",	--2826
		x"7b",	--2827
		x"1f",	--2828
		x"05",	--2829
		x"12",	--2830
		x"0d",	--2831
		x"0c",	--2832
		x"7b",	--2833
		x"fb",	--2834
		x"18",	--2835
		x"09",	--2836
		x"77",	--2837
		x"1f",	--2838
		x"04",	--2839
		x"08",	--2840
		x"09",	--2841
		x"77",	--2842
		x"fc",	--2843
		x"38",	--2844
		x"39",	--2845
		x"08",	--2846
		x"09",	--2847
		x"1e",	--2848
		x"0f",	--2849
		x"08",	--2850
		x"04",	--2851
		x"09",	--2852
		x"02",	--2853
		x"0e",	--2854
		x"0f",	--2855
		x"08",	--2856
		x"09",	--2857
		x"08",	--2858
		x"09",	--2859
		x"0e",	--2860
		x"0f",	--2861
		x"3e",	--2862
		x"7f",	--2863
		x"0f",	--2864
		x"3e",	--2865
		x"40",	--2866
		x"26",	--2867
		x"38",	--2868
		x"3f",	--2869
		x"09",	--2870
		x"0e",	--2871
		x"0f",	--2872
		x"12",	--2873
		x"0f",	--2874
		x"0e",	--2875
		x"12",	--2876
		x"0f",	--2877
		x"0e",	--2878
		x"12",	--2879
		x"0f",	--2880
		x"0e",	--2881
		x"12",	--2882
		x"0f",	--2883
		x"0e",	--2884
		x"12",	--2885
		x"0f",	--2886
		x"0e",	--2887
		x"12",	--2888
		x"0f",	--2889
		x"0e",	--2890
		x"12",	--2891
		x"0f",	--2892
		x"0e",	--2893
		x"3e",	--2894
		x"3f",	--2895
		x"7f",	--2896
		x"5d",	--2897
		x"39",	--2898
		x"00",	--2899
		x"72",	--2900
		x"4d",	--2901
		x"70",	--2902
		x"08",	--2903
		x"09",	--2904
		x"da",	--2905
		x"0f",	--2906
		x"d8",	--2907
		x"0e",	--2908
		x"0f",	--2909
		x"3e",	--2910
		x"80",	--2911
		x"0f",	--2912
		x"0e",	--2913
		x"04",	--2914
		x"38",	--2915
		x"40",	--2916
		x"09",	--2917
		x"d0",	--2918
		x"0f",	--2919
		x"ce",	--2920
		x"f9",	--2921
		x"0b",	--2922
		x"0a",	--2923
		x"2a",	--2924
		x"5b",	--2925
		x"02",	--2926
		x"3b",	--2927
		x"7f",	--2928
		x"1d",	--2929
		x"02",	--2930
		x"12",	--2931
		x"0d",	--2932
		x"12",	--2933
		x"0d",	--2934
		x"12",	--2935
		x"0d",	--2936
		x"12",	--2937
		x"0d",	--2938
		x"12",	--2939
		x"0d",	--2940
		x"12",	--2941
		x"0d",	--2942
		x"12",	--2943
		x"0d",	--2944
		x"4d",	--2945
		x"5f",	--2946
		x"03",	--2947
		x"3f",	--2948
		x"80",	--2949
		x"0f",	--2950
		x"0f",	--2951
		x"ce",	--2952
		x"01",	--2953
		x"0d",	--2954
		x"2d",	--2955
		x"0a",	--2956
		x"51",	--2957
		x"be",	--2958
		x"82",	--2959
		x"02",	--2960
		x"0c",	--2961
		x"0d",	--2962
		x"0c",	--2963
		x"0d",	--2964
		x"0c",	--2965
		x"0d",	--2966
		x"0c",	--2967
		x"0d",	--2968
		x"0c",	--2969
		x"0d",	--2970
		x"0c",	--2971
		x"0d",	--2972
		x"0c",	--2973
		x"0d",	--2974
		x"0c",	--2975
		x"0d",	--2976
		x"fe",	--2977
		x"03",	--2978
		x"00",	--2979
		x"3d",	--2980
		x"00",	--2981
		x"0b",	--2982
		x"3f",	--2983
		x"81",	--2984
		x"0c",	--2985
		x"0d",	--2986
		x"0a",	--2987
		x"3f",	--2988
		x"3d",	--2989
		x"00",	--2990
		x"f9",	--2991
		x"8e",	--2992
		x"02",	--2993
		x"8e",	--2994
		x"04",	--2995
		x"8e",	--2996
		x"06",	--2997
		x"3a",	--2998
		x"3b",	--2999
		x"30",	--3000
		x"3d",	--3001
		x"ff",	--3002
		x"2a",	--3003
		x"3d",	--3004
		x"81",	--3005
		x"8e",	--3006
		x"02",	--3007
		x"fe",	--3008
		x"03",	--3009
		x"00",	--3010
		x"0c",	--3011
		x"0d",	--3012
		x"0c",	--3013
		x"0d",	--3014
		x"0c",	--3015
		x"0d",	--3016
		x"0c",	--3017
		x"0d",	--3018
		x"0c",	--3019
		x"0d",	--3020
		x"0c",	--3021
		x"0d",	--3022
		x"0c",	--3023
		x"0d",	--3024
		x"0c",	--3025
		x"0d",	--3026
		x"0a",	--3027
		x"0b",	--3028
		x"0a",	--3029
		x"3b",	--3030
		x"00",	--3031
		x"8e",	--3032
		x"04",	--3033
		x"8e",	--3034
		x"06",	--3035
		x"3a",	--3036
		x"3b",	--3037
		x"30",	--3038
		x"0b",	--3039
		x"ad",	--3040
		x"ee",	--3041
		x"00",	--3042
		x"3a",	--3043
		x"3b",	--3044
		x"30",	--3045
		x"0a",	--3046
		x"0c",	--3047
		x"0c",	--3048
		x"0d",	--3049
		x"0c",	--3050
		x"3d",	--3051
		x"10",	--3052
		x"0c",	--3053
		x"02",	--3054
		x"0d",	--3055
		x"08",	--3056
		x"de",	--3057
		x"00",	--3058
		x"e4",	--3059
		x"0b",	--3060
		x"f2",	--3061
		x"ee",	--3062
		x"00",	--3063
		x"e3",	--3064
		x"ce",	--3065
		x"00",	--3066
		x"dc",	--3067
		x"0b",	--3068
		x"6d",	--3069
		x"6d",	--3070
		x"12",	--3071
		x"6c",	--3072
		x"6c",	--3073
		x"0f",	--3074
		x"6d",	--3075
		x"41",	--3076
		x"6c",	--3077
		x"11",	--3078
		x"6d",	--3079
		x"0d",	--3080
		x"6c",	--3081
		x"14",	--3082
		x"5d",	--3083
		x"01",	--3084
		x"5d",	--3085
		x"01",	--3086
		x"14",	--3087
		x"4d",	--3088
		x"09",	--3089
		x"1e",	--3090
		x"0f",	--3091
		x"3b",	--3092
		x"30",	--3093
		x"6c",	--3094
		x"28",	--3095
		x"ce",	--3096
		x"01",	--3097
		x"f7",	--3098
		x"3e",	--3099
		x"0f",	--3100
		x"3b",	--3101
		x"30",	--3102
		x"cf",	--3103
		x"01",	--3104
		x"f0",	--3105
		x"3e",	--3106
		x"f8",	--3107
		x"1b",	--3108
		x"02",	--3109
		x"1c",	--3110
		x"02",	--3111
		x"0c",	--3112
		x"e6",	--3113
		x"0b",	--3114
		x"16",	--3115
		x"1b",	--3116
		x"04",	--3117
		x"1f",	--3118
		x"06",	--3119
		x"1c",	--3120
		x"04",	--3121
		x"1e",	--3122
		x"06",	--3123
		x"0e",	--3124
		x"da",	--3125
		x"0f",	--3126
		x"02",	--3127
		x"0c",	--3128
		x"d6",	--3129
		x"0f",	--3130
		x"06",	--3131
		x"0e",	--3132
		x"02",	--3133
		x"0b",	--3134
		x"02",	--3135
		x"0e",	--3136
		x"d1",	--3137
		x"4d",	--3138
		x"ce",	--3139
		x"3e",	--3140
		x"d6",	--3141
		x"6c",	--3142
		x"d7",	--3143
		x"5e",	--3144
		x"01",	--3145
		x"5f",	--3146
		x"01",	--3147
		x"0e",	--3148
		x"c5",	--3149
		x"0d",	--3150
		x"0f",	--3151
		x"04",	--3152
		x"3d",	--3153
		x"03",	--3154
		x"3f",	--3155
		x"1f",	--3156
		x"0e",	--3157
		x"03",	--3158
		x"5d",	--3159
		x"3e",	--3160
		x"1e",	--3161
		x"0d",	--3162
		x"b0",	--3163
		x"22",	--3164
		x"3d",	--3165
		x"6d",	--3166
		x"02",	--3167
		x"3e",	--3168
		x"1e",	--3169
		x"5d",	--3170
		x"02",	--3171
		x"3f",	--3172
		x"1f",	--3173
		x"30",	--3174
		x"b0",	--3175
		x"9c",	--3176
		x"0f",	--3177
		x"30",	--3178
		x"0b",	--3179
		x"0b",	--3180
		x"0f",	--3181
		x"06",	--3182
		x"3b",	--3183
		x"03",	--3184
		x"3e",	--3185
		x"3f",	--3186
		x"1e",	--3187
		x"0f",	--3188
		x"0d",	--3189
		x"05",	--3190
		x"5b",	--3191
		x"3c",	--3192
		x"3d",	--3193
		x"1c",	--3194
		x"0d",	--3195
		x"b0",	--3196
		x"44",	--3197
		x"6b",	--3198
		x"04",	--3199
		x"3c",	--3200
		x"3d",	--3201
		x"1c",	--3202
		x"0d",	--3203
		x"5b",	--3204
		x"04",	--3205
		x"3e",	--3206
		x"3f",	--3207
		x"1e",	--3208
		x"0f",	--3209
		x"3b",	--3210
		x"30",	--3211
		x"b0",	--3212
		x"d6",	--3213
		x"0e",	--3214
		x"0f",	--3215
		x"30",	--3216
		x"7c",	--3217
		x"10",	--3218
		x"0d",	--3219
		x"0e",	--3220
		x"0f",	--3221
		x"0e",	--3222
		x"0e",	--3223
		x"02",	--3224
		x"0e",	--3225
		x"1f",	--3226
		x"1c",	--3227
		x"f8",	--3228
		x"30",	--3229
		x"b0",	--3230
		x"22",	--3231
		x"0f",	--3232
		x"30",	--3233
		x"0b",	--3234
		x"0a",	--3235
		x"09",	--3236
		x"79",	--3237
		x"20",	--3238
		x"0a",	--3239
		x"0b",	--3240
		x"0c",	--3241
		x"0d",	--3242
		x"0e",	--3243
		x"0f",	--3244
		x"0c",	--3245
		x"0d",	--3246
		x"0d",	--3247
		x"06",	--3248
		x"02",	--3249
		x"0c",	--3250
		x"03",	--3251
		x"0c",	--3252
		x"0d",	--3253
		x"1e",	--3254
		x"19",	--3255
		x"f2",	--3256
		x"39",	--3257
		x"3a",	--3258
		x"3b",	--3259
		x"30",	--3260
		x"b0",	--3261
		x"44",	--3262
		x"0e",	--3263
		x"0f",	--3264
		x"30",	--3265
		x"00",	--3266
		x"32",	--3267
		x"f0",	--3268
		x"fd",	--3269
		x"57",	--3270
		x"69",	--3271
		x"69",	--3272
		x"67",	--3273
		x"66",	--3274
		x"72",	--3275
		x"61",	--3276
		x"6e",	--3277
		x"77",	--3278
		x"2e",	--3279
		x"69",	--3280
		x"20",	--3281
		x"69",	--3282
		x"65",	--3283
		x"0a",	--3284
		x"57",	--3285
		x"20",	--3286
		x"68",	--3287
		x"75",	--3288
		x"64",	--3289
		x"6e",	--3290
		x"74",	--3291
		x"73",	--3292
		x"65",	--3293
		x"74",	--3294
		x"61",	--3295
		x"0d",	--3296
		x"00",	--3297
		x"72",	--3298
		x"6f",	--3299
		x"3a",	--3300
		x"6d",	--3301
		x"73",	--3302
		x"69",	--3303
		x"67",	--3304
		x"61",	--3305
		x"67",	--3306
		x"6d",	--3307
		x"6e",	--3308
		x"0d",	--3309
		x"00",	--3310
		x"6f",	--3311
		x"72",	--3312
		x"63",	--3313
		x"20",	--3314
		x"73",	--3315
		x"67",	--3316
		x"3a",	--3317
		x"0a",	--3318
		x"09",	--3319
		x"73",	--3320
		x"4c",	--3321
		x"46",	--3322
		x"20",	--3323
		x"49",	--3324
		x"48",	--3325
		x"0d",	--3326
		x"00",	--3327
		x"64",	--3328
		x"25",	--3329
		x"0d",	--3330
		x"00",	--3331
		x"77",	--3332
		x"25",	--3333
		x"20",	--3334
		x"77",	--3335
		x"25",	--3336
		x"0d",	--3337
		x"00",	--3338
		x"48",	--3339
		x"70",	--3340
		x"76",	--3341
		x"7e",	--3342
		x"86",	--3343
		x"8e",	--3344
		x"60",	--3345
		x"68",	--3346
		x"0d",	--3347
		x"3d",	--3348
		x"3d",	--3349
		x"3d",	--3350
		x"20",	--3351
		x"61",	--3352
		x"63",	--3353
		x"6c",	--3354
		x"4d",	--3355
		x"55",	--3356
		x"3d",	--3357
		x"3d",	--3358
		x"3d",	--3359
		x"0d",	--3360
		x"00",	--3361
		x"72",	--3362
		x"74",	--3363
		x"00",	--3364
		x"65",	--3365
		x"64",	--3366
		x"70",	--3367
		x"6d",	--3368
		x"65",	--3369
		x"63",	--3370
		x"64",	--3371
		x"72",	--3372
		x"62",	--3373
		x"6f",	--3374
		x"6c",	--3375
		x"61",	--3376
		x"65",	--3377
		x"00",	--3378
		x"0a",	--3379
		x"08",	--3380
		x"08",	--3381
		x"25",	--3382
		x"00",	--3383
		x"77",	--3384
		x"69",	--3385
		x"65",	--3386
		x"0d",	--3387
		x"65",	--3388
		x"72",	--3389
		x"72",	--3390
		x"20",	--3391
		x"69",	--3392
		x"73",	--3393
		x"6e",	--3394
		x"20",	--3395
		x"72",	--3396
		x"75",	--3397
		x"65",	--3398
		x"74",	--3399
		x"0a",	--3400
		x"63",	--3401
		x"72",	--3402
		x"65",	--3403
		x"74",	--3404
		x"75",	--3405
		x"61",	--3406
		x"65",	--3407
		x"0d",	--3408
		x"00",	--3409
		x"25",	--3410
		x"20",	--3411
		x"45",	--3412
		x"49",	--3413
		x"54",	--3414
		x"52",	--3415
		x"56",	--3416
		x"4c",	--3417
		x"45",	--3418
		x"0a",	--3419
		x"72",	--3420
		x"25",	--3421
		x"20",	--3422
		x"3d",	--3423
		x"64",	--3424
		x"0a",	--3425
		x"09",	--3426
		x"73",	--3427
		x"52",	--3428
		x"47",	--3429
		x"53",	--3430
		x"45",	--3431
		x"0d",	--3432
		x"00",	--3433
		x"65",	--3434
		x"64",	--3435
		x"0d",	--3436
		x"25",	--3437
		x"20",	--3438
		x"73",	--3439
		x"6e",	--3440
		x"74",	--3441
		x"61",	--3442
		x"6e",	--3443
		x"6d",	--3444
		x"65",	--3445
		x"0d",	--3446
		x"00",	--3447
		x"63",	--3448
		x"25",	--3449
		x"0d",	--3450
		x"00",	--3451
		x"63",	--3452
		x"20",	--3453
		x"6f",	--3454
		x"73",	--3455
		x"63",	--3456
		x"20",	--3457
		x"6f",	--3458
		x"6d",	--3459
		x"6e",	--3460
		x"0d",	--3461
		x"00",	--3462
		x"2c",	--3463
		x"5a",	--3464
		x"5a",	--3465
		x"5a",	--3466
		x"5a",	--3467
		x"5a",	--3468
		x"5a",	--3469
		x"5a",	--3470
		x"5a",	--3471
		x"5a",	--3472
		x"5a",	--3473
		x"5a",	--3474
		x"5a",	--3475
		x"5a",	--3476
		x"5a",	--3477
		x"5a",	--3478
		x"5a",	--3479
		x"5a",	--3480
		x"5a",	--3481
		x"5a",	--3482
		x"5a",	--3483
		x"5a",	--3484
		x"5a",	--3485
		x"5a",	--3486
		x"5a",	--3487
		x"5a",	--3488
		x"5a",	--3489
		x"5a",	--3490
		x"5a",	--3491
		x"1e",	--3492
		x"5a",	--3493
		x"5a",	--3494
		x"5a",	--3495
		x"5a",	--3496
		x"5a",	--3497
		x"5a",	--3498
		x"5a",	--3499
		x"5a",	--3500
		x"5a",	--3501
		x"5a",	--3502
		x"5a",	--3503
		x"5a",	--3504
		x"5a",	--3505
		x"5a",	--3506
		x"5a",	--3507
		x"5a",	--3508
		x"5a",	--3509
		x"5a",	--3510
		x"5a",	--3511
		x"5a",	--3512
		x"5a",	--3513
		x"5a",	--3514
		x"5a",	--3515
		x"5a",	--3516
		x"5a",	--3517
		x"5a",	--3518
		x"5a",	--3519
		x"5a",	--3520
		x"5a",	--3521
		x"5a",	--3522
		x"5a",	--3523
		x"10",	--3524
		x"02",	--3525
		x"f4",	--3526
		x"5a",	--3527
		x"5a",	--3528
		x"5a",	--3529
		x"5a",	--3530
		x"5a",	--3531
		x"5a",	--3532
		x"5a",	--3533
		x"dc",	--3534
		x"5a",	--3535
		x"ca",	--3536
		x"5a",	--3537
		x"5a",	--3538
		x"5a",	--3539
		x"5a",	--3540
		x"ae",	--3541
		x"5a",	--3542
		x"5a",	--3543
		x"5a",	--3544
		x"a0",	--3545
		x"8e",	--3546
		x"30",	--3547
		x"32",	--3548
		x"34",	--3549
		x"36",	--3550
		x"38",	--3551
		x"61",	--3552
		x"63",	--3553
		x"65",	--3554
		x"00",	--3555
		x"00",	--3556
		x"00",	--3557
		x"00",	--3558
		x"00",	--3559
		x"00",	--3560
		x"02",	--3561
		x"03",	--3562
		x"03",	--3563
		x"04",	--3564
		x"04",	--3565
		x"04",	--3566
		x"04",	--3567
		x"05",	--3568
		x"05",	--3569
		x"05",	--3570
		x"05",	--3571
		x"05",	--3572
		x"05",	--3573
		x"05",	--3574
		x"05",	--3575
		x"06",	--3576
		x"06",	--3577
		x"06",	--3578
		x"06",	--3579
		x"06",	--3580
		x"06",	--3581
		x"06",	--3582
		x"06",	--3583
		x"06",	--3584
		x"06",	--3585
		x"06",	--3586
		x"06",	--3587
		x"06",	--3588
		x"06",	--3589
		x"06",	--3590
		x"06",	--3591
		x"07",	--3592
		x"07",	--3593
		x"07",	--3594
		x"07",	--3595
		x"07",	--3596
		x"07",	--3597
		x"07",	--3598
		x"07",	--3599
		x"07",	--3600
		x"07",	--3601
		x"07",	--3602
		x"07",	--3603
		x"07",	--3604
		x"07",	--3605
		x"07",	--3606
		x"07",	--3607
		x"07",	--3608
		x"07",	--3609
		x"07",	--3610
		x"07",	--3611
		x"07",	--3612
		x"07",	--3613
		x"07",	--3614
		x"07",	--3615
		x"07",	--3616
		x"07",	--3617
		x"07",	--3618
		x"07",	--3619
		x"07",	--3620
		x"07",	--3621
		x"07",	--3622
		x"07",	--3623
		x"08",	--3624
		x"08",	--3625
		x"08",	--3626
		x"08",	--3627
		x"08",	--3628
		x"08",	--3629
		x"08",	--3630
		x"08",	--3631
		x"08",	--3632
		x"08",	--3633
		x"08",	--3634
		x"08",	--3635
		x"08",	--3636
		x"08",	--3637
		x"08",	--3638
		x"08",	--3639
		x"08",	--3640
		x"08",	--3641
		x"08",	--3642
		x"08",	--3643
		x"08",	--3644
		x"08",	--3645
		x"08",	--3646
		x"08",	--3647
		x"08",	--3648
		x"08",	--3649
		x"08",	--3650
		x"08",	--3651
		x"08",	--3652
		x"08",	--3653
		x"08",	--3654
		x"08",	--3655
		x"08",	--3656
		x"08",	--3657
		x"08",	--3658
		x"08",	--3659
		x"08",	--3660
		x"08",	--3661
		x"08",	--3662
		x"08",	--3663
		x"08",	--3664
		x"08",	--3665
		x"08",	--3666
		x"08",	--3667
		x"08",	--3668
		x"08",	--3669
		x"08",	--3670
		x"08",	--3671
		x"08",	--3672
		x"08",	--3673
		x"08",	--3674
		x"08",	--3675
		x"08",	--3676
		x"08",	--3677
		x"08",	--3678
		x"08",	--3679
		x"08",	--3680
		x"08",	--3681
		x"08",	--3682
		x"08",	--3683
		x"08",	--3684
		x"08",	--3685
		x"08",	--3686
		x"08",	--3687
		x"ff",	--3688
		x"68",	--3689
		x"6c",	--3690
		x"00",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"c2",	--4080
		x"c2",	--4081
		x"c2",	--4082
		x"c2",	--4083
		x"c2",	--4084
		x"c2",	--4085
		x"c2",	--4086
		x"36",	--4087
		x"ee",	--4088
		x"c2",	--4089
		x"c2",	--4090
		x"c2",	--4091
		x"c2",	--4092
		x"c2",	--4093
		x"c2",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"04",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"04",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fc",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"02",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"04",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"25",	--41
		x"43",	--42
		x"12",	--43
		x"eb",	--44
		x"12",	--45
		x"e6",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"fa",	--50
		x"12",	--51
		x"ea",	--52
		x"53",	--53
		x"40",	--54
		x"fa",	--55
		x"40",	--56
		x"e3",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"e6",	--61
		x"40",	--62
		x"fa",	--63
		x"40",	--64
		x"e4",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"e6",	--69
		x"40",	--70
		x"fa",	--71
		x"40",	--72
		x"e1",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"e6",	--77
		x"40",	--78
		x"fa",	--79
		x"40",	--80
		x"e2",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"e6",	--85
		x"40",	--86
		x"fa",	--87
		x"40",	--88
		x"e1",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"e6",	--93
		x"43",	--94
		x"43",	--95
		x"12",	--96
		x"e6",	--97
		x"43",	--98
		x"40",	--99
		x"4e",	--100
		x"40",	--101
		x"01",	--102
		x"41",	--103
		x"50",	--104
		x"00",	--105
		x"12",	--106
		x"e5",	--107
		x"41",	--108
		x"50",	--109
		x"00",	--110
		x"12",	--111
		x"e5",	--112
		x"43",	--113
		x"40",	--114
		x"4e",	--115
		x"40",	--116
		x"01",	--117
		x"41",	--118
		x"52",	--119
		x"12",	--120
		x"e5",	--121
		x"41",	--122
		x"52",	--123
		x"12",	--124
		x"e5",	--125
		x"41",	--126
		x"52",	--127
		x"41",	--128
		x"50",	--129
		x"00",	--130
		x"12",	--131
		x"e1",	--132
		x"40",	--133
		x"01",	--134
		x"41",	--135
		x"53",	--136
		x"12",	--137
		x"e8",	--138
		x"40",	--139
		x"01",	--140
		x"41",	--141
		x"12",	--142
		x"e8",	--143
		x"41",	--144
		x"41",	--145
		x"53",	--146
		x"12",	--147
		x"e2",	--148
		x"12",	--149
		x"e7",	--150
		x"43",	--151
		x"40",	--152
		x"e3",	--153
		x"12",	--154
		x"e7",	--155
		x"43",	--156
		x"12",	--157
		x"e7",	--158
		x"40",	--159
		x"ff",	--160
		x"00",	--161
		x"d2",	--162
		x"43",	--163
		x"12",	--164
		x"eb",	--165
		x"93",	--166
		x"27",	--167
		x"12",	--168
		x"eb",	--169
		x"92",	--170
		x"24",	--171
		x"90",	--172
		x"00",	--173
		x"20",	--174
		x"12",	--175
		x"fa",	--176
		x"12",	--177
		x"ea",	--178
		x"53",	--179
		x"40",	--180
		x"00",	--181
		x"51",	--182
		x"5f",	--183
		x"43",	--184
		x"00",	--185
		x"4f",	--186
		x"41",	--187
		x"00",	--188
		x"12",	--189
		x"e6",	--190
		x"43",	--191
		x"3f",	--192
		x"93",	--193
		x"27",	--194
		x"53",	--195
		x"12",	--196
		x"fa",	--197
		x"12",	--198
		x"ea",	--199
		x"53",	--200
		x"3f",	--201
		x"90",	--202
		x"00",	--203
		x"2f",	--204
		x"4f",	--205
		x"11",	--206
		x"12",	--207
		x"12",	--208
		x"fa",	--209
		x"4f",	--210
		x"00",	--211
		x"12",	--212
		x"ea",	--213
		x"52",	--214
		x"40",	--215
		x"00",	--216
		x"51",	--217
		x"5b",	--218
		x"41",	--219
		x"00",	--220
		x"4f",	--221
		x"00",	--222
		x"53",	--223
		x"3f",	--224
		x"40",	--225
		x"f9",	--226
		x"40",	--227
		x"e0",	--228
		x"01",	--229
		x"42",	--230
		x"01",	--231
		x"40",	--232
		x"02",	--233
		x"01",	--234
		x"12",	--235
		x"f9",	--236
		x"12",	--237
		x"ea",	--238
		x"43",	--239
		x"01",	--240
		x"40",	--241
		x"f9",	--242
		x"00",	--243
		x"12",	--244
		x"ea",	--245
		x"53",	--246
		x"43",	--247
		x"41",	--248
		x"4f",	--249
		x"02",	--250
		x"4e",	--251
		x"02",	--252
		x"41",	--253
		x"12",	--254
		x"12",	--255
		x"83",	--256
		x"4e",	--257
		x"93",	--258
		x"24",	--259
		x"38",	--260
		x"41",	--261
		x"4b",	--262
		x"00",	--263
		x"12",	--264
		x"e4",	--265
		x"4f",	--266
		x"41",	--267
		x"4b",	--268
		x"00",	--269
		x"12",	--270
		x"e4",	--271
		x"4f",	--272
		x"12",	--273
		x"12",	--274
		x"12",	--275
		x"f9",	--276
		x"12",	--277
		x"ea",	--278
		x"50",	--279
		x"00",	--280
		x"4a",	--281
		x"43",	--282
		x"12",	--283
		x"f3",	--284
		x"43",	--285
		x"40",	--286
		x"42",	--287
		x"12",	--288
		x"f1",	--289
		x"4e",	--290
		x"4f",	--291
		x"42",	--292
		x"02",	--293
		x"12",	--294
		x"e5",	--295
		x"4b",	--296
		x"43",	--297
		x"12",	--298
		x"f3",	--299
		x"43",	--300
		x"40",	--301
		x"42",	--302
		x"12",	--303
		x"f1",	--304
		x"4e",	--305
		x"4f",	--306
		x"42",	--307
		x"02",	--308
		x"12",	--309
		x"e5",	--310
		x"43",	--311
		x"53",	--312
		x"41",	--313
		x"41",	--314
		x"41",	--315
		x"12",	--316
		x"f9",	--317
		x"12",	--318
		x"ea",	--319
		x"40",	--320
		x"f9",	--321
		x"00",	--322
		x"12",	--323
		x"ea",	--324
		x"4b",	--325
		x"00",	--326
		x"12",	--327
		x"f9",	--328
		x"12",	--329
		x"ea",	--330
		x"52",	--331
		x"43",	--332
		x"3f",	--333
		x"42",	--334
		x"02",	--335
		x"4f",	--336
		x"42",	--337
		x"02",	--338
		x"4f",	--339
		x"12",	--340
		x"12",	--341
		x"00",	--342
		x"12",	--343
		x"12",	--344
		x"00",	--345
		x"12",	--346
		x"fa",	--347
		x"12",	--348
		x"ea",	--349
		x"50",	--350
		x"00",	--351
		x"41",	--352
		x"4f",	--353
		x"02",	--354
		x"4e",	--355
		x"02",	--356
		x"41",	--357
		x"12",	--358
		x"83",	--359
		x"4e",	--360
		x"43",	--361
		x"00",	--362
		x"93",	--363
		x"24",	--364
		x"93",	--365
		x"02",	--366
		x"24",	--367
		x"43",	--368
		x"02",	--369
		x"41",	--370
		x"4b",	--371
		x"00",	--372
		x"12",	--373
		x"e4",	--374
		x"4f",	--375
		x"42",	--376
		x"02",	--377
		x"12",	--378
		x"e7",	--379
		x"43",	--380
		x"53",	--381
		x"41",	--382
		x"41",	--383
		x"93",	--384
		x"02",	--385
		x"24",	--386
		x"43",	--387
		x"02",	--388
		x"42",	--389
		x"02",	--390
		x"12",	--391
		x"e7",	--392
		x"43",	--393
		x"53",	--394
		x"41",	--395
		x"41",	--396
		x"43",	--397
		x"12",	--398
		x"e2",	--399
		x"43",	--400
		x"53",	--401
		x"41",	--402
		x"41",	--403
		x"43",	--404
		x"40",	--405
		x"e2",	--406
		x"12",	--407
		x"e7",	--408
		x"4f",	--409
		x"02",	--410
		x"3f",	--411
		x"42",	--412
		x"02",	--413
		x"92",	--414
		x"2c",	--415
		x"4e",	--416
		x"5f",	--417
		x"4f",	--418
		x"fa",	--419
		x"43",	--420
		x"00",	--421
		x"90",	--422
		x"00",	--423
		x"38",	--424
		x"43",	--425
		x"02",	--426
		x"41",	--427
		x"53",	--428
		x"4e",	--429
		x"02",	--430
		x"41",	--431
		x"40",	--432
		x"00",	--433
		x"00",	--434
		x"3f",	--435
		x"40",	--436
		x"00",	--437
		x"00",	--438
		x"3f",	--439
		x"42",	--440
		x"00",	--441
		x"3f",	--442
		x"40",	--443
		x"00",	--444
		x"00",	--445
		x"3f",	--446
		x"40",	--447
		x"00",	--448
		x"00",	--449
		x"3f",	--450
		x"40",	--451
		x"00",	--452
		x"00",	--453
		x"3f",	--454
		x"40",	--455
		x"00",	--456
		x"00",	--457
		x"3f",	--458
		x"42",	--459
		x"00",	--460
		x"4e",	--461
		x"be",	--462
		x"20",	--463
		x"df",	--464
		x"00",	--465
		x"41",	--466
		x"cf",	--467
		x"00",	--468
		x"41",	--469
		x"12",	--470
		x"12",	--471
		x"83",	--472
		x"4f",	--473
		x"4e",	--474
		x"12",	--475
		x"fa",	--476
		x"12",	--477
		x"ea",	--478
		x"53",	--479
		x"90",	--480
		x"00",	--481
		x"38",	--482
		x"41",	--483
		x"4b",	--484
		x"00",	--485
		x"12",	--486
		x"e4",	--487
		x"4f",	--488
		x"41",	--489
		x"4b",	--490
		x"00",	--491
		x"12",	--492
		x"e4",	--493
		x"4f",	--494
		x"12",	--495
		x"12",	--496
		x"12",	--497
		x"fa",	--498
		x"12",	--499
		x"ea",	--500
		x"50",	--501
		x"00",	--502
		x"4b",	--503
		x"00",	--504
		x"43",	--505
		x"53",	--506
		x"41",	--507
		x"41",	--508
		x"41",	--509
		x"12",	--510
		x"fa",	--511
		x"12",	--512
		x"ea",	--513
		x"40",	--514
		x"fa",	--515
		x"00",	--516
		x"12",	--517
		x"ea",	--518
		x"4b",	--519
		x"00",	--520
		x"12",	--521
		x"fa",	--522
		x"12",	--523
		x"ea",	--524
		x"52",	--525
		x"43",	--526
		x"3f",	--527
		x"12",	--528
		x"83",	--529
		x"4e",	--530
		x"93",	--531
		x"24",	--532
		x"38",	--533
		x"12",	--534
		x"fa",	--535
		x"12",	--536
		x"ea",	--537
		x"53",	--538
		x"41",	--539
		x"4b",	--540
		x"00",	--541
		x"12",	--542
		x"e4",	--543
		x"12",	--544
		x"12",	--545
		x"12",	--546
		x"fa",	--547
		x"12",	--548
		x"ea",	--549
		x"50",	--550
		x"00",	--551
		x"43",	--552
		x"53",	--553
		x"41",	--554
		x"41",	--555
		x"12",	--556
		x"fa",	--557
		x"12",	--558
		x"ea",	--559
		x"40",	--560
		x"fa",	--561
		x"00",	--562
		x"12",	--563
		x"ea",	--564
		x"4b",	--565
		x"00",	--566
		x"12",	--567
		x"fa",	--568
		x"12",	--569
		x"ea",	--570
		x"52",	--571
		x"43",	--572
		x"3f",	--573
		x"12",	--574
		x"12",	--575
		x"43",	--576
		x"00",	--577
		x"4f",	--578
		x"93",	--579
		x"24",	--580
		x"53",	--581
		x"43",	--582
		x"43",	--583
		x"3c",	--584
		x"90",	--585
		x"00",	--586
		x"2c",	--587
		x"5c",	--588
		x"5c",	--589
		x"5c",	--590
		x"5c",	--591
		x"11",	--592
		x"5d",	--593
		x"50",	--594
		x"ff",	--595
		x"43",	--596
		x"4f",	--597
		x"93",	--598
		x"24",	--599
		x"90",	--600
		x"00",	--601
		x"24",	--602
		x"4d",	--603
		x"50",	--604
		x"ff",	--605
		x"93",	--606
		x"23",	--607
		x"90",	--608
		x"00",	--609
		x"2c",	--610
		x"5c",	--611
		x"4c",	--612
		x"5b",	--613
		x"5b",	--614
		x"5b",	--615
		x"11",	--616
		x"5d",	--617
		x"50",	--618
		x"ff",	--619
		x"4f",	--620
		x"93",	--621
		x"23",	--622
		x"43",	--623
		x"00",	--624
		x"4c",	--625
		x"41",	--626
		x"41",	--627
		x"41",	--628
		x"43",	--629
		x"3f",	--630
		x"4d",	--631
		x"50",	--632
		x"ff",	--633
		x"90",	--634
		x"00",	--635
		x"2c",	--636
		x"5c",	--637
		x"5c",	--638
		x"5c",	--639
		x"5c",	--640
		x"11",	--641
		x"5d",	--642
		x"50",	--643
		x"ff",	--644
		x"43",	--645
		x"3f",	--646
		x"4d",	--647
		x"50",	--648
		x"ff",	--649
		x"90",	--650
		x"00",	--651
		x"2c",	--652
		x"5c",	--653
		x"5c",	--654
		x"5c",	--655
		x"5c",	--656
		x"11",	--657
		x"5d",	--658
		x"50",	--659
		x"ff",	--660
		x"43",	--661
		x"3f",	--662
		x"11",	--663
		x"12",	--664
		x"12",	--665
		x"fa",	--666
		x"12",	--667
		x"ea",	--668
		x"52",	--669
		x"43",	--670
		x"4c",	--671
		x"41",	--672
		x"41",	--673
		x"41",	--674
		x"43",	--675
		x"3f",	--676
		x"12",	--677
		x"12",	--678
		x"4e",	--679
		x"4c",	--680
		x"4e",	--681
		x"00",	--682
		x"4d",	--683
		x"00",	--684
		x"4c",	--685
		x"00",	--686
		x"4d",	--687
		x"43",	--688
		x"40",	--689
		x"36",	--690
		x"40",	--691
		x"01",	--692
		x"12",	--693
		x"f8",	--694
		x"4e",	--695
		x"00",	--696
		x"12",	--697
		x"c2",	--698
		x"43",	--699
		x"4a",	--700
		x"01",	--701
		x"40",	--702
		x"00",	--703
		x"01",	--704
		x"42",	--705
		x"01",	--706
		x"00",	--707
		x"41",	--708
		x"43",	--709
		x"41",	--710
		x"41",	--711
		x"41",	--712
		x"12",	--713
		x"12",	--714
		x"12",	--715
		x"43",	--716
		x"00",	--717
		x"40",	--718
		x"3f",	--719
		x"00",	--720
		x"4f",	--721
		x"4b",	--722
		x"00",	--723
		x"43",	--724
		x"12",	--725
		x"f3",	--726
		x"43",	--727
		x"40",	--728
		x"3f",	--729
		x"12",	--730
		x"ef",	--731
		x"4e",	--732
		x"4f",	--733
		x"4b",	--734
		x"00",	--735
		x"43",	--736
		x"12",	--737
		x"f3",	--738
		x"4e",	--739
		x"4f",	--740
		x"48",	--741
		x"49",	--742
		x"12",	--743
		x"ee",	--744
		x"12",	--745
		x"eb",	--746
		x"4e",	--747
		x"00",	--748
		x"43",	--749
		x"00",	--750
		x"41",	--751
		x"41",	--752
		x"41",	--753
		x"41",	--754
		x"12",	--755
		x"12",	--756
		x"12",	--757
		x"4d",	--758
		x"4e",	--759
		x"4d",	--760
		x"00",	--761
		x"4e",	--762
		x"00",	--763
		x"4f",	--764
		x"49",	--765
		x"00",	--766
		x"43",	--767
		x"12",	--768
		x"f3",	--769
		x"4e",	--770
		x"4f",	--771
		x"4a",	--772
		x"4b",	--773
		x"12",	--774
		x"ef",	--775
		x"4e",	--776
		x"4f",	--777
		x"49",	--778
		x"00",	--779
		x"43",	--780
		x"12",	--781
		x"f3",	--782
		x"4e",	--783
		x"4f",	--784
		x"4a",	--785
		x"4b",	--786
		x"12",	--787
		x"ee",	--788
		x"12",	--789
		x"eb",	--790
		x"4e",	--791
		x"00",	--792
		x"41",	--793
		x"41",	--794
		x"41",	--795
		x"41",	--796
		x"12",	--797
		x"12",	--798
		x"93",	--799
		x"02",	--800
		x"38",	--801
		x"40",	--802
		x"02",	--803
		x"43",	--804
		x"12",	--805
		x"4b",	--806
		x"ff",	--807
		x"11",	--808
		x"12",	--809
		x"12",	--810
		x"fa",	--811
		x"12",	--812
		x"ea",	--813
		x"50",	--814
		x"00",	--815
		x"53",	--816
		x"50",	--817
		x"00",	--818
		x"92",	--819
		x"02",	--820
		x"3b",	--821
		x"43",	--822
		x"41",	--823
		x"41",	--824
		x"41",	--825
		x"42",	--826
		x"02",	--827
		x"90",	--828
		x"00",	--829
		x"34",	--830
		x"4e",	--831
		x"5f",	--832
		x"5e",	--833
		x"5f",	--834
		x"50",	--835
		x"02",	--836
		x"40",	--837
		x"00",	--838
		x"00",	--839
		x"40",	--840
		x"e6",	--841
		x"00",	--842
		x"40",	--843
		x"02",	--844
		x"00",	--845
		x"53",	--846
		x"4e",	--847
		x"02",	--848
		x"41",	--849
		x"12",	--850
		x"42",	--851
		x"02",	--852
		x"90",	--853
		x"00",	--854
		x"34",	--855
		x"4b",	--856
		x"5c",	--857
		x"5b",	--858
		x"5c",	--859
		x"50",	--860
		x"02",	--861
		x"4f",	--862
		x"00",	--863
		x"4e",	--864
		x"00",	--865
		x"4d",	--866
		x"00",	--867
		x"53",	--868
		x"4b",	--869
		x"02",	--870
		x"43",	--871
		x"41",	--872
		x"41",	--873
		x"43",	--874
		x"3f",	--875
		x"12",	--876
		x"50",	--877
		x"ff",	--878
		x"42",	--879
		x"02",	--880
		x"93",	--881
		x"38",	--882
		x"92",	--883
		x"02",	--884
		x"24",	--885
		x"40",	--886
		x"02",	--887
		x"43",	--888
		x"3c",	--889
		x"50",	--890
		x"00",	--891
		x"9f",	--892
		x"ff",	--893
		x"24",	--894
		x"53",	--895
		x"9b",	--896
		x"23",	--897
		x"12",	--898
		x"fa",	--899
		x"12",	--900
		x"ea",	--901
		x"53",	--902
		x"43",	--903
		x"50",	--904
		x"00",	--905
		x"41",	--906
		x"41",	--907
		x"43",	--908
		x"4e",	--909
		x"00",	--910
		x"4e",	--911
		x"93",	--912
		x"24",	--913
		x"53",	--914
		x"43",	--915
		x"3c",	--916
		x"4e",	--917
		x"93",	--918
		x"24",	--919
		x"53",	--920
		x"92",	--921
		x"34",	--922
		x"90",	--923
		x"00",	--924
		x"23",	--925
		x"43",	--926
		x"ff",	--927
		x"4f",	--928
		x"5d",	--929
		x"51",	--930
		x"4e",	--931
		x"00",	--932
		x"53",	--933
		x"4e",	--934
		x"93",	--935
		x"23",	--936
		x"4c",	--937
		x"5e",	--938
		x"5e",	--939
		x"5c",	--940
		x"50",	--941
		x"02",	--942
		x"41",	--943
		x"12",	--944
		x"00",	--945
		x"50",	--946
		x"00",	--947
		x"41",	--948
		x"41",	--949
		x"43",	--950
		x"3f",	--951
		x"d0",	--952
		x"02",	--953
		x"01",	--954
		x"40",	--955
		x"0b",	--956
		x"01",	--957
		x"43",	--958
		x"41",	--959
		x"12",	--960
		x"4f",	--961
		x"42",	--962
		x"02",	--963
		x"90",	--964
		x"00",	--965
		x"34",	--966
		x"4f",	--967
		x"5c",	--968
		x"4c",	--969
		x"5d",	--970
		x"5d",	--971
		x"5c",	--972
		x"50",	--973
		x"02",	--974
		x"43",	--975
		x"00",	--976
		x"43",	--977
		x"00",	--978
		x"4b",	--979
		x"00",	--980
		x"4e",	--981
		x"00",	--982
		x"4f",	--983
		x"53",	--984
		x"4e",	--985
		x"02",	--986
		x"41",	--987
		x"41",	--988
		x"43",	--989
		x"3f",	--990
		x"5f",	--991
		x"4f",	--992
		x"5d",	--993
		x"5d",	--994
		x"5f",	--995
		x"50",	--996
		x"02",	--997
		x"43",	--998
		x"00",	--999
		x"4e",	--1000
		x"00",	--1001
		x"43",	--1002
		x"00",	--1003
		x"43",	--1004
		x"41",	--1005
		x"5f",	--1006
		x"4f",	--1007
		x"5e",	--1008
		x"5e",	--1009
		x"5f",	--1010
		x"43",	--1011
		x"02",	--1012
		x"43",	--1013
		x"41",	--1014
		x"12",	--1015
		x"12",	--1016
		x"12",	--1017
		x"12",	--1018
		x"12",	--1019
		x"12",	--1020
		x"93",	--1021
		x"02",	--1022
		x"38",	--1023
		x"40",	--1024
		x"02",	--1025
		x"43",	--1026
		x"3c",	--1027
		x"53",	--1028
		x"4f",	--1029
		x"00",	--1030
		x"53",	--1031
		x"50",	--1032
		x"00",	--1033
		x"92",	--1034
		x"02",	--1035
		x"34",	--1036
		x"93",	--1037
		x"ff",	--1038
		x"27",	--1039
		x"4b",	--1040
		x"9b",	--1041
		x"00",	--1042
		x"2b",	--1043
		x"43",	--1044
		x"00",	--1045
		x"4b",	--1046
		x"00",	--1047
		x"12",	--1048
		x"00",	--1049
		x"53",	--1050
		x"50",	--1051
		x"00",	--1052
		x"92",	--1053
		x"02",	--1054
		x"3b",	--1055
		x"f0",	--1056
		x"ff",	--1057
		x"01",	--1058
		x"41",	--1059
		x"41",	--1060
		x"41",	--1061
		x"41",	--1062
		x"41",	--1063
		x"41",	--1064
		x"13",	--1065
		x"4e",	--1066
		x"00",	--1067
		x"43",	--1068
		x"41",	--1069
		x"4f",	--1070
		x"4f",	--1071
		x"41",	--1072
		x"42",	--1073
		x"00",	--1074
		x"f2",	--1075
		x"23",	--1076
		x"4f",	--1077
		x"00",	--1078
		x"43",	--1079
		x"41",	--1080
		x"f0",	--1081
		x"00",	--1082
		x"4f",	--1083
		x"fb",	--1084
		x"11",	--1085
		x"12",	--1086
		x"e8",	--1087
		x"41",	--1088
		x"12",	--1089
		x"4f",	--1090
		x"4f",	--1091
		x"11",	--1092
		x"11",	--1093
		x"11",	--1094
		x"11",	--1095
		x"4e",	--1096
		x"12",	--1097
		x"e8",	--1098
		x"4b",	--1099
		x"12",	--1100
		x"e8",	--1101
		x"41",	--1102
		x"41",	--1103
		x"12",	--1104
		x"12",	--1105
		x"4f",	--1106
		x"40",	--1107
		x"00",	--1108
		x"4a",	--1109
		x"4b",	--1110
		x"f0",	--1111
		x"00",	--1112
		x"24",	--1113
		x"11",	--1114
		x"53",	--1115
		x"23",	--1116
		x"f3",	--1117
		x"24",	--1118
		x"40",	--1119
		x"00",	--1120
		x"12",	--1121
		x"e8",	--1122
		x"53",	--1123
		x"93",	--1124
		x"23",	--1125
		x"41",	--1126
		x"41",	--1127
		x"41",	--1128
		x"40",	--1129
		x"00",	--1130
		x"3f",	--1131
		x"12",	--1132
		x"4f",	--1133
		x"4f",	--1134
		x"10",	--1135
		x"11",	--1136
		x"4e",	--1137
		x"12",	--1138
		x"e8",	--1139
		x"4b",	--1140
		x"12",	--1141
		x"e8",	--1142
		x"41",	--1143
		x"41",	--1144
		x"12",	--1145
		x"12",	--1146
		x"4e",	--1147
		x"4f",	--1148
		x"4f",	--1149
		x"10",	--1150
		x"11",	--1151
		x"4d",	--1152
		x"12",	--1153
		x"e8",	--1154
		x"4b",	--1155
		x"12",	--1156
		x"e8",	--1157
		x"4b",	--1158
		x"4a",	--1159
		x"10",	--1160
		x"10",	--1161
		x"ec",	--1162
		x"ec",	--1163
		x"4d",	--1164
		x"12",	--1165
		x"e8",	--1166
		x"4a",	--1167
		x"12",	--1168
		x"e8",	--1169
		x"41",	--1170
		x"41",	--1171
		x"41",	--1172
		x"12",	--1173
		x"12",	--1174
		x"12",	--1175
		x"4f",	--1176
		x"93",	--1177
		x"24",	--1178
		x"4e",	--1179
		x"53",	--1180
		x"43",	--1181
		x"4a",	--1182
		x"5b",	--1183
		x"4d",	--1184
		x"11",	--1185
		x"12",	--1186
		x"e8",	--1187
		x"99",	--1188
		x"24",	--1189
		x"53",	--1190
		x"b0",	--1191
		x"00",	--1192
		x"20",	--1193
		x"40",	--1194
		x"00",	--1195
		x"12",	--1196
		x"e8",	--1197
		x"3f",	--1198
		x"40",	--1199
		x"00",	--1200
		x"12",	--1201
		x"e8",	--1202
		x"3f",	--1203
		x"41",	--1204
		x"41",	--1205
		x"41",	--1206
		x"41",	--1207
		x"12",	--1208
		x"12",	--1209
		x"12",	--1210
		x"4f",	--1211
		x"93",	--1212
		x"24",	--1213
		x"4e",	--1214
		x"53",	--1215
		x"43",	--1216
		x"4a",	--1217
		x"11",	--1218
		x"12",	--1219
		x"e8",	--1220
		x"99",	--1221
		x"24",	--1222
		x"53",	--1223
		x"b0",	--1224
		x"00",	--1225
		x"23",	--1226
		x"40",	--1227
		x"00",	--1228
		x"12",	--1229
		x"e8",	--1230
		x"4a",	--1231
		x"11",	--1232
		x"12",	--1233
		x"e8",	--1234
		x"99",	--1235
		x"23",	--1236
		x"41",	--1237
		x"41",	--1238
		x"41",	--1239
		x"41",	--1240
		x"12",	--1241
		x"12",	--1242
		x"12",	--1243
		x"50",	--1244
		x"ff",	--1245
		x"4f",	--1246
		x"93",	--1247
		x"38",	--1248
		x"90",	--1249
		x"00",	--1250
		x"38",	--1251
		x"43",	--1252
		x"41",	--1253
		x"59",	--1254
		x"40",	--1255
		x"00",	--1256
		x"4b",	--1257
		x"12",	--1258
		x"f8",	--1259
		x"50",	--1260
		x"00",	--1261
		x"4f",	--1262
		x"00",	--1263
		x"53",	--1264
		x"40",	--1265
		x"00",	--1266
		x"4b",	--1267
		x"12",	--1268
		x"f8",	--1269
		x"4f",	--1270
		x"90",	--1271
		x"00",	--1272
		x"37",	--1273
		x"49",	--1274
		x"53",	--1275
		x"51",	--1276
		x"40",	--1277
		x"00",	--1278
		x"4b",	--1279
		x"12",	--1280
		x"f8",	--1281
		x"50",	--1282
		x"00",	--1283
		x"4f",	--1284
		x"00",	--1285
		x"53",	--1286
		x"41",	--1287
		x"5a",	--1288
		x"4f",	--1289
		x"11",	--1290
		x"12",	--1291
		x"e8",	--1292
		x"93",	--1293
		x"23",	--1294
		x"50",	--1295
		x"00",	--1296
		x"41",	--1297
		x"41",	--1298
		x"41",	--1299
		x"41",	--1300
		x"40",	--1301
		x"00",	--1302
		x"12",	--1303
		x"e8",	--1304
		x"e3",	--1305
		x"53",	--1306
		x"3f",	--1307
		x"43",	--1308
		x"43",	--1309
		x"3f",	--1310
		x"12",	--1311
		x"12",	--1312
		x"12",	--1313
		x"41",	--1314
		x"52",	--1315
		x"4b",	--1316
		x"49",	--1317
		x"93",	--1318
		x"20",	--1319
		x"3c",	--1320
		x"11",	--1321
		x"12",	--1322
		x"e8",	--1323
		x"49",	--1324
		x"4a",	--1325
		x"53",	--1326
		x"4a",	--1327
		x"00",	--1328
		x"93",	--1329
		x"24",	--1330
		x"90",	--1331
		x"00",	--1332
		x"23",	--1333
		x"49",	--1334
		x"53",	--1335
		x"49",	--1336
		x"00",	--1337
		x"50",	--1338
		x"ff",	--1339
		x"90",	--1340
		x"00",	--1341
		x"2f",	--1342
		x"4f",	--1343
		x"5f",	--1344
		x"4f",	--1345
		x"fb",	--1346
		x"41",	--1347
		x"41",	--1348
		x"41",	--1349
		x"41",	--1350
		x"4b",	--1351
		x"52",	--1352
		x"4b",	--1353
		x"00",	--1354
		x"4b",	--1355
		x"12",	--1356
		x"e9",	--1357
		x"49",	--1358
		x"3f",	--1359
		x"4b",	--1360
		x"53",	--1361
		x"4b",	--1362
		x"12",	--1363
		x"e8",	--1364
		x"49",	--1365
		x"3f",	--1366
		x"4b",	--1367
		x"53",	--1368
		x"4f",	--1369
		x"49",	--1370
		x"93",	--1371
		x"27",	--1372
		x"53",	--1373
		x"11",	--1374
		x"12",	--1375
		x"e8",	--1376
		x"49",	--1377
		x"93",	--1378
		x"23",	--1379
		x"3f",	--1380
		x"4b",	--1381
		x"52",	--1382
		x"4b",	--1383
		x"00",	--1384
		x"4b",	--1385
		x"12",	--1386
		x"e9",	--1387
		x"49",	--1388
		x"3f",	--1389
		x"4b",	--1390
		x"53",	--1391
		x"4b",	--1392
		x"4e",	--1393
		x"10",	--1394
		x"11",	--1395
		x"10",	--1396
		x"11",	--1397
		x"12",	--1398
		x"e8",	--1399
		x"49",	--1400
		x"3f",	--1401
		x"4b",	--1402
		x"53",	--1403
		x"4b",	--1404
		x"12",	--1405
		x"e9",	--1406
		x"49",	--1407
		x"3f",	--1408
		x"4b",	--1409
		x"53",	--1410
		x"4b",	--1411
		x"12",	--1412
		x"e8",	--1413
		x"49",	--1414
		x"3f",	--1415
		x"4b",	--1416
		x"53",	--1417
		x"4b",	--1418
		x"12",	--1419
		x"e8",	--1420
		x"49",	--1421
		x"3f",	--1422
		x"4b",	--1423
		x"53",	--1424
		x"4b",	--1425
		x"12",	--1426
		x"e8",	--1427
		x"49",	--1428
		x"3f",	--1429
		x"40",	--1430
		x"00",	--1431
		x"12",	--1432
		x"e8",	--1433
		x"3f",	--1434
		x"12",	--1435
		x"12",	--1436
		x"42",	--1437
		x"02",	--1438
		x"42",	--1439
		x"00",	--1440
		x"04",	--1441
		x"42",	--1442
		x"02",	--1443
		x"90",	--1444
		x"00",	--1445
		x"34",	--1446
		x"53",	--1447
		x"02",	--1448
		x"42",	--1449
		x"02",	--1450
		x"42",	--1451
		x"02",	--1452
		x"9f",	--1453
		x"20",	--1454
		x"53",	--1455
		x"02",	--1456
		x"40",	--1457
		x"00",	--1458
		x"00",	--1459
		x"41",	--1460
		x"41",	--1461
		x"c0",	--1462
		x"00",	--1463
		x"00",	--1464
		x"13",	--1465
		x"43",	--1466
		x"02",	--1467
		x"3f",	--1468
		x"40",	--1469
		x"09",	--1470
		x"00",	--1471
		x"40",	--1472
		x"00",	--1473
		x"00",	--1474
		x"41",	--1475
		x"42",	--1476
		x"02",	--1477
		x"42",	--1478
		x"02",	--1479
		x"9f",	--1480
		x"38",	--1481
		x"42",	--1482
		x"02",	--1483
		x"82",	--1484
		x"02",	--1485
		x"41",	--1486
		x"42",	--1487
		x"02",	--1488
		x"42",	--1489
		x"02",	--1490
		x"40",	--1491
		x"00",	--1492
		x"8d",	--1493
		x"8e",	--1494
		x"41",	--1495
		x"42",	--1496
		x"02",	--1497
		x"4f",	--1498
		x"04",	--1499
		x"42",	--1500
		x"02",	--1501
		x"42",	--1502
		x"02",	--1503
		x"9e",	--1504
		x"24",	--1505
		x"42",	--1506
		x"02",	--1507
		x"90",	--1508
		x"00",	--1509
		x"38",	--1510
		x"43",	--1511
		x"02",	--1512
		x"41",	--1513
		x"53",	--1514
		x"02",	--1515
		x"41",	--1516
		x"43",	--1517
		x"41",	--1518
		x"12",	--1519
		x"12",	--1520
		x"4e",	--1521
		x"4f",	--1522
		x"43",	--1523
		x"40",	--1524
		x"4f",	--1525
		x"12",	--1526
		x"f2",	--1527
		x"93",	--1528
		x"34",	--1529
		x"4a",	--1530
		x"4b",	--1531
		x"12",	--1532
		x"f3",	--1533
		x"41",	--1534
		x"41",	--1535
		x"41",	--1536
		x"43",	--1537
		x"40",	--1538
		x"4f",	--1539
		x"4a",	--1540
		x"4b",	--1541
		x"12",	--1542
		x"ee",	--1543
		x"12",	--1544
		x"f3",	--1545
		x"53",	--1546
		x"60",	--1547
		x"80",	--1548
		x"41",	--1549
		x"41",	--1550
		x"41",	--1551
		x"12",	--1552
		x"12",	--1553
		x"12",	--1554
		x"12",	--1555
		x"12",	--1556
		x"12",	--1557
		x"12",	--1558
		x"12",	--1559
		x"50",	--1560
		x"ff",	--1561
		x"4d",	--1562
		x"4f",	--1563
		x"93",	--1564
		x"28",	--1565
		x"4e",	--1566
		x"93",	--1567
		x"28",	--1568
		x"92",	--1569
		x"20",	--1570
		x"40",	--1571
		x"ee",	--1572
		x"92",	--1573
		x"24",	--1574
		x"93",	--1575
		x"24",	--1576
		x"93",	--1577
		x"24",	--1578
		x"4f",	--1579
		x"00",	--1580
		x"00",	--1581
		x"4e",	--1582
		x"00",	--1583
		x"4f",	--1584
		x"00",	--1585
		x"4f",	--1586
		x"00",	--1587
		x"4e",	--1588
		x"00",	--1589
		x"4e",	--1590
		x"00",	--1591
		x"41",	--1592
		x"8b",	--1593
		x"4c",	--1594
		x"93",	--1595
		x"38",	--1596
		x"90",	--1597
		x"00",	--1598
		x"34",	--1599
		x"93",	--1600
		x"38",	--1601
		x"46",	--1602
		x"00",	--1603
		x"47",	--1604
		x"00",	--1605
		x"49",	--1606
		x"f0",	--1607
		x"00",	--1608
		x"24",	--1609
		x"46",	--1610
		x"47",	--1611
		x"c3",	--1612
		x"10",	--1613
		x"10",	--1614
		x"53",	--1615
		x"23",	--1616
		x"4a",	--1617
		x"00",	--1618
		x"4b",	--1619
		x"00",	--1620
		x"43",	--1621
		x"43",	--1622
		x"f0",	--1623
		x"00",	--1624
		x"24",	--1625
		x"5c",	--1626
		x"6d",	--1627
		x"53",	--1628
		x"23",	--1629
		x"53",	--1630
		x"63",	--1631
		x"f6",	--1632
		x"f7",	--1633
		x"43",	--1634
		x"43",	--1635
		x"93",	--1636
		x"20",	--1637
		x"93",	--1638
		x"24",	--1639
		x"41",	--1640
		x"00",	--1641
		x"41",	--1642
		x"00",	--1643
		x"da",	--1644
		x"db",	--1645
		x"4f",	--1646
		x"00",	--1647
		x"9e",	--1648
		x"00",	--1649
		x"20",	--1650
		x"4f",	--1651
		x"00",	--1652
		x"41",	--1653
		x"00",	--1654
		x"46",	--1655
		x"47",	--1656
		x"54",	--1657
		x"65",	--1658
		x"4e",	--1659
		x"00",	--1660
		x"4f",	--1661
		x"00",	--1662
		x"40",	--1663
		x"00",	--1664
		x"00",	--1665
		x"93",	--1666
		x"38",	--1667
		x"48",	--1668
		x"50",	--1669
		x"00",	--1670
		x"41",	--1671
		x"41",	--1672
		x"41",	--1673
		x"41",	--1674
		x"41",	--1675
		x"41",	--1676
		x"41",	--1677
		x"41",	--1678
		x"41",	--1679
		x"91",	--1680
		x"38",	--1681
		x"4b",	--1682
		x"00",	--1683
		x"43",	--1684
		x"43",	--1685
		x"4f",	--1686
		x"00",	--1687
		x"9e",	--1688
		x"00",	--1689
		x"27",	--1690
		x"93",	--1691
		x"24",	--1692
		x"46",	--1693
		x"47",	--1694
		x"84",	--1695
		x"75",	--1696
		x"93",	--1697
		x"38",	--1698
		x"43",	--1699
		x"00",	--1700
		x"41",	--1701
		x"00",	--1702
		x"4e",	--1703
		x"00",	--1704
		x"4f",	--1705
		x"00",	--1706
		x"4e",	--1707
		x"4f",	--1708
		x"53",	--1709
		x"63",	--1710
		x"90",	--1711
		x"3f",	--1712
		x"28",	--1713
		x"90",	--1714
		x"40",	--1715
		x"2c",	--1716
		x"93",	--1717
		x"2c",	--1718
		x"48",	--1719
		x"00",	--1720
		x"53",	--1721
		x"5e",	--1722
		x"6f",	--1723
		x"4b",	--1724
		x"53",	--1725
		x"4e",	--1726
		x"4f",	--1727
		x"53",	--1728
		x"63",	--1729
		x"90",	--1730
		x"3f",	--1731
		x"2b",	--1732
		x"24",	--1733
		x"4e",	--1734
		x"00",	--1735
		x"4f",	--1736
		x"00",	--1737
		x"4a",	--1738
		x"00",	--1739
		x"40",	--1740
		x"00",	--1741
		x"00",	--1742
		x"93",	--1743
		x"37",	--1744
		x"4e",	--1745
		x"4f",	--1746
		x"f3",	--1747
		x"f3",	--1748
		x"c3",	--1749
		x"10",	--1750
		x"10",	--1751
		x"4c",	--1752
		x"4d",	--1753
		x"de",	--1754
		x"df",	--1755
		x"4a",	--1756
		x"00",	--1757
		x"4b",	--1758
		x"00",	--1759
		x"53",	--1760
		x"00",	--1761
		x"48",	--1762
		x"3f",	--1763
		x"93",	--1764
		x"23",	--1765
		x"4f",	--1766
		x"00",	--1767
		x"4f",	--1768
		x"00",	--1769
		x"00",	--1770
		x"4f",	--1771
		x"00",	--1772
		x"00",	--1773
		x"4f",	--1774
		x"00",	--1775
		x"00",	--1776
		x"4e",	--1777
		x"00",	--1778
		x"ff",	--1779
		x"00",	--1780
		x"4e",	--1781
		x"00",	--1782
		x"4d",	--1783
		x"3f",	--1784
		x"43",	--1785
		x"43",	--1786
		x"3f",	--1787
		x"e3",	--1788
		x"53",	--1789
		x"90",	--1790
		x"00",	--1791
		x"37",	--1792
		x"3f",	--1793
		x"93",	--1794
		x"2b",	--1795
		x"3f",	--1796
		x"44",	--1797
		x"45",	--1798
		x"86",	--1799
		x"77",	--1800
		x"3f",	--1801
		x"4e",	--1802
		x"3f",	--1803
		x"43",	--1804
		x"00",	--1805
		x"41",	--1806
		x"00",	--1807
		x"e3",	--1808
		x"e3",	--1809
		x"53",	--1810
		x"63",	--1811
		x"4e",	--1812
		x"00",	--1813
		x"4f",	--1814
		x"00",	--1815
		x"3f",	--1816
		x"93",	--1817
		x"27",	--1818
		x"59",	--1819
		x"00",	--1820
		x"44",	--1821
		x"00",	--1822
		x"45",	--1823
		x"00",	--1824
		x"49",	--1825
		x"f0",	--1826
		x"00",	--1827
		x"24",	--1828
		x"4d",	--1829
		x"44",	--1830
		x"45",	--1831
		x"c3",	--1832
		x"10",	--1833
		x"10",	--1834
		x"53",	--1835
		x"23",	--1836
		x"4c",	--1837
		x"00",	--1838
		x"4d",	--1839
		x"00",	--1840
		x"43",	--1841
		x"43",	--1842
		x"f0",	--1843
		x"00",	--1844
		x"24",	--1845
		x"5c",	--1846
		x"6d",	--1847
		x"53",	--1848
		x"23",	--1849
		x"53",	--1850
		x"63",	--1851
		x"f4",	--1852
		x"f5",	--1853
		x"43",	--1854
		x"43",	--1855
		x"93",	--1856
		x"20",	--1857
		x"93",	--1858
		x"20",	--1859
		x"43",	--1860
		x"43",	--1861
		x"41",	--1862
		x"00",	--1863
		x"41",	--1864
		x"00",	--1865
		x"da",	--1866
		x"db",	--1867
		x"3f",	--1868
		x"43",	--1869
		x"43",	--1870
		x"3f",	--1871
		x"92",	--1872
		x"23",	--1873
		x"9e",	--1874
		x"00",	--1875
		x"00",	--1876
		x"27",	--1877
		x"40",	--1878
		x"fb",	--1879
		x"3f",	--1880
		x"50",	--1881
		x"ff",	--1882
		x"4e",	--1883
		x"00",	--1884
		x"4f",	--1885
		x"00",	--1886
		x"4c",	--1887
		x"00",	--1888
		x"4d",	--1889
		x"00",	--1890
		x"41",	--1891
		x"50",	--1892
		x"00",	--1893
		x"41",	--1894
		x"52",	--1895
		x"12",	--1896
		x"f6",	--1897
		x"41",	--1898
		x"50",	--1899
		x"00",	--1900
		x"41",	--1901
		x"12",	--1902
		x"f6",	--1903
		x"41",	--1904
		x"52",	--1905
		x"41",	--1906
		x"50",	--1907
		x"00",	--1908
		x"41",	--1909
		x"50",	--1910
		x"00",	--1911
		x"12",	--1912
		x"ec",	--1913
		x"12",	--1914
		x"f4",	--1915
		x"50",	--1916
		x"00",	--1917
		x"41",	--1918
		x"50",	--1919
		x"ff",	--1920
		x"4e",	--1921
		x"00",	--1922
		x"4f",	--1923
		x"00",	--1924
		x"4c",	--1925
		x"00",	--1926
		x"4d",	--1927
		x"00",	--1928
		x"41",	--1929
		x"50",	--1930
		x"00",	--1931
		x"41",	--1932
		x"52",	--1933
		x"12",	--1934
		x"f6",	--1935
		x"41",	--1936
		x"50",	--1937
		x"00",	--1938
		x"41",	--1939
		x"12",	--1940
		x"f6",	--1941
		x"e3",	--1942
		x"00",	--1943
		x"41",	--1944
		x"52",	--1945
		x"41",	--1946
		x"50",	--1947
		x"00",	--1948
		x"41",	--1949
		x"50",	--1950
		x"00",	--1951
		x"12",	--1952
		x"ec",	--1953
		x"12",	--1954
		x"f4",	--1955
		x"50",	--1956
		x"00",	--1957
		x"41",	--1958
		x"12",	--1959
		x"12",	--1960
		x"12",	--1961
		x"12",	--1962
		x"12",	--1963
		x"12",	--1964
		x"12",	--1965
		x"12",	--1966
		x"50",	--1967
		x"ff",	--1968
		x"4e",	--1969
		x"00",	--1970
		x"4f",	--1971
		x"00",	--1972
		x"4c",	--1973
		x"00",	--1974
		x"4d",	--1975
		x"00",	--1976
		x"41",	--1977
		x"50",	--1978
		x"00",	--1979
		x"41",	--1980
		x"52",	--1981
		x"12",	--1982
		x"f6",	--1983
		x"41",	--1984
		x"50",	--1985
		x"00",	--1986
		x"41",	--1987
		x"12",	--1988
		x"f6",	--1989
		x"41",	--1990
		x"00",	--1991
		x"93",	--1992
		x"28",	--1993
		x"41",	--1994
		x"00",	--1995
		x"93",	--1996
		x"28",	--1997
		x"92",	--1998
		x"24",	--1999
		x"92",	--2000
		x"24",	--2001
		x"93",	--2002
		x"24",	--2003
		x"93",	--2004
		x"24",	--2005
		x"41",	--2006
		x"00",	--2007
		x"41",	--2008
		x"00",	--2009
		x"41",	--2010
		x"00",	--2011
		x"41",	--2012
		x"00",	--2013
		x"40",	--2014
		x"00",	--2015
		x"43",	--2016
		x"43",	--2017
		x"43",	--2018
		x"43",	--2019
		x"43",	--2020
		x"00",	--2021
		x"43",	--2022
		x"00",	--2023
		x"43",	--2024
		x"43",	--2025
		x"4c",	--2026
		x"00",	--2027
		x"3c",	--2028
		x"58",	--2029
		x"69",	--2030
		x"c3",	--2031
		x"10",	--2032
		x"10",	--2033
		x"53",	--2034
		x"00",	--2035
		x"24",	--2036
		x"b3",	--2037
		x"24",	--2038
		x"58",	--2039
		x"69",	--2040
		x"56",	--2041
		x"67",	--2042
		x"43",	--2043
		x"43",	--2044
		x"99",	--2045
		x"28",	--2046
		x"24",	--2047
		x"43",	--2048
		x"43",	--2049
		x"5c",	--2050
		x"6d",	--2051
		x"56",	--2052
		x"67",	--2053
		x"93",	--2054
		x"37",	--2055
		x"d3",	--2056
		x"d3",	--2057
		x"3f",	--2058
		x"98",	--2059
		x"2b",	--2060
		x"3f",	--2061
		x"4a",	--2062
		x"00",	--2063
		x"4b",	--2064
		x"00",	--2065
		x"4f",	--2066
		x"41",	--2067
		x"00",	--2068
		x"51",	--2069
		x"00",	--2070
		x"4a",	--2071
		x"53",	--2072
		x"46",	--2073
		x"00",	--2074
		x"43",	--2075
		x"91",	--2076
		x"00",	--2077
		x"00",	--2078
		x"24",	--2079
		x"4d",	--2080
		x"00",	--2081
		x"93",	--2082
		x"38",	--2083
		x"90",	--2084
		x"40",	--2085
		x"2c",	--2086
		x"41",	--2087
		x"00",	--2088
		x"53",	--2089
		x"41",	--2090
		x"00",	--2091
		x"41",	--2092
		x"00",	--2093
		x"4d",	--2094
		x"5e",	--2095
		x"6f",	--2096
		x"93",	--2097
		x"38",	--2098
		x"5a",	--2099
		x"6b",	--2100
		x"53",	--2101
		x"90",	--2102
		x"40",	--2103
		x"2b",	--2104
		x"4a",	--2105
		x"00",	--2106
		x"4b",	--2107
		x"00",	--2108
		x"4c",	--2109
		x"00",	--2110
		x"4e",	--2111
		x"4f",	--2112
		x"f0",	--2113
		x"00",	--2114
		x"f3",	--2115
		x"90",	--2116
		x"00",	--2117
		x"24",	--2118
		x"4e",	--2119
		x"00",	--2120
		x"4f",	--2121
		x"00",	--2122
		x"40",	--2123
		x"00",	--2124
		x"00",	--2125
		x"41",	--2126
		x"52",	--2127
		x"12",	--2128
		x"f4",	--2129
		x"50",	--2130
		x"00",	--2131
		x"41",	--2132
		x"41",	--2133
		x"41",	--2134
		x"41",	--2135
		x"41",	--2136
		x"41",	--2137
		x"41",	--2138
		x"41",	--2139
		x"41",	--2140
		x"d3",	--2141
		x"d3",	--2142
		x"3f",	--2143
		x"50",	--2144
		x"00",	--2145
		x"4a",	--2146
		x"b3",	--2147
		x"24",	--2148
		x"41",	--2149
		x"00",	--2150
		x"41",	--2151
		x"00",	--2152
		x"c3",	--2153
		x"10",	--2154
		x"10",	--2155
		x"4c",	--2156
		x"4d",	--2157
		x"d3",	--2158
		x"d0",	--2159
		x"80",	--2160
		x"46",	--2161
		x"00",	--2162
		x"47",	--2163
		x"00",	--2164
		x"c3",	--2165
		x"10",	--2166
		x"10",	--2167
		x"53",	--2168
		x"93",	--2169
		x"3b",	--2170
		x"48",	--2171
		x"00",	--2172
		x"3f",	--2173
		x"93",	--2174
		x"24",	--2175
		x"43",	--2176
		x"91",	--2177
		x"00",	--2178
		x"00",	--2179
		x"24",	--2180
		x"4f",	--2181
		x"00",	--2182
		x"41",	--2183
		x"50",	--2184
		x"00",	--2185
		x"3f",	--2186
		x"93",	--2187
		x"23",	--2188
		x"4e",	--2189
		x"4f",	--2190
		x"f0",	--2191
		x"00",	--2192
		x"f3",	--2193
		x"93",	--2194
		x"23",	--2195
		x"93",	--2196
		x"23",	--2197
		x"93",	--2198
		x"00",	--2199
		x"20",	--2200
		x"93",	--2201
		x"00",	--2202
		x"27",	--2203
		x"50",	--2204
		x"00",	--2205
		x"63",	--2206
		x"f0",	--2207
		x"ff",	--2208
		x"f3",	--2209
		x"3f",	--2210
		x"43",	--2211
		x"3f",	--2212
		x"43",	--2213
		x"3f",	--2214
		x"43",	--2215
		x"91",	--2216
		x"00",	--2217
		x"00",	--2218
		x"24",	--2219
		x"4f",	--2220
		x"00",	--2221
		x"41",	--2222
		x"50",	--2223
		x"00",	--2224
		x"3f",	--2225
		x"43",	--2226
		x"3f",	--2227
		x"93",	--2228
		x"23",	--2229
		x"40",	--2230
		x"fb",	--2231
		x"3f",	--2232
		x"12",	--2233
		x"12",	--2234
		x"12",	--2235
		x"12",	--2236
		x"12",	--2237
		x"50",	--2238
		x"ff",	--2239
		x"4e",	--2240
		x"00",	--2241
		x"4f",	--2242
		x"00",	--2243
		x"4c",	--2244
		x"00",	--2245
		x"4d",	--2246
		x"00",	--2247
		x"41",	--2248
		x"50",	--2249
		x"00",	--2250
		x"41",	--2251
		x"52",	--2252
		x"12",	--2253
		x"f6",	--2254
		x"41",	--2255
		x"52",	--2256
		x"41",	--2257
		x"12",	--2258
		x"f6",	--2259
		x"41",	--2260
		x"00",	--2261
		x"93",	--2262
		x"28",	--2263
		x"41",	--2264
		x"00",	--2265
		x"93",	--2266
		x"28",	--2267
		x"e1",	--2268
		x"00",	--2269
		x"00",	--2270
		x"92",	--2271
		x"24",	--2272
		x"93",	--2273
		x"24",	--2274
		x"92",	--2275
		x"24",	--2276
		x"93",	--2277
		x"24",	--2278
		x"41",	--2279
		x"00",	--2280
		x"81",	--2281
		x"00",	--2282
		x"4d",	--2283
		x"00",	--2284
		x"41",	--2285
		x"00",	--2286
		x"41",	--2287
		x"00",	--2288
		x"41",	--2289
		x"00",	--2290
		x"41",	--2291
		x"00",	--2292
		x"99",	--2293
		x"2c",	--2294
		x"5e",	--2295
		x"6f",	--2296
		x"53",	--2297
		x"4d",	--2298
		x"00",	--2299
		x"40",	--2300
		x"00",	--2301
		x"43",	--2302
		x"40",	--2303
		x"40",	--2304
		x"43",	--2305
		x"43",	--2306
		x"3c",	--2307
		x"dc",	--2308
		x"dd",	--2309
		x"88",	--2310
		x"79",	--2311
		x"c3",	--2312
		x"10",	--2313
		x"10",	--2314
		x"5e",	--2315
		x"6f",	--2316
		x"53",	--2317
		x"24",	--2318
		x"99",	--2319
		x"2b",	--2320
		x"23",	--2321
		x"98",	--2322
		x"2b",	--2323
		x"3f",	--2324
		x"9f",	--2325
		x"2b",	--2326
		x"98",	--2327
		x"2f",	--2328
		x"3f",	--2329
		x"4a",	--2330
		x"4b",	--2331
		x"f0",	--2332
		x"00",	--2333
		x"f3",	--2334
		x"90",	--2335
		x"00",	--2336
		x"24",	--2337
		x"4a",	--2338
		x"00",	--2339
		x"4b",	--2340
		x"00",	--2341
		x"41",	--2342
		x"50",	--2343
		x"00",	--2344
		x"12",	--2345
		x"f4",	--2346
		x"50",	--2347
		x"00",	--2348
		x"41",	--2349
		x"41",	--2350
		x"41",	--2351
		x"41",	--2352
		x"41",	--2353
		x"41",	--2354
		x"42",	--2355
		x"00",	--2356
		x"41",	--2357
		x"50",	--2358
		x"00",	--2359
		x"3f",	--2360
		x"9e",	--2361
		x"23",	--2362
		x"40",	--2363
		x"fb",	--2364
		x"3f",	--2365
		x"93",	--2366
		x"23",	--2367
		x"4a",	--2368
		x"4b",	--2369
		x"f0",	--2370
		x"00",	--2371
		x"f3",	--2372
		x"93",	--2373
		x"23",	--2374
		x"93",	--2375
		x"23",	--2376
		x"93",	--2377
		x"20",	--2378
		x"93",	--2379
		x"27",	--2380
		x"50",	--2381
		x"00",	--2382
		x"63",	--2383
		x"f0",	--2384
		x"ff",	--2385
		x"f3",	--2386
		x"3f",	--2387
		x"43",	--2388
		x"00",	--2389
		x"43",	--2390
		x"00",	--2391
		x"43",	--2392
		x"00",	--2393
		x"41",	--2394
		x"50",	--2395
		x"00",	--2396
		x"3f",	--2397
		x"41",	--2398
		x"52",	--2399
		x"3f",	--2400
		x"50",	--2401
		x"ff",	--2402
		x"4e",	--2403
		x"00",	--2404
		x"4f",	--2405
		x"00",	--2406
		x"4c",	--2407
		x"00",	--2408
		x"4d",	--2409
		x"00",	--2410
		x"41",	--2411
		x"50",	--2412
		x"00",	--2413
		x"41",	--2414
		x"52",	--2415
		x"12",	--2416
		x"f6",	--2417
		x"41",	--2418
		x"52",	--2419
		x"41",	--2420
		x"12",	--2421
		x"f6",	--2422
		x"93",	--2423
		x"00",	--2424
		x"28",	--2425
		x"93",	--2426
		x"00",	--2427
		x"28",	--2428
		x"41",	--2429
		x"52",	--2430
		x"41",	--2431
		x"50",	--2432
		x"00",	--2433
		x"12",	--2434
		x"f7",	--2435
		x"50",	--2436
		x"00",	--2437
		x"41",	--2438
		x"43",	--2439
		x"3f",	--2440
		x"50",	--2441
		x"ff",	--2442
		x"4e",	--2443
		x"00",	--2444
		x"4f",	--2445
		x"00",	--2446
		x"41",	--2447
		x"52",	--2448
		x"41",	--2449
		x"12",	--2450
		x"f6",	--2451
		x"41",	--2452
		x"00",	--2453
		x"93",	--2454
		x"24",	--2455
		x"28",	--2456
		x"92",	--2457
		x"24",	--2458
		x"41",	--2459
		x"00",	--2460
		x"93",	--2461
		x"38",	--2462
		x"90",	--2463
		x"00",	--2464
		x"38",	--2465
		x"93",	--2466
		x"00",	--2467
		x"20",	--2468
		x"43",	--2469
		x"40",	--2470
		x"7f",	--2471
		x"50",	--2472
		x"00",	--2473
		x"41",	--2474
		x"41",	--2475
		x"00",	--2476
		x"41",	--2477
		x"00",	--2478
		x"40",	--2479
		x"00",	--2480
		x"8d",	--2481
		x"4c",	--2482
		x"f0",	--2483
		x"00",	--2484
		x"20",	--2485
		x"93",	--2486
		x"00",	--2487
		x"27",	--2488
		x"e3",	--2489
		x"e3",	--2490
		x"53",	--2491
		x"63",	--2492
		x"50",	--2493
		x"00",	--2494
		x"41",	--2495
		x"43",	--2496
		x"43",	--2497
		x"50",	--2498
		x"00",	--2499
		x"41",	--2500
		x"c3",	--2501
		x"10",	--2502
		x"10",	--2503
		x"53",	--2504
		x"23",	--2505
		x"3f",	--2506
		x"43",	--2507
		x"40",	--2508
		x"80",	--2509
		x"50",	--2510
		x"00",	--2511
		x"41",	--2512
		x"12",	--2513
		x"12",	--2514
		x"12",	--2515
		x"12",	--2516
		x"82",	--2517
		x"4e",	--2518
		x"4f",	--2519
		x"43",	--2520
		x"00",	--2521
		x"93",	--2522
		x"20",	--2523
		x"93",	--2524
		x"20",	--2525
		x"43",	--2526
		x"00",	--2527
		x"41",	--2528
		x"12",	--2529
		x"f4",	--2530
		x"52",	--2531
		x"41",	--2532
		x"41",	--2533
		x"41",	--2534
		x"41",	--2535
		x"41",	--2536
		x"40",	--2537
		x"00",	--2538
		x"00",	--2539
		x"40",	--2540
		x"00",	--2541
		x"00",	--2542
		x"4a",	--2543
		x"00",	--2544
		x"4b",	--2545
		x"00",	--2546
		x"4a",	--2547
		x"4b",	--2548
		x"12",	--2549
		x"f4",	--2550
		x"53",	--2551
		x"93",	--2552
		x"38",	--2553
		x"27",	--2554
		x"4a",	--2555
		x"00",	--2556
		x"4b",	--2557
		x"00",	--2558
		x"4f",	--2559
		x"f0",	--2560
		x"00",	--2561
		x"20",	--2562
		x"40",	--2563
		x"00",	--2564
		x"8f",	--2565
		x"4e",	--2566
		x"00",	--2567
		x"3f",	--2568
		x"51",	--2569
		x"00",	--2570
		x"00",	--2571
		x"61",	--2572
		x"00",	--2573
		x"00",	--2574
		x"53",	--2575
		x"23",	--2576
		x"3f",	--2577
		x"4f",	--2578
		x"e3",	--2579
		x"53",	--2580
		x"43",	--2581
		x"43",	--2582
		x"4e",	--2583
		x"f0",	--2584
		x"00",	--2585
		x"24",	--2586
		x"5c",	--2587
		x"6d",	--2588
		x"53",	--2589
		x"23",	--2590
		x"53",	--2591
		x"63",	--2592
		x"fa",	--2593
		x"fb",	--2594
		x"43",	--2595
		x"43",	--2596
		x"93",	--2597
		x"20",	--2598
		x"93",	--2599
		x"20",	--2600
		x"43",	--2601
		x"43",	--2602
		x"f0",	--2603
		x"00",	--2604
		x"20",	--2605
		x"48",	--2606
		x"49",	--2607
		x"da",	--2608
		x"db",	--2609
		x"4d",	--2610
		x"00",	--2611
		x"4e",	--2612
		x"00",	--2613
		x"40",	--2614
		x"00",	--2615
		x"8f",	--2616
		x"4e",	--2617
		x"00",	--2618
		x"3f",	--2619
		x"c3",	--2620
		x"10",	--2621
		x"10",	--2622
		x"53",	--2623
		x"23",	--2624
		x"3f",	--2625
		x"12",	--2626
		x"12",	--2627
		x"12",	--2628
		x"93",	--2629
		x"2c",	--2630
		x"90",	--2631
		x"01",	--2632
		x"28",	--2633
		x"40",	--2634
		x"00",	--2635
		x"43",	--2636
		x"42",	--2637
		x"4e",	--2638
		x"4f",	--2639
		x"49",	--2640
		x"93",	--2641
		x"20",	--2642
		x"50",	--2643
		x"fb",	--2644
		x"4c",	--2645
		x"43",	--2646
		x"8e",	--2647
		x"7f",	--2648
		x"4a",	--2649
		x"41",	--2650
		x"41",	--2651
		x"41",	--2652
		x"41",	--2653
		x"90",	--2654
		x"01",	--2655
		x"28",	--2656
		x"42",	--2657
		x"43",	--2658
		x"40",	--2659
		x"00",	--2660
		x"4e",	--2661
		x"4f",	--2662
		x"49",	--2663
		x"93",	--2664
		x"27",	--2665
		x"c3",	--2666
		x"10",	--2667
		x"10",	--2668
		x"53",	--2669
		x"23",	--2670
		x"3f",	--2671
		x"40",	--2672
		x"00",	--2673
		x"43",	--2674
		x"40",	--2675
		x"00",	--2676
		x"3f",	--2677
		x"40",	--2678
		x"00",	--2679
		x"43",	--2680
		x"43",	--2681
		x"3f",	--2682
		x"12",	--2683
		x"12",	--2684
		x"12",	--2685
		x"12",	--2686
		x"12",	--2687
		x"4f",	--2688
		x"4f",	--2689
		x"00",	--2690
		x"4f",	--2691
		x"00",	--2692
		x"4d",	--2693
		x"00",	--2694
		x"4d",	--2695
		x"93",	--2696
		x"28",	--2697
		x"92",	--2698
		x"24",	--2699
		x"93",	--2700
		x"24",	--2701
		x"93",	--2702
		x"24",	--2703
		x"4d",	--2704
		x"00",	--2705
		x"90",	--2706
		x"ff",	--2707
		x"38",	--2708
		x"90",	--2709
		x"00",	--2710
		x"34",	--2711
		x"4e",	--2712
		x"4f",	--2713
		x"f0",	--2714
		x"00",	--2715
		x"f3",	--2716
		x"90",	--2717
		x"00",	--2718
		x"24",	--2719
		x"50",	--2720
		x"00",	--2721
		x"63",	--2722
		x"93",	--2723
		x"38",	--2724
		x"4b",	--2725
		x"50",	--2726
		x"00",	--2727
		x"c3",	--2728
		x"10",	--2729
		x"10",	--2730
		x"c3",	--2731
		x"10",	--2732
		x"10",	--2733
		x"c3",	--2734
		x"10",	--2735
		x"10",	--2736
		x"c3",	--2737
		x"10",	--2738
		x"10",	--2739
		x"c3",	--2740
		x"10",	--2741
		x"10",	--2742
		x"c3",	--2743
		x"10",	--2744
		x"10",	--2745
		x"c3",	--2746
		x"10",	--2747
		x"10",	--2748
		x"f3",	--2749
		x"f0",	--2750
		x"00",	--2751
		x"4d",	--2752
		x"3c",	--2753
		x"93",	--2754
		x"23",	--2755
		x"43",	--2756
		x"43",	--2757
		x"43",	--2758
		x"4d",	--2759
		x"5d",	--2760
		x"5d",	--2761
		x"5d",	--2762
		x"5d",	--2763
		x"5d",	--2764
		x"5d",	--2765
		x"5d",	--2766
		x"4f",	--2767
		x"f0",	--2768
		x"00",	--2769
		x"dd",	--2770
		x"4a",	--2771
		x"11",	--2772
		x"43",	--2773
		x"10",	--2774
		x"4c",	--2775
		x"df",	--2776
		x"4d",	--2777
		x"41",	--2778
		x"41",	--2779
		x"41",	--2780
		x"41",	--2781
		x"41",	--2782
		x"41",	--2783
		x"93",	--2784
		x"23",	--2785
		x"4e",	--2786
		x"4f",	--2787
		x"f0",	--2788
		x"00",	--2789
		x"f3",	--2790
		x"93",	--2791
		x"20",	--2792
		x"93",	--2793
		x"27",	--2794
		x"50",	--2795
		x"00",	--2796
		x"63",	--2797
		x"3f",	--2798
		x"c3",	--2799
		x"10",	--2800
		x"10",	--2801
		x"4b",	--2802
		x"50",	--2803
		x"00",	--2804
		x"3f",	--2805
		x"43",	--2806
		x"43",	--2807
		x"43",	--2808
		x"3f",	--2809
		x"d3",	--2810
		x"d0",	--2811
		x"00",	--2812
		x"f3",	--2813
		x"f0",	--2814
		x"00",	--2815
		x"43",	--2816
		x"3f",	--2817
		x"40",	--2818
		x"ff",	--2819
		x"8b",	--2820
		x"90",	--2821
		x"00",	--2822
		x"34",	--2823
		x"4e",	--2824
		x"4f",	--2825
		x"47",	--2826
		x"f0",	--2827
		x"00",	--2828
		x"24",	--2829
		x"c3",	--2830
		x"10",	--2831
		x"10",	--2832
		x"53",	--2833
		x"23",	--2834
		x"43",	--2835
		x"43",	--2836
		x"f0",	--2837
		x"00",	--2838
		x"24",	--2839
		x"58",	--2840
		x"69",	--2841
		x"53",	--2842
		x"23",	--2843
		x"53",	--2844
		x"63",	--2845
		x"fe",	--2846
		x"ff",	--2847
		x"43",	--2848
		x"43",	--2849
		x"93",	--2850
		x"20",	--2851
		x"93",	--2852
		x"20",	--2853
		x"43",	--2854
		x"43",	--2855
		x"4e",	--2856
		x"4f",	--2857
		x"dc",	--2858
		x"dd",	--2859
		x"48",	--2860
		x"49",	--2861
		x"f0",	--2862
		x"00",	--2863
		x"f3",	--2864
		x"90",	--2865
		x"00",	--2866
		x"24",	--2867
		x"50",	--2868
		x"00",	--2869
		x"63",	--2870
		x"48",	--2871
		x"49",	--2872
		x"c3",	--2873
		x"10",	--2874
		x"10",	--2875
		x"c3",	--2876
		x"10",	--2877
		x"10",	--2878
		x"c3",	--2879
		x"10",	--2880
		x"10",	--2881
		x"c3",	--2882
		x"10",	--2883
		x"10",	--2884
		x"c3",	--2885
		x"10",	--2886
		x"10",	--2887
		x"c3",	--2888
		x"10",	--2889
		x"10",	--2890
		x"c3",	--2891
		x"10",	--2892
		x"10",	--2893
		x"f3",	--2894
		x"f0",	--2895
		x"00",	--2896
		x"43",	--2897
		x"90",	--2898
		x"40",	--2899
		x"2f",	--2900
		x"43",	--2901
		x"3f",	--2902
		x"43",	--2903
		x"43",	--2904
		x"3f",	--2905
		x"93",	--2906
		x"23",	--2907
		x"48",	--2908
		x"49",	--2909
		x"f0",	--2910
		x"00",	--2911
		x"f3",	--2912
		x"93",	--2913
		x"24",	--2914
		x"50",	--2915
		x"00",	--2916
		x"63",	--2917
		x"3f",	--2918
		x"93",	--2919
		x"27",	--2920
		x"3f",	--2921
		x"12",	--2922
		x"12",	--2923
		x"4f",	--2924
		x"4f",	--2925
		x"00",	--2926
		x"f0",	--2927
		x"00",	--2928
		x"4f",	--2929
		x"00",	--2930
		x"c3",	--2931
		x"10",	--2932
		x"c3",	--2933
		x"10",	--2934
		x"c3",	--2935
		x"10",	--2936
		x"c3",	--2937
		x"10",	--2938
		x"c3",	--2939
		x"10",	--2940
		x"c3",	--2941
		x"10",	--2942
		x"c3",	--2943
		x"10",	--2944
		x"4d",	--2945
		x"4f",	--2946
		x"00",	--2947
		x"b0",	--2948
		x"00",	--2949
		x"43",	--2950
		x"6f",	--2951
		x"4f",	--2952
		x"00",	--2953
		x"93",	--2954
		x"20",	--2955
		x"93",	--2956
		x"24",	--2957
		x"40",	--2958
		x"ff",	--2959
		x"00",	--2960
		x"4a",	--2961
		x"4b",	--2962
		x"5c",	--2963
		x"6d",	--2964
		x"5c",	--2965
		x"6d",	--2966
		x"5c",	--2967
		x"6d",	--2968
		x"5c",	--2969
		x"6d",	--2970
		x"5c",	--2971
		x"6d",	--2972
		x"5c",	--2973
		x"6d",	--2974
		x"5c",	--2975
		x"6d",	--2976
		x"40",	--2977
		x"00",	--2978
		x"00",	--2979
		x"90",	--2980
		x"40",	--2981
		x"2c",	--2982
		x"40",	--2983
		x"ff",	--2984
		x"5c",	--2985
		x"6d",	--2986
		x"4f",	--2987
		x"53",	--2988
		x"90",	--2989
		x"40",	--2990
		x"2b",	--2991
		x"4a",	--2992
		x"00",	--2993
		x"4c",	--2994
		x"00",	--2995
		x"4d",	--2996
		x"00",	--2997
		x"41",	--2998
		x"41",	--2999
		x"41",	--3000
		x"90",	--3001
		x"00",	--3002
		x"24",	--3003
		x"50",	--3004
		x"ff",	--3005
		x"4d",	--3006
		x"00",	--3007
		x"40",	--3008
		x"00",	--3009
		x"00",	--3010
		x"4a",	--3011
		x"4b",	--3012
		x"5c",	--3013
		x"6d",	--3014
		x"5c",	--3015
		x"6d",	--3016
		x"5c",	--3017
		x"6d",	--3018
		x"5c",	--3019
		x"6d",	--3020
		x"5c",	--3021
		x"6d",	--3022
		x"5c",	--3023
		x"6d",	--3024
		x"5c",	--3025
		x"6d",	--3026
		x"4c",	--3027
		x"4d",	--3028
		x"d3",	--3029
		x"d0",	--3030
		x"40",	--3031
		x"4a",	--3032
		x"00",	--3033
		x"4b",	--3034
		x"00",	--3035
		x"41",	--3036
		x"41",	--3037
		x"41",	--3038
		x"93",	--3039
		x"23",	--3040
		x"43",	--3041
		x"00",	--3042
		x"41",	--3043
		x"41",	--3044
		x"41",	--3045
		x"93",	--3046
		x"24",	--3047
		x"4a",	--3048
		x"4b",	--3049
		x"f3",	--3050
		x"f0",	--3051
		x"00",	--3052
		x"93",	--3053
		x"20",	--3054
		x"93",	--3055
		x"24",	--3056
		x"43",	--3057
		x"00",	--3058
		x"3f",	--3059
		x"93",	--3060
		x"23",	--3061
		x"42",	--3062
		x"00",	--3063
		x"3f",	--3064
		x"43",	--3065
		x"00",	--3066
		x"3f",	--3067
		x"12",	--3068
		x"4f",	--3069
		x"93",	--3070
		x"28",	--3071
		x"4e",	--3072
		x"93",	--3073
		x"28",	--3074
		x"92",	--3075
		x"24",	--3076
		x"92",	--3077
		x"24",	--3078
		x"93",	--3079
		x"24",	--3080
		x"93",	--3081
		x"24",	--3082
		x"4f",	--3083
		x"00",	--3084
		x"9e",	--3085
		x"00",	--3086
		x"24",	--3087
		x"93",	--3088
		x"20",	--3089
		x"43",	--3090
		x"4e",	--3091
		x"41",	--3092
		x"41",	--3093
		x"93",	--3094
		x"24",	--3095
		x"93",	--3096
		x"00",	--3097
		x"23",	--3098
		x"43",	--3099
		x"4e",	--3100
		x"41",	--3101
		x"41",	--3102
		x"93",	--3103
		x"00",	--3104
		x"27",	--3105
		x"43",	--3106
		x"3f",	--3107
		x"4f",	--3108
		x"00",	--3109
		x"4e",	--3110
		x"00",	--3111
		x"9b",	--3112
		x"3b",	--3113
		x"9c",	--3114
		x"38",	--3115
		x"4f",	--3116
		x"00",	--3117
		x"4f",	--3118
		x"00",	--3119
		x"4e",	--3120
		x"00",	--3121
		x"4e",	--3122
		x"00",	--3123
		x"9f",	--3124
		x"2b",	--3125
		x"9e",	--3126
		x"28",	--3127
		x"9b",	--3128
		x"2b",	--3129
		x"9e",	--3130
		x"28",	--3131
		x"9f",	--3132
		x"28",	--3133
		x"9c",	--3134
		x"28",	--3135
		x"43",	--3136
		x"3f",	--3137
		x"93",	--3138
		x"23",	--3139
		x"43",	--3140
		x"3f",	--3141
		x"92",	--3142
		x"23",	--3143
		x"4e",	--3144
		x"00",	--3145
		x"4f",	--3146
		x"00",	--3147
		x"8f",	--3148
		x"3f",	--3149
		x"43",	--3150
		x"93",	--3151
		x"34",	--3152
		x"40",	--3153
		x"00",	--3154
		x"e3",	--3155
		x"53",	--3156
		x"93",	--3157
		x"34",	--3158
		x"e3",	--3159
		x"e3",	--3160
		x"53",	--3161
		x"12",	--3162
		x"12",	--3163
		x"f9",	--3164
		x"41",	--3165
		x"b3",	--3166
		x"24",	--3167
		x"e3",	--3168
		x"53",	--3169
		x"b3",	--3170
		x"24",	--3171
		x"e3",	--3172
		x"53",	--3173
		x"41",	--3174
		x"12",	--3175
		x"f8",	--3176
		x"4e",	--3177
		x"41",	--3178
		x"12",	--3179
		x"43",	--3180
		x"93",	--3181
		x"34",	--3182
		x"40",	--3183
		x"00",	--3184
		x"e3",	--3185
		x"e3",	--3186
		x"53",	--3187
		x"63",	--3188
		x"93",	--3189
		x"34",	--3190
		x"e3",	--3191
		x"e3",	--3192
		x"e3",	--3193
		x"53",	--3194
		x"63",	--3195
		x"12",	--3196
		x"f9",	--3197
		x"b3",	--3198
		x"24",	--3199
		x"e3",	--3200
		x"e3",	--3201
		x"53",	--3202
		x"63",	--3203
		x"b3",	--3204
		x"24",	--3205
		x"e3",	--3206
		x"e3",	--3207
		x"53",	--3208
		x"63",	--3209
		x"41",	--3210
		x"41",	--3211
		x"12",	--3212
		x"f8",	--3213
		x"4c",	--3214
		x"4d",	--3215
		x"41",	--3216
		x"40",	--3217
		x"00",	--3218
		x"4e",	--3219
		x"43",	--3220
		x"5f",	--3221
		x"6e",	--3222
		x"9d",	--3223
		x"28",	--3224
		x"8d",	--3225
		x"d3",	--3226
		x"83",	--3227
		x"23",	--3228
		x"41",	--3229
		x"12",	--3230
		x"f9",	--3231
		x"4e",	--3232
		x"41",	--3233
		x"12",	--3234
		x"12",	--3235
		x"12",	--3236
		x"40",	--3237
		x"00",	--3238
		x"4c",	--3239
		x"4d",	--3240
		x"43",	--3241
		x"43",	--3242
		x"5e",	--3243
		x"6f",	--3244
		x"6c",	--3245
		x"6d",	--3246
		x"9b",	--3247
		x"28",	--3248
		x"20",	--3249
		x"9a",	--3250
		x"28",	--3251
		x"8a",	--3252
		x"7b",	--3253
		x"d3",	--3254
		x"83",	--3255
		x"23",	--3256
		x"41",	--3257
		x"41",	--3258
		x"41",	--3259
		x"41",	--3260
		x"12",	--3261
		x"f9",	--3262
		x"4c",	--3263
		x"4d",	--3264
		x"41",	--3265
		x"13",	--3266
		x"d0",	--3267
		x"00",	--3268
		x"3f",	--3269
		x"61",	--3270
		x"74",	--3271
		x"6e",	--3272
		x"20",	--3273
		x"6f",	--3274
		x"20",	--3275
		x"20",	--3276
		x"65",	--3277
		x"20",	--3278
		x"62",	--3279
		x"6e",	--3280
		x"66",	--3281
		x"6c",	--3282
		x"0d",	--3283
		x"00",	--3284
		x"65",	--3285
		x"73",	--3286
		x"6f",	--3287
		x"6c",	--3288
		x"20",	--3289
		x"6f",	--3290
		x"20",	--3291
		x"65",	--3292
		x"20",	--3293
		x"68",	--3294
		x"74",	--3295
		x"0a",	--3296
		x"65",	--3297
		x"72",	--3298
		x"72",	--3299
		x"20",	--3300
		x"69",	--3301
		x"73",	--3302
		x"6e",	--3303
		x"20",	--3304
		x"72",	--3305
		x"75",	--3306
		x"65",	--3307
		x"74",	--3308
		x"0a",	--3309
		x"63",	--3310
		x"72",	--3311
		x"65",	--3312
		x"74",	--3313
		x"75",	--3314
		x"61",	--3315
		x"65",	--3316
		x"0d",	--3317
		x"00",	--3318
		x"25",	--3319
		x"20",	--3320
		x"45",	--3321
		x"54",	--3322
		x"52",	--3323
		x"47",	--3324
		x"54",	--3325
		x"0a",	--3326
		x"25",	--3327
		x"20",	--3328
		x"64",	--3329
		x"0a",	--3330
		x"25",	--3331
		x"20",	--3332
		x"77",	--3333
		x"25",	--3334
		x"20",	--3335
		x"77",	--3336
		x"0a",	--3337
		x"00",	--3338
		x"e3",	--3339
		x"e3",	--3340
		x"e3",	--3341
		x"e3",	--3342
		x"e3",	--3343
		x"e3",	--3344
		x"e3",	--3345
		x"e3",	--3346
		x"0a",	--3347
		x"3d",	--3348
		x"3d",	--3349
		x"3d",	--3350
		x"4d",	--3351
		x"72",	--3352
		x"65",	--3353
		x"20",	--3354
		x"43",	--3355
		x"20",	--3356
		x"3d",	--3357
		x"3d",	--3358
		x"3d",	--3359
		x"0a",	--3360
		x"77",	--3361
		x"69",	--3362
		x"65",	--3363
		x"72",	--3364
		x"61",	--3365
		x"00",	--3366
		x"77",	--3367
		x"00",	--3368
		x"6e",	--3369
		x"6f",	--3370
		x"65",	--3371
		x"00",	--3372
		x"6f",	--3373
		x"74",	--3374
		x"6f",	--3375
		x"64",	--3376
		x"72",	--3377
		x"0d",	--3378
		x"00",	--3379
		x"20",	--3380
		x"00",	--3381
		x"63",	--3382
		x"00",	--3383
		x"72",	--3384
		x"74",	--3385
		x"0a",	--3386
		x"00",	--3387
		x"72",	--3388
		x"6f",	--3389
		x"3a",	--3390
		x"6d",	--3391
		x"73",	--3392
		x"69",	--3393
		x"67",	--3394
		x"61",	--3395
		x"67",	--3396
		x"6d",	--3397
		x"6e",	--3398
		x"0d",	--3399
		x"00",	--3400
		x"6f",	--3401
		x"72",	--3402
		x"63",	--3403
		x"20",	--3404
		x"73",	--3405
		x"67",	--3406
		x"3a",	--3407
		x"0a",	--3408
		x"09",	--3409
		x"73",	--3410
		x"52",	--3411
		x"47",	--3412
		x"53",	--3413
		x"45",	--3414
		x"20",	--3415
		x"41",	--3416
		x"55",	--3417
		x"0d",	--3418
		x"00",	--3419
		x"3d",	--3420
		x"64",	--3421
		x"76",	--3422
		x"25",	--3423
		x"0d",	--3424
		x"00",	--3425
		x"25",	--3426
		x"20",	--3427
		x"45",	--3428
		x"49",	--3429
		x"54",	--3430
		x"52",	--3431
		x"0a",	--3432
		x"72",	--3433
		x"61",	--3434
		x"0a",	--3435
		x"00",	--3436
		x"63",	--3437
		x"69",	--3438
		x"20",	--3439
		x"6f",	--3440
		x"20",	--3441
		x"20",	--3442
		x"75",	--3443
		x"62",	--3444
		x"72",	--3445
		x"0a",	--3446
		x"25",	--3447
		x"20",	--3448
		x"73",	--3449
		x"0a",	--3450
		x"25",	--3451
		x"3a",	--3452
		x"6e",	--3453
		x"20",	--3454
		x"75",	--3455
		x"68",	--3456
		x"63",	--3457
		x"6d",	--3458
		x"61",	--3459
		x"64",	--3460
		x"0a",	--3461
		x"00",	--3462
		x"eb",	--3463
		x"ea",	--3464
		x"ea",	--3465
		x"ea",	--3466
		x"ea",	--3467
		x"ea",	--3468
		x"ea",	--3469
		x"ea",	--3470
		x"ea",	--3471
		x"ea",	--3472
		x"ea",	--3473
		x"ea",	--3474
		x"ea",	--3475
		x"ea",	--3476
		x"ea",	--3477
		x"ea",	--3478
		x"ea",	--3479
		x"ea",	--3480
		x"ea",	--3481
		x"ea",	--3482
		x"ea",	--3483
		x"ea",	--3484
		x"ea",	--3485
		x"ea",	--3486
		x"ea",	--3487
		x"ea",	--3488
		x"ea",	--3489
		x"ea",	--3490
		x"ea",	--3491
		x"eb",	--3492
		x"ea",	--3493
		x"ea",	--3494
		x"ea",	--3495
		x"ea",	--3496
		x"ea",	--3497
		x"ea",	--3498
		x"ea",	--3499
		x"ea",	--3500
		x"ea",	--3501
		x"ea",	--3502
		x"ea",	--3503
		x"ea",	--3504
		x"ea",	--3505
		x"ea",	--3506
		x"ea",	--3507
		x"ea",	--3508
		x"ea",	--3509
		x"ea",	--3510
		x"ea",	--3511
		x"ea",	--3512
		x"ea",	--3513
		x"ea",	--3514
		x"ea",	--3515
		x"ea",	--3516
		x"ea",	--3517
		x"ea",	--3518
		x"ea",	--3519
		x"ea",	--3520
		x"ea",	--3521
		x"ea",	--3522
		x"ea",	--3523
		x"eb",	--3524
		x"eb",	--3525
		x"ea",	--3526
		x"ea",	--3527
		x"ea",	--3528
		x"ea",	--3529
		x"ea",	--3530
		x"ea",	--3531
		x"ea",	--3532
		x"ea",	--3533
		x"ea",	--3534
		x"ea",	--3535
		x"ea",	--3536
		x"ea",	--3537
		x"ea",	--3538
		x"ea",	--3539
		x"ea",	--3540
		x"ea",	--3541
		x"ea",	--3542
		x"ea",	--3543
		x"ea",	--3544
		x"ea",	--3545
		x"ea",	--3546
		x"31",	--3547
		x"33",	--3548
		x"35",	--3549
		x"37",	--3550
		x"39",	--3551
		x"62",	--3552
		x"64",	--3553
		x"66",	--3554
		x"00",	--3555
		x"00",	--3556
		x"00",	--3557
		x"00",	--3558
		x"00",	--3559
		x"01",	--3560
		x"02",	--3561
		x"03",	--3562
		x"03",	--3563
		x"04",	--3564
		x"04",	--3565
		x"04",	--3566
		x"04",	--3567
		x"05",	--3568
		x"05",	--3569
		x"05",	--3570
		x"05",	--3571
		x"05",	--3572
		x"05",	--3573
		x"05",	--3574
		x"05",	--3575
		x"06",	--3576
		x"06",	--3577
		x"06",	--3578
		x"06",	--3579
		x"06",	--3580
		x"06",	--3581
		x"06",	--3582
		x"06",	--3583
		x"06",	--3584
		x"06",	--3585
		x"06",	--3586
		x"06",	--3587
		x"06",	--3588
		x"06",	--3589
		x"06",	--3590
		x"06",	--3591
		x"07",	--3592
		x"07",	--3593
		x"07",	--3594
		x"07",	--3595
		x"07",	--3596
		x"07",	--3597
		x"07",	--3598
		x"07",	--3599
		x"07",	--3600
		x"07",	--3601
		x"07",	--3602
		x"07",	--3603
		x"07",	--3604
		x"07",	--3605
		x"07",	--3606
		x"07",	--3607
		x"07",	--3608
		x"07",	--3609
		x"07",	--3610
		x"07",	--3611
		x"07",	--3612
		x"07",	--3613
		x"07",	--3614
		x"07",	--3615
		x"07",	--3616
		x"07",	--3617
		x"07",	--3618
		x"07",	--3619
		x"07",	--3620
		x"07",	--3621
		x"07",	--3622
		x"07",	--3623
		x"08",	--3624
		x"08",	--3625
		x"08",	--3626
		x"08",	--3627
		x"08",	--3628
		x"08",	--3629
		x"08",	--3630
		x"08",	--3631
		x"08",	--3632
		x"08",	--3633
		x"08",	--3634
		x"08",	--3635
		x"08",	--3636
		x"08",	--3637
		x"08",	--3638
		x"08",	--3639
		x"08",	--3640
		x"08",	--3641
		x"08",	--3642
		x"08",	--3643
		x"08",	--3644
		x"08",	--3645
		x"08",	--3646
		x"08",	--3647
		x"08",	--3648
		x"08",	--3649
		x"08",	--3650
		x"08",	--3651
		x"08",	--3652
		x"08",	--3653
		x"08",	--3654
		x"08",	--3655
		x"08",	--3656
		x"08",	--3657
		x"08",	--3658
		x"08",	--3659
		x"08",	--3660
		x"08",	--3661
		x"08",	--3662
		x"08",	--3663
		x"08",	--3664
		x"08",	--3665
		x"08",	--3666
		x"08",	--3667
		x"08",	--3668
		x"08",	--3669
		x"08",	--3670
		x"08",	--3671
		x"08",	--3672
		x"08",	--3673
		x"08",	--3674
		x"08",	--3675
		x"08",	--3676
		x"08",	--3677
		x"08",	--3678
		x"08",	--3679
		x"08",	--3680
		x"08",	--3681
		x"08",	--3682
		x"08",	--3683
		x"08",	--3684
		x"08",	--3685
		x"08",	--3686
		x"08",	--3687
		x"ff",	--3688
		x"65",	--3689
		x"70",	--3690
		x"00",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"eb",	--4087
		x"e7",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
