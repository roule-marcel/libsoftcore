library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"2e",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"0e",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"2e",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"86",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"20",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"2e",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"0e",	--29
		x"f9",	--30
		x"31",	--31
		x"64",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"30",	--44
		x"b0",	--45
		x"b2",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"7c",	--50
		x"b0",	--51
		x"f4",	--52
		x"21",	--53
		x"3d",	--54
		x"99",	--55
		x"3e",	--56
		x"24",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"e2",	--61
		x"3d",	--62
		x"aa",	--63
		x"3e",	--64
		x"62",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"e2",	--69
		x"3d",	--70
		x"b0",	--71
		x"3e",	--72
		x"d6",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"e2",	--77
		x"3d",	--78
		x"b5",	--79
		x"3e",	--80
		x"52",	--81
		x"7f",	--82
		x"61",	--83
		x"b0",	--84
		x"e2",	--85
		x"3d",	--86
		x"bc",	--87
		x"3e",	--88
		x"da",	--89
		x"7f",	--90
		x"70",	--91
		x"b0",	--92
		x"e2",	--93
		x"3d",	--94
		x"c0",	--95
		x"3e",	--96
		x"1a",	--97
		x"7f",	--98
		x"65",	--99
		x"b0",	--100
		x"e2",	--101
		x"3d",	--102
		x"c8",	--103
		x"3e",	--104
		x"f8",	--105
		x"7f",	--106
		x"73",	--107
		x"b0",	--108
		x"e2",	--109
		x"3d",	--110
		x"d9",	--111
		x"3e",	--112
		x"20",	--113
		x"7f",	--114
		x"63",	--115
		x"b0",	--116
		x"e2",	--117
		x"3d",	--118
		x"ed",	--119
		x"3e",	--120
		x"2e",	--121
		x"7f",	--122
		x"62",	--123
		x"b0",	--124
		x"e2",	--125
		x"0e",	--126
		x"0f",	--127
		x"b0",	--128
		x"78",	--129
		x"2c",	--130
		x"3d",	--131
		x"20",	--132
		x"3e",	--133
		x"80",	--134
		x"0f",	--135
		x"3f",	--136
		x"10",	--137
		x"b0",	--138
		x"80",	--139
		x"0f",	--140
		x"3f",	--141
		x"10",	--142
		x"b0",	--143
		x"c8",	--144
		x"2c",	--145
		x"3d",	--146
		x"20",	--147
		x"3e",	--148
		x"88",	--149
		x"0f",	--150
		x"3f",	--151
		x"06",	--152
		x"b0",	--153
		x"80",	--154
		x"0f",	--155
		x"3f",	--156
		x"06",	--157
		x"b0",	--158
		x"c8",	--159
		x"0e",	--160
		x"3e",	--161
		x"06",	--162
		x"0f",	--163
		x"3f",	--164
		x"10",	--165
		x"b0",	--166
		x"d0",	--167
		x"3e",	--168
		x"98",	--169
		x"0f",	--170
		x"2f",	--171
		x"b0",	--172
		x"d6",	--173
		x"3e",	--174
		x"9c",	--175
		x"0f",	--176
		x"2f",	--177
		x"b0",	--178
		x"d6",	--179
		x"0e",	--180
		x"2e",	--181
		x"0f",	--182
		x"2f",	--183
		x"b0",	--184
		x"06",	--185
		x"0e",	--186
		x"3e",	--187
		x"06",	--188
		x"0f",	--189
		x"3f",	--190
		x"10",	--191
		x"b0",	--192
		x"10",	--193
		x"b0",	--194
		x"ae",	--195
		x"3e",	--196
		x"a0",	--197
		x"0f",	--198
		x"b0",	--199
		x"ee",	--200
		x"0f",	--201
		x"b0",	--202
		x"4c",	--203
		x"3d",	--204
		x"64",	--205
		x"3e",	--206
		x"2a",	--207
		x"0f",	--208
		x"b0",	--209
		x"02",	--210
		x"30",	--211
		x"a0",	--212
		x"03",	--213
		x"03",	--214
		x"03",	--215
		x"30",	--216
		x"d1",	--217
		x"30",	--218
		x"17",	--219
		x"30",	--220
		x"1d",	--221
		x"30",	--222
		x"52",	--223
		x"3c",	--224
		x"32",	--225
		x"0d",	--226
		x"3d",	--227
		x"14",	--228
		x"0e",	--229
		x"3e",	--230
		x"20",	--231
		x"0f",	--232
		x"3f",	--233
		x"7e",	--234
		x"b0",	--235
		x"e8",	--236
		x"31",	--237
		x"10",	--238
		x"30",	--239
		x"a0",	--240
		x"03",	--241
		x"03",	--242
		x"03",	--243
		x"30",	--244
		x"d1",	--245
		x"30",	--246
		x"17",	--247
		x"30",	--248
		x"1d",	--249
		x"30",	--250
		x"52",	--251
		x"3c",	--252
		x"32",	--253
		x"0d",	--254
		x"3d",	--255
		x"12",	--256
		x"0e",	--257
		x"3e",	--258
		x"16",	--259
		x"0f",	--260
		x"3f",	--261
		x"52",	--262
		x"b0",	--263
		x"e8",	--264
		x"31",	--265
		x"10",	--266
		x"0e",	--267
		x"3e",	--268
		x"42",	--269
		x"0f",	--270
		x"3f",	--271
		x"6e",	--272
		x"b0",	--273
		x"ee",	--274
		x"b0",	--275
		x"c6",	--276
		x"f2",	--277
		x"80",	--278
		x"19",	--279
		x"32",	--280
		x"0b",	--281
		x"0a",	--282
		x"05",	--283
		x"1b",	--284
		x"03",	--285
		x"2b",	--286
		x"01",	--287
		x"0b",	--288
		x"b0",	--289
		x"4e",	--290
		x"0f",	--291
		x"fc",	--292
		x"b0",	--293
		x"76",	--294
		x"0b",	--295
		x"3e",	--296
		x"7f",	--297
		x"0d",	--298
		x"06",	--299
		x"7f",	--300
		x"1b",	--301
		x"ed",	--302
		x"7f",	--303
		x"1c",	--304
		x"12",	--305
		x"30",	--306
		x"f8",	--307
		x"b0",	--308
		x"f4",	--309
		x"21",	--310
		x"3f",	--311
		x"1a",	--312
		x"0f",	--313
		x"0a",	--314
		x"ca",	--315
		x"00",	--316
		x"0e",	--317
		x"5f",	--318
		x"1a",	--319
		x"b0",	--320
		x"16",	--321
		x"0a",	--322
		x"dd",	--323
		x"0a",	--324
		x"db",	--325
		x"3a",	--326
		x"30",	--327
		x"fb",	--328
		x"b0",	--329
		x"f4",	--330
		x"21",	--331
		x"d4",	--332
		x"3a",	--333
		x"28",	--334
		x"d1",	--335
		x"82",	--336
		x"10",	--337
		x"0c",	--338
		x"4e",	--339
		x"8e",	--340
		x"0e",	--341
		x"30",	--342
		x"ff",	--343
		x"81",	--344
		x"9e",	--345
		x"b0",	--346
		x"f4",	--347
		x"21",	--348
		x"1f",	--349
		x"9a",	--350
		x"3e",	--351
		x"1a",	--352
		x"0e",	--353
		x"0e",	--354
		x"ce",	--355
		x"00",	--356
		x"1a",	--357
		x"ba",	--358
		x"1b",	--359
		x"04",	--360
		x"7f",	--361
		x"5b",	--362
		x"b5",	--363
		x"b1",	--364
		x"2b",	--365
		x"b2",	--366
		x"7f",	--367
		x"42",	--368
		x"17",	--369
		x"7f",	--370
		x"43",	--371
		x"04",	--372
		x"7f",	--373
		x"41",	--374
		x"a8",	--375
		x"07",	--376
		x"7f",	--377
		x"43",	--378
		x"16",	--379
		x"7f",	--380
		x"44",	--381
		x"a1",	--382
		x"1b",	--383
		x"30",	--384
		x"02",	--385
		x"b0",	--386
		x"f4",	--387
		x"21",	--388
		x"b0",	--389
		x"80",	--390
		x"0b",	--391
		x"98",	--392
		x"30",	--393
		x"07",	--394
		x"b0",	--395
		x"f4",	--396
		x"21",	--397
		x"b0",	--398
		x"a8",	--399
		x"0b",	--400
		x"8f",	--401
		x"30",	--402
		x"0e",	--403
		x"b0",	--404
		x"f4",	--405
		x"21",	--406
		x"b0",	--407
		x"d0",	--408
		x"0b",	--409
		x"86",	--410
		x"30",	--411
		x"16",	--412
		x"b0",	--413
		x"f4",	--414
		x"21",	--415
		x"b0",	--416
		x"f8",	--417
		x"0b",	--418
		x"7d",	--419
		x"30",	--420
		x"72",	--421
		x"82",	--422
		x"20",	--423
		x"30",	--424
		x"0b",	--425
		x"0a",	--426
		x"21",	--427
		x"0a",	--428
		x"0b",	--429
		x"2f",	--430
		x"1b",	--431
		x"0e",	--432
		x"1f",	--433
		x"02",	--434
		x"b0",	--435
		x"32",	--436
		x"0d",	--437
		x"2a",	--438
		x"18",	--439
		x"0e",	--440
		x"1f",	--441
		x"04",	--442
		x"81",	--443
		x"02",	--444
		x"b0",	--445
		x"32",	--446
		x"0e",	--447
		x"1d",	--448
		x"02",	--449
		x"1f",	--450
		x"20",	--451
		x"b0",	--452
		x"02",	--453
		x"0f",	--454
		x"21",	--455
		x"3a",	--456
		x"3b",	--457
		x"30",	--458
		x"3d",	--459
		x"64",	--460
		x"3e",	--461
		x"2a",	--462
		x"f2",	--463
		x"3e",	--464
		x"2a",	--465
		x"ef",	--466
		x"0e",	--467
		x"1f",	--468
		x"24",	--469
		x"b0",	--470
		x"7c",	--471
		x"0e",	--472
		x"1f",	--473
		x"22",	--474
		x"b0",	--475
		x"7c",	--476
		x"30",	--477
		x"7a",	--478
		x"b0",	--479
		x"f4",	--480
		x"21",	--481
		x"30",	--482
		x"b2",	--483
		x"00",	--484
		x"09",	--485
		x"1f",	--486
		x"24",	--487
		x"b0",	--488
		x"38",	--489
		x"1f",	--490
		x"22",	--491
		x"b0",	--492
		x"38",	--493
		x"30",	--494
		x"0e",	--495
		x"3f",	--496
		x"a6",	--497
		x"b0",	--498
		x"be",	--499
		x"82",	--500
		x"00",	--501
		x"ef",	--502
		x"82",	--503
		x"24",	--504
		x"82",	--505
		x"22",	--506
		x"30",	--507
		x"0b",	--508
		x"0a",	--509
		x"21",	--510
		x"0b",	--511
		x"3f",	--512
		x"03",	--513
		x"30",	--514
		x"23",	--515
		x"0e",	--516
		x"1f",	--517
		x"02",	--518
		x"b0",	--519
		x"00",	--520
		x"0a",	--521
		x"0e",	--522
		x"1f",	--523
		x"04",	--524
		x"b0",	--525
		x"00",	--526
		x"0b",	--527
		x"0f",	--528
		x"0a",	--529
		x"30",	--530
		x"ad",	--531
		x"b0",	--532
		x"f4",	--533
		x"31",	--534
		x"06",	--535
		x"0e",	--536
		x"1f",	--537
		x"24",	--538
		x"b0",	--539
		x"7c",	--540
		x"0e",	--541
		x"1f",	--542
		x"22",	--543
		x"b0",	--544
		x"7c",	--545
		x"0f",	--546
		x"21",	--547
		x"3a",	--548
		x"3b",	--549
		x"30",	--550
		x"0e",	--551
		x"1f",	--552
		x"06",	--553
		x"b0",	--554
		x"32",	--555
		x"1d",	--556
		x"0e",	--557
		x"1f",	--558
		x"00",	--559
		x"b0",	--560
		x"02",	--561
		x"d1",	--562
		x"30",	--563
		x"81",	--564
		x"b0",	--565
		x"f4",	--566
		x"a1",	--567
		x"00",	--568
		x"30",	--569
		x"92",	--570
		x"b0",	--571
		x"f4",	--572
		x"21",	--573
		x"3f",	--574
		x"e3",	--575
		x"3e",	--576
		x"9c",	--577
		x"1f",	--578
		x"24",	--579
		x"b0",	--580
		x"7c",	--581
		x"3e",	--582
		x"64",	--583
		x"1f",	--584
		x"22",	--585
		x"b0",	--586
		x"7c",	--587
		x"1d",	--588
		x"3e",	--589
		x"c8",	--590
		x"1f",	--591
		x"00",	--592
		x"b0",	--593
		x"02",	--594
		x"30",	--595
		x"3e",	--596
		x"64",	--597
		x"1f",	--598
		x"24",	--599
		x"b0",	--600
		x"7c",	--601
		x"3e",	--602
		x"9c",	--603
		x"1f",	--604
		x"22",	--605
		x"b0",	--606
		x"7c",	--607
		x"1d",	--608
		x"3e",	--609
		x"c8",	--610
		x"1f",	--611
		x"00",	--612
		x"b0",	--613
		x"02",	--614
		x"30",	--615
		x"3e",	--616
		x"c4",	--617
		x"1f",	--618
		x"24",	--619
		x"b0",	--620
		x"7c",	--621
		x"3e",	--622
		x"c4",	--623
		x"1f",	--624
		x"22",	--625
		x"b0",	--626
		x"7c",	--627
		x"1d",	--628
		x"3e",	--629
		x"c8",	--630
		x"1f",	--631
		x"00",	--632
		x"b0",	--633
		x"02",	--634
		x"30",	--635
		x"3e",	--636
		x"3c",	--637
		x"1f",	--638
		x"24",	--639
		x"b0",	--640
		x"7c",	--641
		x"3e",	--642
		x"3c",	--643
		x"1f",	--644
		x"22",	--645
		x"b0",	--646
		x"7c",	--647
		x"1d",	--648
		x"3e",	--649
		x"c8",	--650
		x"1f",	--651
		x"00",	--652
		x"b0",	--653
		x"02",	--654
		x"30",	--655
		x"30",	--656
		x"b5",	--657
		x"b0",	--658
		x"f4",	--659
		x"21",	--660
		x"0f",	--661
		x"30",	--662
		x"b2",	--663
		x"00",	--664
		x"92",	--665
		x"b2",	--666
		x"30",	--667
		x"94",	--668
		x"b2",	--669
		x"41",	--670
		x"96",	--671
		x"30",	--672
		x"cb",	--673
		x"b0",	--674
		x"f4",	--675
		x"92",	--676
		x"90",	--677
		x"b1",	--678
		x"e9",	--679
		x"00",	--680
		x"b0",	--681
		x"f4",	--682
		x"21",	--683
		x"0f",	--684
		x"30",	--685
		x"0b",	--686
		x"0a",	--687
		x"09",	--688
		x"09",	--689
		x"1f",	--690
		x"22",	--691
		x"b0",	--692
		x"de",	--693
		x"0a",	--694
		x"0b",	--695
		x"1e",	--696
		x"24",	--697
		x"1f",	--698
		x"26",	--699
		x"b0",	--700
		x"78",	--701
		x"89",	--702
		x"24",	--703
		x"89",	--704
		x"26",	--705
		x"0d",	--706
		x"0e",	--707
		x"0f",	--708
		x"b0",	--709
		x"44",	--710
		x"0c",	--711
		x"3d",	--712
		x"00",	--713
		x"b0",	--714
		x"78",	--715
		x"0a",	--716
		x"0b",	--717
		x"3c",	--718
		x"66",	--719
		x"3d",	--720
		x"66",	--721
		x"b0",	--722
		x"88",	--723
		x"0f",	--724
		x"01",	--725
		x"18",	--726
		x"3c",	--727
		x"cd",	--728
		x"3d",	--729
		x"cc",	--730
		x"0e",	--731
		x"0f",	--732
		x"b0",	--733
		x"28",	--734
		x"0f",	--735
		x"04",	--736
		x"3a",	--737
		x"cd",	--738
		x"3b",	--739
		x"cc",	--740
		x"0d",	--741
		x"0e",	--742
		x"1f",	--743
		x"20",	--744
		x"b0",	--745
		x"1c",	--746
		x"39",	--747
		x"3a",	--748
		x"3b",	--749
		x"30",	--750
		x"3a",	--751
		x"66",	--752
		x"3b",	--753
		x"66",	--754
		x"f1",	--755
		x"0b",	--756
		x"0a",	--757
		x"0b",	--758
		x"0a",	--759
		x"8f",	--760
		x"20",	--761
		x"8f",	--762
		x"22",	--763
		x"11",	--764
		x"16",	--765
		x"11",	--766
		x"16",	--767
		x"11",	--768
		x"16",	--769
		x"11",	--770
		x"16",	--771
		x"11",	--772
		x"16",	--773
		x"11",	--774
		x"16",	--775
		x"1d",	--776
		x"12",	--777
		x"1e",	--778
		x"14",	--779
		x"b0",	--780
		x"aa",	--781
		x"31",	--782
		x"0c",	--783
		x"8b",	--784
		x"28",	--785
		x"0e",	--786
		x"3f",	--787
		x"5c",	--788
		x"b0",	--789
		x"be",	--790
		x"8b",	--791
		x"2a",	--792
		x"3a",	--793
		x"3b",	--794
		x"30",	--795
		x"0b",	--796
		x"0b",	--797
		x"1f",	--798
		x"22",	--799
		x"b0",	--800
		x"de",	--801
		x"8b",	--802
		x"24",	--803
		x"8b",	--804
		x"26",	--805
		x"0d",	--806
		x"1e",	--807
		x"28",	--808
		x"1f",	--809
		x"2a",	--810
		x"b0",	--811
		x"02",	--812
		x"3b",	--813
		x"30",	--814
		x"0b",	--815
		x"0b",	--816
		x"0d",	--817
		x"3e",	--818
		x"00",	--819
		x"1f",	--820
		x"20",	--821
		x"b0",	--822
		x"1c",	--823
		x"1f",	--824
		x"2a",	--825
		x"b0",	--826
		x"2a",	--827
		x"3b",	--828
		x"30",	--829
		x"0b",	--830
		x"0b",	--831
		x"0d",	--832
		x"8d",	--833
		x"8d",	--834
		x"8d",	--835
		x"8d",	--836
		x"0f",	--837
		x"b0",	--838
		x"78",	--839
		x"0d",	--840
		x"0e",	--841
		x"0f",	--842
		x"b0",	--843
		x"30",	--844
		x"3b",	--845
		x"30",	--846
		x"0b",	--847
		x"0a",	--848
		x"0a",	--849
		x"3b",	--850
		x"00",	--851
		x"0d",	--852
		x"0e",	--853
		x"1f",	--854
		x"68",	--855
		x"b0",	--856
		x"1c",	--857
		x"0d",	--858
		x"0e",	--859
		x"1f",	--860
		x"66",	--861
		x"b0",	--862
		x"1c",	--863
		x"30",	--864
		x"02",	--865
		x"b0",	--866
		x"f4",	--867
		x"21",	--868
		x"3a",	--869
		x"3b",	--870
		x"30",	--871
		x"82",	--872
		x"68",	--873
		x"82",	--874
		x"66",	--875
		x"30",	--876
		x"0b",	--877
		x"0a",	--878
		x"21",	--879
		x"0a",	--880
		x"0b",	--881
		x"b2",	--882
		x"02",	--883
		x"4e",	--884
		x"3a",	--885
		x"03",	--886
		x"53",	--887
		x"3e",	--888
		x"0e",	--889
		x"1f",	--890
		x"02",	--891
		x"b0",	--892
		x"32",	--893
		x"0a",	--894
		x"0e",	--895
		x"1f",	--896
		x"04",	--897
		x"b0",	--898
		x"32",	--899
		x"0b",	--900
		x"0f",	--901
		x"0a",	--902
		x"30",	--903
		x"4f",	--904
		x"b0",	--905
		x"f4",	--906
		x"31",	--907
		x"06",	--908
		x"0e",	--909
		x"0f",	--910
		x"b0",	--911
		x"ae",	--912
		x"0c",	--913
		x"3d",	--914
		x"c8",	--915
		x"b0",	--916
		x"38",	--917
		x"0c",	--918
		x"0d",	--919
		x"0e",	--920
		x"3f",	--921
		x"80",	--922
		x"b0",	--923
		x"c4",	--924
		x"0d",	--925
		x"0e",	--926
		x"1f",	--927
		x"68",	--928
		x"b0",	--929
		x"1c",	--930
		x"0e",	--931
		x"0f",	--932
		x"b0",	--933
		x"ae",	--934
		x"0c",	--935
		x"3d",	--936
		x"c8",	--937
		x"b0",	--938
		x"38",	--939
		x"0d",	--940
		x"0e",	--941
		x"1f",	--942
		x"66",	--943
		x"b0",	--944
		x"1c",	--945
		x"0f",	--946
		x"21",	--947
		x"3a",	--948
		x"3b",	--949
		x"30",	--950
		x"0e",	--951
		x"1f",	--952
		x"06",	--953
		x"b0",	--954
		x"32",	--955
		x"1d",	--956
		x"0e",	--957
		x"1f",	--958
		x"02",	--959
		x"b0",	--960
		x"02",	--961
		x"b6",	--962
		x"0e",	--963
		x"3f",	--964
		x"9e",	--965
		x"b0",	--966
		x"be",	--967
		x"82",	--968
		x"02",	--969
		x"aa",	--970
		x"30",	--971
		x"09",	--972
		x"b0",	--973
		x"f4",	--974
		x"b1",	--975
		x"23",	--976
		x"00",	--977
		x"b0",	--978
		x"f4",	--979
		x"a1",	--980
		x"00",	--981
		x"30",	--982
		x"34",	--983
		x"b0",	--984
		x"f4",	--985
		x"21",	--986
		x"3f",	--987
		x"d6",	--988
		x"0b",	--989
		x"0a",	--990
		x"1f",	--991
		x"6c",	--992
		x"b0",	--993
		x"de",	--994
		x"0a",	--995
		x"0b",	--996
		x"1f",	--997
		x"6a",	--998
		x"b0",	--999
		x"de",	--1000
		x"0b",	--1001
		x"0a",	--1002
		x"3e",	--1003
		x"3f",	--1004
		x"1e",	--1005
		x"0f",	--1006
		x"0f",	--1007
		x"0e",	--1008
		x"30",	--1009
		x"57",	--1010
		x"30",	--1011
		x"26",	--1012
		x"b0",	--1013
		x"06",	--1014
		x"31",	--1015
		x"0c",	--1016
		x"30",	--1017
		x"26",	--1018
		x"30",	--1019
		x"5f",	--1020
		x"b0",	--1021
		x"f4",	--1022
		x"21",	--1023
		x"3a",	--1024
		x"3b",	--1025
		x"30",	--1026
		x"82",	--1027
		x"6a",	--1028
		x"82",	--1029
		x"6c",	--1030
		x"30",	--1031
		x"82",	--1032
		x"68",	--1033
		x"82",	--1034
		x"66",	--1035
		x"30",	--1036
		x"0b",	--1037
		x"0a",	--1038
		x"09",	--1039
		x"08",	--1040
		x"21",	--1041
		x"0a",	--1042
		x"0b",	--1043
		x"81",	--1044
		x"00",	--1045
		x"1f",	--1046
		x"1c",	--1047
		x"b2",	--1048
		x"04",	--1049
		x"6f",	--1050
		x"92",	--1051
		x"0e",	--1052
		x"0e",	--1053
		x"1f",	--1054
		x"02",	--1055
		x"b0",	--1056
		x"32",	--1057
		x"08",	--1058
		x"3a",	--1059
		x"03",	--1060
		x"1e",	--1061
		x"09",	--1062
		x"0d",	--1063
		x"0e",	--1064
		x"1f",	--1065
		x"04",	--1066
		x"b0",	--1067
		x"02",	--1068
		x"0f",	--1069
		x"21",	--1070
		x"38",	--1071
		x"39",	--1072
		x"3a",	--1073
		x"3b",	--1074
		x"30",	--1075
		x"82",	--1076
		x"0e",	--1077
		x"49",	--1078
		x"82",	--1079
		x"0e",	--1080
		x"1f",	--1081
		x"04",	--1082
		x"b0",	--1083
		x"2a",	--1084
		x"0f",	--1085
		x"21",	--1086
		x"38",	--1087
		x"39",	--1088
		x"3a",	--1089
		x"3b",	--1090
		x"30",	--1091
		x"0e",	--1092
		x"1f",	--1093
		x"04",	--1094
		x"b0",	--1095
		x"32",	--1096
		x"09",	--1097
		x"3a",	--1098
		x"05",	--1099
		x"da",	--1100
		x"0e",	--1101
		x"1f",	--1102
		x"06",	--1103
		x"b0",	--1104
		x"32",	--1105
		x"0a",	--1106
		x"0e",	--1107
		x"1f",	--1108
		x"08",	--1109
		x"b0",	--1110
		x"32",	--1111
		x"0b",	--1112
		x"0f",	--1113
		x"0a",	--1114
		x"30",	--1115
		x"64",	--1116
		x"b0",	--1117
		x"f4",	--1118
		x"31",	--1119
		x"06",	--1120
		x"0e",	--1121
		x"0f",	--1122
		x"b0",	--1123
		x"ae",	--1124
		x"0c",	--1125
		x"3d",	--1126
		x"c8",	--1127
		x"b0",	--1128
		x"38",	--1129
		x"0d",	--1130
		x"0e",	--1131
		x"1f",	--1132
		x"68",	--1133
		x"b0",	--1134
		x"1c",	--1135
		x"0e",	--1136
		x"0f",	--1137
		x"b0",	--1138
		x"ae",	--1139
		x"0c",	--1140
		x"3d",	--1141
		x"c8",	--1142
		x"b0",	--1143
		x"38",	--1144
		x"0d",	--1145
		x"0e",	--1146
		x"1f",	--1147
		x"66",	--1148
		x"b0",	--1149
		x"1c",	--1150
		x"a7",	--1151
		x"0f",	--1152
		x"b0",	--1153
		x"ba",	--1154
		x"0f",	--1155
		x"21",	--1156
		x"38",	--1157
		x"39",	--1158
		x"3a",	--1159
		x"3b",	--1160
		x"30",	--1161
		x"0e",	--1162
		x"3f",	--1163
		x"ba",	--1164
		x"b0",	--1165
		x"be",	--1166
		x"82",	--1167
		x"04",	--1168
		x"89",	--1169
		x"1f",	--1170
		x"82",	--1171
		x"10",	--1172
		x"01",	--1173
		x"0f",	--1174
		x"82",	--1175
		x"10",	--1176
		x"0f",	--1177
		x"30",	--1178
		x"5e",	--1179
		x"19",	--1180
		x"4e",	--1181
		x"0f",	--1182
		x"03",	--1183
		x"c2",	--1184
		x"19",	--1185
		x"30",	--1186
		x"c2",	--1187
		x"19",	--1188
		x"30",	--1189
		x"1e",	--1190
		x"12",	--1191
		x"3e",	--1192
		x"06",	--1193
		x"0f",	--1194
		x"0f",	--1195
		x"10",	--1196
		x"6c",	--1197
		x"c2",	--1198
		x"19",	--1199
		x"3e",	--1200
		x"07",	--1201
		x"03",	--1202
		x"82",	--1203
		x"12",	--1204
		x"30",	--1205
		x"1e",	--1206
		x"82",	--1207
		x"12",	--1208
		x"30",	--1209
		x"f2",	--1210
		x"0e",	--1211
		x"19",	--1212
		x"f2",	--1213
		x"f2",	--1214
		x"0a",	--1215
		x"19",	--1216
		x"ee",	--1217
		x"e2",	--1218
		x"19",	--1219
		x"eb",	--1220
		x"f2",	--1221
		x"0d",	--1222
		x"19",	--1223
		x"e7",	--1224
		x"f2",	--1225
		x"09",	--1226
		x"19",	--1227
		x"e3",	--1228
		x"f2",	--1229
		x"03",	--1230
		x"19",	--1231
		x"df",	--1232
		x"f2",	--1233
		x"07",	--1234
		x"19",	--1235
		x"db",	--1236
		x"8f",	--1237
		x"00",	--1238
		x"8f",	--1239
		x"02",	--1240
		x"9f",	--1241
		x"02",	--1242
		x"04",	--1243
		x"9f",	--1244
		x"04",	--1245
		x"06",	--1246
		x"9f",	--1247
		x"06",	--1248
		x"08",	--1249
		x"9f",	--1250
		x"08",	--1251
		x"0a",	--1252
		x"9f",	--1253
		x"0a",	--1254
		x"10",	--1255
		x"9f",	--1256
		x"0c",	--1257
		x"12",	--1258
		x"8f",	--1259
		x"14",	--1260
		x"8f",	--1261
		x"16",	--1262
		x"8f",	--1263
		x"0c",	--1264
		x"8f",	--1265
		x"0e",	--1266
		x"8f",	--1267
		x"18",	--1268
		x"8f",	--1269
		x"1a",	--1270
		x"8f",	--1271
		x"1c",	--1272
		x"8f",	--1273
		x"1e",	--1274
		x"30",	--1275
		x"8f",	--1276
		x"0c",	--1277
		x"8f",	--1278
		x"0e",	--1279
		x"8f",	--1280
		x"18",	--1281
		x"8f",	--1282
		x"1a",	--1283
		x"8f",	--1284
		x"1c",	--1285
		x"8f",	--1286
		x"1e",	--1287
		x"30",	--1288
		x"8f",	--1289
		x"00",	--1290
		x"8f",	--1291
		x"02",	--1292
		x"30",	--1293
		x"8f",	--1294
		x"04",	--1295
		x"8f",	--1296
		x"06",	--1297
		x"30",	--1298
		x"8f",	--1299
		x"08",	--1300
		x"8f",	--1301
		x"0a",	--1302
		x"30",	--1303
		x"8f",	--1304
		x"0c",	--1305
		x"8f",	--1306
		x"0e",	--1307
		x"30",	--1308
		x"8f",	--1309
		x"10",	--1310
		x"8f",	--1311
		x"12",	--1312
		x"30",	--1313
		x"0b",	--1314
		x"0a",	--1315
		x"09",	--1316
		x"07",	--1317
		x"06",	--1318
		x"05",	--1319
		x"04",	--1320
		x"09",	--1321
		x"04",	--1322
		x"05",	--1323
		x"16",	--1324
		x"14",	--1325
		x"17",	--1326
		x"16",	--1327
		x"1a",	--1328
		x"0c",	--1329
		x"1b",	--1330
		x"0e",	--1331
		x"0c",	--1332
		x"0d",	--1333
		x"0e",	--1334
		x"0f",	--1335
		x"b0",	--1336
		x"28",	--1337
		x"1c",	--1338
		x"10",	--1339
		x"1d",	--1340
		x"12",	--1341
		x"0f",	--1342
		x"5b",	--1343
		x"0e",	--1344
		x"0f",	--1345
		x"b0",	--1346
		x"78",	--1347
		x"06",	--1348
		x"07",	--1349
		x"89",	--1350
		x"14",	--1351
		x"89",	--1352
		x"16",	--1353
		x"0c",	--1354
		x"0d",	--1355
		x"0e",	--1356
		x"0f",	--1357
		x"b0",	--1358
		x"28",	--1359
		x"0f",	--1360
		x"5c",	--1361
		x"89",	--1362
		x"14",	--1363
		x"89",	--1364
		x"16",	--1365
		x"0c",	--1366
		x"0d",	--1367
		x"0e",	--1368
		x"0f",	--1369
		x"b0",	--1370
		x"c4",	--1371
		x"0a",	--1372
		x"0b",	--1373
		x"1c",	--1374
		x"18",	--1375
		x"1d",	--1376
		x"1a",	--1377
		x"b0",	--1378
		x"78",	--1379
		x"06",	--1380
		x"07",	--1381
		x"89",	--1382
		x"18",	--1383
		x"89",	--1384
		x"1a",	--1385
		x"2c",	--1386
		x"1d",	--1387
		x"02",	--1388
		x"0e",	--1389
		x"0f",	--1390
		x"b0",	--1391
		x"14",	--1392
		x"04",	--1393
		x"05",	--1394
		x"1c",	--1395
		x"04",	--1396
		x"1d",	--1397
		x"06",	--1398
		x"0e",	--1399
		x"0f",	--1400
		x"b0",	--1401
		x"14",	--1402
		x"0c",	--1403
		x"0d",	--1404
		x"b0",	--1405
		x"78",	--1406
		x"06",	--1407
		x"07",	--1408
		x"1c",	--1409
		x"1c",	--1410
		x"1d",	--1411
		x"1e",	--1412
		x"0e",	--1413
		x"0f",	--1414
		x"b0",	--1415
		x"c4",	--1416
		x"1c",	--1417
		x"08",	--1418
		x"1d",	--1419
		x"0a",	--1420
		x"b0",	--1421
		x"14",	--1422
		x"0c",	--1423
		x"0d",	--1424
		x"b0",	--1425
		x"78",	--1426
		x"34",	--1427
		x"35",	--1428
		x"36",	--1429
		x"37",	--1430
		x"39",	--1431
		x"3a",	--1432
		x"3b",	--1433
		x"30",	--1434
		x"0e",	--1435
		x"0f",	--1436
		x"b0",	--1437
		x"c4",	--1438
		x"06",	--1439
		x"07",	--1440
		x"89",	--1441
		x"14",	--1442
		x"89",	--1443
		x"16",	--1444
		x"0c",	--1445
		x"0d",	--1446
		x"0e",	--1447
		x"0f",	--1448
		x"b0",	--1449
		x"88",	--1450
		x"0f",	--1451
		x"01",	--1452
		x"a4",	--1453
		x"0a",	--1454
		x"0b",	--1455
		x"a5",	--1456
		x"0b",	--1457
		x"0a",	--1458
		x"21",	--1459
		x"0a",	--1460
		x"0b",	--1461
		x"30",	--1462
		x"1e",	--1463
		x"b0",	--1464
		x"f4",	--1465
		x"21",	--1466
		x"3a",	--1467
		x"03",	--1468
		x"1b",	--1469
		x"0e",	--1470
		x"1f",	--1471
		x"02",	--1472
		x"b0",	--1473
		x"32",	--1474
		x"0a",	--1475
		x"0e",	--1476
		x"1f",	--1477
		x"04",	--1478
		x"b0",	--1479
		x"32",	--1480
		x"0b",	--1481
		x"0f",	--1482
		x"0a",	--1483
		x"30",	--1484
		x"66",	--1485
		x"b0",	--1486
		x"f4",	--1487
		x"31",	--1488
		x"06",	--1489
		x"8a",	--1490
		x"00",	--1491
		x"0f",	--1492
		x"21",	--1493
		x"3a",	--1494
		x"3b",	--1495
		x"30",	--1496
		x"30",	--1497
		x"26",	--1498
		x"b0",	--1499
		x"f4",	--1500
		x"b1",	--1501
		x"40",	--1502
		x"00",	--1503
		x"b0",	--1504
		x"f4",	--1505
		x"a1",	--1506
		x"00",	--1507
		x"30",	--1508
		x"51",	--1509
		x"b0",	--1510
		x"f4",	--1511
		x"21",	--1512
		x"3f",	--1513
		x"ea",	--1514
		x"0b",	--1515
		x"21",	--1516
		x"0b",	--1517
		x"1f",	--1518
		x"17",	--1519
		x"16",	--1520
		x"30",	--1521
		x"81",	--1522
		x"b0",	--1523
		x"f4",	--1524
		x"21",	--1525
		x"0e",	--1526
		x"1f",	--1527
		x"02",	--1528
		x"b0",	--1529
		x"32",	--1530
		x"2f",	--1531
		x"0f",	--1532
		x"30",	--1533
		x"66",	--1534
		x"b0",	--1535
		x"f4",	--1536
		x"31",	--1537
		x"06",	--1538
		x"0f",	--1539
		x"21",	--1540
		x"3b",	--1541
		x"30",	--1542
		x"30",	--1543
		x"26",	--1544
		x"b0",	--1545
		x"f4",	--1546
		x"b1",	--1547
		x"40",	--1548
		x"00",	--1549
		x"b0",	--1550
		x"f4",	--1551
		x"a1",	--1552
		x"00",	--1553
		x"30",	--1554
		x"72",	--1555
		x"b0",	--1556
		x"f4",	--1557
		x"21",	--1558
		x"3f",	--1559
		x"eb",	--1560
		x"0b",	--1561
		x"0a",	--1562
		x"8e",	--1563
		x"00",	--1564
		x"6d",	--1565
		x"4d",	--1566
		x"5e",	--1567
		x"1f",	--1568
		x"0a",	--1569
		x"0c",	--1570
		x"0f",	--1571
		x"7b",	--1572
		x"0a",	--1573
		x"2b",	--1574
		x"0c",	--1575
		x"0c",	--1576
		x"0c",	--1577
		x"0c",	--1578
		x"8d",	--1579
		x"0c",	--1580
		x"3c",	--1581
		x"d0",	--1582
		x"1a",	--1583
		x"7d",	--1584
		x"4d",	--1585
		x"17",	--1586
		x"7d",	--1587
		x"78",	--1588
		x"1a",	--1589
		x"4b",	--1590
		x"7b",	--1591
		x"d0",	--1592
		x"0a",	--1593
		x"e9",	--1594
		x"7b",	--1595
		x"0a",	--1596
		x"34",	--1597
		x"0c",	--1598
		x"0b",	--1599
		x"0b",	--1600
		x"0b",	--1601
		x"0c",	--1602
		x"8d",	--1603
		x"0c",	--1604
		x"3c",	--1605
		x"d0",	--1606
		x"7d",	--1607
		x"4d",	--1608
		x"e9",	--1609
		x"9e",	--1610
		x"00",	--1611
		x"0f",	--1612
		x"3a",	--1613
		x"3b",	--1614
		x"30",	--1615
		x"1a",	--1616
		x"de",	--1617
		x"4b",	--1618
		x"7b",	--1619
		x"9f",	--1620
		x"7b",	--1621
		x"06",	--1622
		x"0a",	--1623
		x"0c",	--1624
		x"0c",	--1625
		x"0c",	--1626
		x"0c",	--1627
		x"8d",	--1628
		x"0c",	--1629
		x"3c",	--1630
		x"a9",	--1631
		x"1a",	--1632
		x"ce",	--1633
		x"4b",	--1634
		x"7b",	--1635
		x"bf",	--1636
		x"7b",	--1637
		x"06",	--1638
		x"0a",	--1639
		x"0c",	--1640
		x"0c",	--1641
		x"0c",	--1642
		x"0c",	--1643
		x"8d",	--1644
		x"0c",	--1645
		x"3c",	--1646
		x"c9",	--1647
		x"1a",	--1648
		x"be",	--1649
		x"8d",	--1650
		x"0d",	--1651
		x"30",	--1652
		x"88",	--1653
		x"b0",	--1654
		x"f4",	--1655
		x"21",	--1656
		x"0c",	--1657
		x"0f",	--1658
		x"3a",	--1659
		x"3b",	--1660
		x"30",	--1661
		x"0c",	--1662
		x"ca",	--1663
		x"0b",	--1664
		x"0a",	--1665
		x"8e",	--1666
		x"00",	--1667
		x"6b",	--1668
		x"4b",	--1669
		x"37",	--1670
		x"1f",	--1671
		x"1a",	--1672
		x"0c",	--1673
		x"12",	--1674
		x"4d",	--1675
		x"7d",	--1676
		x"d0",	--1677
		x"7d",	--1678
		x"0a",	--1679
		x"22",	--1680
		x"0c",	--1681
		x"0d",	--1682
		x"0d",	--1683
		x"0d",	--1684
		x"0c",	--1685
		x"8b",	--1686
		x"0c",	--1687
		x"3c",	--1688
		x"d0",	--1689
		x"7b",	--1690
		x"4b",	--1691
		x"07",	--1692
		x"7b",	--1693
		x"2d",	--1694
		x"eb",	--1695
		x"3a",	--1696
		x"7b",	--1697
		x"4b",	--1698
		x"f9",	--1699
		x"02",	--1700
		x"32",	--1701
		x"03",	--1702
		x"82",	--1703
		x"32",	--1704
		x"82",	--1705
		x"38",	--1706
		x"1f",	--1707
		x"3a",	--1708
		x"32",	--1709
		x"9e",	--1710
		x"00",	--1711
		x"3a",	--1712
		x"3b",	--1713
		x"30",	--1714
		x"8b",	--1715
		x"0b",	--1716
		x"30",	--1717
		x"88",	--1718
		x"b0",	--1719
		x"f4",	--1720
		x"21",	--1721
		x"0f",	--1722
		x"3a",	--1723
		x"3b",	--1724
		x"30",	--1725
		x"0f",	--1726
		x"ee",	--1727
		x"0b",	--1728
		x"0a",	--1729
		x"0b",	--1730
		x"0a",	--1731
		x"8f",	--1732
		x"00",	--1733
		x"8f",	--1734
		x"02",	--1735
		x"8f",	--1736
		x"04",	--1737
		x"0c",	--1738
		x"0d",	--1739
		x"3e",	--1740
		x"00",	--1741
		x"3f",	--1742
		x"6e",	--1743
		x"b0",	--1744
		x"14",	--1745
		x"8b",	--1746
		x"02",	--1747
		x"02",	--1748
		x"32",	--1749
		x"03",	--1750
		x"82",	--1751
		x"32",	--1752
		x"b2",	--1753
		x"18",	--1754
		x"38",	--1755
		x"9b",	--1756
		x"3a",	--1757
		x"06",	--1758
		x"32",	--1759
		x"0f",	--1760
		x"3a",	--1761
		x"3b",	--1762
		x"30",	--1763
		x"0b",	--1764
		x"09",	--1765
		x"08",	--1766
		x"8f",	--1767
		x"06",	--1768
		x"bf",	--1769
		x"00",	--1770
		x"08",	--1771
		x"2b",	--1772
		x"1e",	--1773
		x"02",	--1774
		x"0f",	--1775
		x"b0",	--1776
		x"ae",	--1777
		x"0c",	--1778
		x"3d",	--1779
		x"00",	--1780
		x"b0",	--1781
		x"14",	--1782
		x"08",	--1783
		x"09",	--1784
		x"1e",	--1785
		x"06",	--1786
		x"0f",	--1787
		x"b0",	--1788
		x"ae",	--1789
		x"0c",	--1790
		x"0d",	--1791
		x"0e",	--1792
		x"0f",	--1793
		x"b0",	--1794
		x"c4",	--1795
		x"b0",	--1796
		x"a4",	--1797
		x"8b",	--1798
		x"04",	--1799
		x"9b",	--1800
		x"00",	--1801
		x"38",	--1802
		x"39",	--1803
		x"3b",	--1804
		x"30",	--1805
		x"0b",	--1806
		x"0a",	--1807
		x"09",	--1808
		x"0a",	--1809
		x"0b",	--1810
		x"8f",	--1811
		x"06",	--1812
		x"8f",	--1813
		x"08",	--1814
		x"29",	--1815
		x"1e",	--1816
		x"02",	--1817
		x"0f",	--1818
		x"b0",	--1819
		x"ae",	--1820
		x"0c",	--1821
		x"0d",	--1822
		x"0e",	--1823
		x"0f",	--1824
		x"b0",	--1825
		x"14",	--1826
		x"0a",	--1827
		x"0b",	--1828
		x"1e",	--1829
		x"06",	--1830
		x"0f",	--1831
		x"b0",	--1832
		x"ae",	--1833
		x"0c",	--1834
		x"0d",	--1835
		x"0e",	--1836
		x"0f",	--1837
		x"b0",	--1838
		x"c4",	--1839
		x"b0",	--1840
		x"a4",	--1841
		x"89",	--1842
		x"04",	--1843
		x"39",	--1844
		x"3a",	--1845
		x"3b",	--1846
		x"30",	--1847
		x"2f",	--1848
		x"8f",	--1849
		x"04",	--1850
		x"30",	--1851
		x"0b",	--1852
		x"0a",	--1853
		x"92",	--1854
		x"14",	--1855
		x"14",	--1856
		x"3b",	--1857
		x"72",	--1858
		x"0a",	--1859
		x"2b",	--1860
		x"5f",	--1861
		x"fc",	--1862
		x"8f",	--1863
		x"0f",	--1864
		x"30",	--1865
		x"9d",	--1866
		x"b0",	--1867
		x"f4",	--1868
		x"31",	--1869
		x"06",	--1870
		x"1a",	--1871
		x"3b",	--1872
		x"06",	--1873
		x"1a",	--1874
		x"14",	--1875
		x"ef",	--1876
		x"0f",	--1877
		x"3a",	--1878
		x"3b",	--1879
		x"30",	--1880
		x"1e",	--1881
		x"14",	--1882
		x"3e",	--1883
		x"20",	--1884
		x"12",	--1885
		x"0f",	--1886
		x"0f",	--1887
		x"0f",	--1888
		x"0f",	--1889
		x"3f",	--1890
		x"6e",	--1891
		x"ff",	--1892
		x"68",	--1893
		x"00",	--1894
		x"bf",	--1895
		x"78",	--1896
		x"02",	--1897
		x"bf",	--1898
		x"06",	--1899
		x"04",	--1900
		x"1e",	--1901
		x"82",	--1902
		x"14",	--1903
		x"30",	--1904
		x"0b",	--1905
		x"1b",	--1906
		x"14",	--1907
		x"3b",	--1908
		x"20",	--1909
		x"12",	--1910
		x"0c",	--1911
		x"0c",	--1912
		x"0c",	--1913
		x"0c",	--1914
		x"3c",	--1915
		x"6e",	--1916
		x"cc",	--1917
		x"00",	--1918
		x"8c",	--1919
		x"02",	--1920
		x"8c",	--1921
		x"04",	--1922
		x"1b",	--1923
		x"82",	--1924
		x"14",	--1925
		x"0f",	--1926
		x"3b",	--1927
		x"30",	--1928
		x"3f",	--1929
		x"fc",	--1930
		x"0b",	--1931
		x"31",	--1932
		x"f0",	--1933
		x"1b",	--1934
		x"14",	--1935
		x"1b",	--1936
		x"0f",	--1937
		x"5f",	--1938
		x"6e",	--1939
		x"16",	--1940
		x"3d",	--1941
		x"74",	--1942
		x"0c",	--1943
		x"05",	--1944
		x"3d",	--1945
		x"06",	--1946
		x"cd",	--1947
		x"fa",	--1948
		x"0e",	--1949
		x"1c",	--1950
		x"0c",	--1951
		x"f8",	--1952
		x"30",	--1953
		x"a5",	--1954
		x"b0",	--1955
		x"f4",	--1956
		x"21",	--1957
		x"3f",	--1958
		x"31",	--1959
		x"10",	--1960
		x"3b",	--1961
		x"30",	--1962
		x"0c",	--1963
		x"81",	--1964
		x"00",	--1965
		x"6d",	--1966
		x"4d",	--1967
		x"24",	--1968
		x"1e",	--1969
		x"1f",	--1970
		x"06",	--1971
		x"6d",	--1972
		x"4d",	--1973
		x"11",	--1974
		x"1e",	--1975
		x"3f",	--1976
		x"0e",	--1977
		x"7d",	--1978
		x"20",	--1979
		x"f7",	--1980
		x"ce",	--1981
		x"ff",	--1982
		x"0d",	--1983
		x"0d",	--1984
		x"0d",	--1985
		x"8d",	--1986
		x"00",	--1987
		x"1f",	--1988
		x"6d",	--1989
		x"4d",	--1990
		x"ef",	--1991
		x"0e",	--1992
		x"0e",	--1993
		x"0c",	--1994
		x"0c",	--1995
		x"3c",	--1996
		x"6e",	--1997
		x"0e",	--1998
		x"9c",	--1999
		x"02",	--2000
		x"31",	--2001
		x"10",	--2002
		x"3b",	--2003
		x"30",	--2004
		x"1f",	--2005
		x"f1",	--2006
		x"b2",	--2007
		x"d2",	--2008
		x"60",	--2009
		x"b2",	--2010
		x"b8",	--2011
		x"72",	--2012
		x"0f",	--2013
		x"30",	--2014
		x"0b",	--2015
		x"0b",	--2016
		x"1f",	--2017
		x"16",	--2018
		x"3f",	--2019
		x"20",	--2020
		x"19",	--2021
		x"0c",	--2022
		x"0c",	--2023
		x"0d",	--2024
		x"0d",	--2025
		x"0d",	--2026
		x"0d",	--2027
		x"0d",	--2028
		x"3d",	--2029
		x"2e",	--2030
		x"8d",	--2031
		x"00",	--2032
		x"8d",	--2033
		x"02",	--2034
		x"8d",	--2035
		x"08",	--2036
		x"8d",	--2037
		x"0a",	--2038
		x"8d",	--2039
		x"0c",	--2040
		x"0e",	--2041
		x"1e",	--2042
		x"82",	--2043
		x"16",	--2044
		x"3b",	--2045
		x"30",	--2046
		x"3f",	--2047
		x"fc",	--2048
		x"0f",	--2049
		x"0c",	--2050
		x"0c",	--2051
		x"0c",	--2052
		x"0c",	--2053
		x"0c",	--2054
		x"3c",	--2055
		x"2e",	--2056
		x"8c",	--2057
		x"02",	--2058
		x"8c",	--2059
		x"04",	--2060
		x"8c",	--2061
		x"06",	--2062
		x"8c",	--2063
		x"08",	--2064
		x"9c",	--2065
		x"00",	--2066
		x"0f",	--2067
		x"30",	--2068
		x"0f",	--2069
		x"0e",	--2070
		x"0e",	--2071
		x"0e",	--2072
		x"0e",	--2073
		x"0e",	--2074
		x"8e",	--2075
		x"2e",	--2076
		x"0f",	--2077
		x"30",	--2078
		x"0f",	--2079
		x"0e",	--2080
		x"0d",	--2081
		x"0c",	--2082
		x"0b",	--2083
		x"0a",	--2084
		x"09",	--2085
		x"08",	--2086
		x"07",	--2087
		x"92",	--2088
		x"16",	--2089
		x"33",	--2090
		x"3a",	--2091
		x"2e",	--2092
		x"0b",	--2093
		x"2b",	--2094
		x"08",	--2095
		x"38",	--2096
		x"07",	--2097
		x"37",	--2098
		x"06",	--2099
		x"09",	--2100
		x"0f",	--2101
		x"1f",	--2102
		x"8b",	--2103
		x"00",	--2104
		x"19",	--2105
		x"3a",	--2106
		x"0e",	--2107
		x"3b",	--2108
		x"0e",	--2109
		x"38",	--2110
		x"0e",	--2111
		x"37",	--2112
		x"0e",	--2113
		x"19",	--2114
		x"16",	--2115
		x"19",	--2116
		x"8a",	--2117
		x"00",	--2118
		x"f1",	--2119
		x"2f",	--2120
		x"1f",	--2121
		x"02",	--2122
		x"ea",	--2123
		x"8b",	--2124
		x"00",	--2125
		x"1f",	--2126
		x"0a",	--2127
		x"9b",	--2128
		x"08",	--2129
		x"88",	--2130
		x"00",	--2131
		x"e4",	--2132
		x"2f",	--2133
		x"1f",	--2134
		x"87",	--2135
		x"00",	--2136
		x"2f",	--2137
		x"de",	--2138
		x"8a",	--2139
		x"00",	--2140
		x"db",	--2141
		x"b2",	--2142
		x"fe",	--2143
		x"60",	--2144
		x"37",	--2145
		x"38",	--2146
		x"39",	--2147
		x"3a",	--2148
		x"3b",	--2149
		x"3c",	--2150
		x"3d",	--2151
		x"3e",	--2152
		x"3f",	--2153
		x"00",	--2154
		x"8f",	--2155
		x"00",	--2156
		x"0f",	--2157
		x"30",	--2158
		x"2f",	--2159
		x"2e",	--2160
		x"1f",	--2161
		x"02",	--2162
		x"30",	--2163
		x"8f",	--2164
		x"00",	--2165
		x"30",	--2166
		x"8f",	--2167
		x"00",	--2168
		x"3f",	--2169
		x"e8",	--2170
		x"b0",	--2171
		x"be",	--2172
		x"82",	--2173
		x"0c",	--2174
		x"0f",	--2175
		x"30",	--2176
		x"0c",	--2177
		x"2f",	--2178
		x"8f",	--2179
		x"00",	--2180
		x"1d",	--2181
		x"0e",	--2182
		x"1f",	--2183
		x"0c",	--2184
		x"b0",	--2185
		x"02",	--2186
		x"30",	--2187
		x"5e",	--2188
		x"81",	--2189
		x"3e",	--2190
		x"fc",	--2191
		x"c2",	--2192
		x"84",	--2193
		x"0f",	--2194
		x"30",	--2195
		x"3f",	--2196
		x"0f",	--2197
		x"5f",	--2198
		x"64",	--2199
		x"8f",	--2200
		x"b0",	--2201
		x"18",	--2202
		x"30",	--2203
		x"0b",	--2204
		x"0b",	--2205
		x"0e",	--2206
		x"0e",	--2207
		x"0e",	--2208
		x"0e",	--2209
		x"0e",	--2210
		x"0f",	--2211
		x"b0",	--2212
		x"28",	--2213
		x"0f",	--2214
		x"b0",	--2215
		x"28",	--2216
		x"3b",	--2217
		x"30",	--2218
		x"0b",	--2219
		x"0a",	--2220
		x"0a",	--2221
		x"3b",	--2222
		x"07",	--2223
		x"0e",	--2224
		x"4d",	--2225
		x"7d",	--2226
		x"0f",	--2227
		x"03",	--2228
		x"0e",	--2229
		x"7d",	--2230
		x"fd",	--2231
		x"1e",	--2232
		x"0a",	--2233
		x"3f",	--2234
		x"31",	--2235
		x"b0",	--2236
		x"18",	--2237
		x"3b",	--2238
		x"3b",	--2239
		x"ef",	--2240
		x"3a",	--2241
		x"3b",	--2242
		x"30",	--2243
		x"3f",	--2244
		x"30",	--2245
		x"f5",	--2246
		x"0b",	--2247
		x"0b",	--2248
		x"0e",	--2249
		x"8e",	--2250
		x"8e",	--2251
		x"0f",	--2252
		x"b0",	--2253
		x"38",	--2254
		x"0f",	--2255
		x"b0",	--2256
		x"38",	--2257
		x"3b",	--2258
		x"30",	--2259
		x"0b",	--2260
		x"0a",	--2261
		x"0a",	--2262
		x"0b",	--2263
		x"0d",	--2264
		x"8d",	--2265
		x"8d",	--2266
		x"0f",	--2267
		x"b0",	--2268
		x"38",	--2269
		x"0f",	--2270
		x"b0",	--2271
		x"38",	--2272
		x"0c",	--2273
		x"0d",	--2274
		x"8d",	--2275
		x"8c",	--2276
		x"4d",	--2277
		x"0d",	--2278
		x"0f",	--2279
		x"b0",	--2280
		x"38",	--2281
		x"0f",	--2282
		x"b0",	--2283
		x"38",	--2284
		x"3a",	--2285
		x"3b",	--2286
		x"30",	--2287
		x"0b",	--2288
		x"0a",	--2289
		x"09",	--2290
		x"0a",	--2291
		x"0e",	--2292
		x"19",	--2293
		x"09",	--2294
		x"39",	--2295
		x"0b",	--2296
		x"0d",	--2297
		x"0d",	--2298
		x"6f",	--2299
		x"8f",	--2300
		x"b0",	--2301
		x"38",	--2302
		x"0b",	--2303
		x"0e",	--2304
		x"1b",	--2305
		x"3b",	--2306
		x"07",	--2307
		x"05",	--2308
		x"3f",	--2309
		x"20",	--2310
		x"b0",	--2311
		x"18",	--2312
		x"ef",	--2313
		x"3f",	--2314
		x"3a",	--2315
		x"b0",	--2316
		x"18",	--2317
		x"ea",	--2318
		x"39",	--2319
		x"3a",	--2320
		x"3b",	--2321
		x"30",	--2322
		x"0b",	--2323
		x"0a",	--2324
		x"09",	--2325
		x"0a",	--2326
		x"0e",	--2327
		x"17",	--2328
		x"09",	--2329
		x"39",	--2330
		x"0b",	--2331
		x"6f",	--2332
		x"8f",	--2333
		x"b0",	--2334
		x"28",	--2335
		x"0b",	--2336
		x"0e",	--2337
		x"1b",	--2338
		x"3b",	--2339
		x"07",	--2340
		x"f6",	--2341
		x"3f",	--2342
		x"20",	--2343
		x"b0",	--2344
		x"18",	--2345
		x"6f",	--2346
		x"8f",	--2347
		x"b0",	--2348
		x"28",	--2349
		x"0b",	--2350
		x"f2",	--2351
		x"39",	--2352
		x"3a",	--2353
		x"3b",	--2354
		x"30",	--2355
		x"0b",	--2356
		x"0a",	--2357
		x"09",	--2358
		x"31",	--2359
		x"ec",	--2360
		x"0b",	--2361
		x"0f",	--2362
		x"34",	--2363
		x"3b",	--2364
		x"0a",	--2365
		x"38",	--2366
		x"09",	--2367
		x"0a",	--2368
		x"0a",	--2369
		x"3e",	--2370
		x"0a",	--2371
		x"0f",	--2372
		x"b0",	--2373
		x"cc",	--2374
		x"7f",	--2375
		x"30",	--2376
		x"ca",	--2377
		x"00",	--2378
		x"19",	--2379
		x"3e",	--2380
		x"0a",	--2381
		x"0f",	--2382
		x"b0",	--2383
		x"9a",	--2384
		x"0b",	--2385
		x"3f",	--2386
		x"0a",	--2387
		x"eb",	--2388
		x"0a",	--2389
		x"1a",	--2390
		x"09",	--2391
		x"3e",	--2392
		x"0a",	--2393
		x"0f",	--2394
		x"b0",	--2395
		x"cc",	--2396
		x"7f",	--2397
		x"30",	--2398
		x"c9",	--2399
		x"00",	--2400
		x"3a",	--2401
		x"0f",	--2402
		x"0f",	--2403
		x"6f",	--2404
		x"8f",	--2405
		x"b0",	--2406
		x"18",	--2407
		x"0a",	--2408
		x"f7",	--2409
		x"31",	--2410
		x"14",	--2411
		x"39",	--2412
		x"3a",	--2413
		x"3b",	--2414
		x"30",	--2415
		x"3f",	--2416
		x"2d",	--2417
		x"b0",	--2418
		x"18",	--2419
		x"3b",	--2420
		x"1b",	--2421
		x"c5",	--2422
		x"1a",	--2423
		x"09",	--2424
		x"dd",	--2425
		x"0b",	--2426
		x"0a",	--2427
		x"09",	--2428
		x"0b",	--2429
		x"3b",	--2430
		x"39",	--2431
		x"6f",	--2432
		x"4f",	--2433
		x"0b",	--2434
		x"1a",	--2435
		x"8f",	--2436
		x"b0",	--2437
		x"18",	--2438
		x"0a",	--2439
		x"09",	--2440
		x"19",	--2441
		x"5f",	--2442
		x"01",	--2443
		x"4f",	--2444
		x"10",	--2445
		x"7f",	--2446
		x"25",	--2447
		x"f3",	--2448
		x"0a",	--2449
		x"1a",	--2450
		x"5f",	--2451
		x"01",	--2452
		x"7f",	--2453
		x"db",	--2454
		x"7f",	--2455
		x"54",	--2456
		x"ee",	--2457
		x"4f",	--2458
		x"0f",	--2459
		x"10",	--2460
		x"bc",	--2461
		x"39",	--2462
		x"3a",	--2463
		x"3b",	--2464
		x"30",	--2465
		x"09",	--2466
		x"29",	--2467
		x"1e",	--2468
		x"02",	--2469
		x"2f",	--2470
		x"b0",	--2471
		x"e0",	--2472
		x"0b",	--2473
		x"dd",	--2474
		x"09",	--2475
		x"29",	--2476
		x"2f",	--2477
		x"b0",	--2478
		x"8e",	--2479
		x"0b",	--2480
		x"d6",	--2481
		x"0f",	--2482
		x"2b",	--2483
		x"29",	--2484
		x"6f",	--2485
		x"4f",	--2486
		x"d0",	--2487
		x"19",	--2488
		x"8f",	--2489
		x"b0",	--2490
		x"18",	--2491
		x"7f",	--2492
		x"4f",	--2493
		x"fa",	--2494
		x"c8",	--2495
		x"09",	--2496
		x"29",	--2497
		x"1e",	--2498
		x"02",	--2499
		x"2f",	--2500
		x"b0",	--2501
		x"26",	--2502
		x"0b",	--2503
		x"bf",	--2504
		x"09",	--2505
		x"29",	--2506
		x"2e",	--2507
		x"0f",	--2508
		x"8f",	--2509
		x"8f",	--2510
		x"8f",	--2511
		x"8f",	--2512
		x"b0",	--2513
		x"a8",	--2514
		x"0b",	--2515
		x"b3",	--2516
		x"09",	--2517
		x"29",	--2518
		x"2f",	--2519
		x"b0",	--2520
		x"68",	--2521
		x"0b",	--2522
		x"ac",	--2523
		x"09",	--2524
		x"29",	--2525
		x"2f",	--2526
		x"b0",	--2527
		x"18",	--2528
		x"0b",	--2529
		x"a5",	--2530
		x"09",	--2531
		x"29",	--2532
		x"2f",	--2533
		x"b0",	--2534
		x"38",	--2535
		x"0b",	--2536
		x"9e",	--2537
		x"09",	--2538
		x"29",	--2539
		x"2f",	--2540
		x"b0",	--2541
		x"56",	--2542
		x"0b",	--2543
		x"97",	--2544
		x"3f",	--2545
		x"25",	--2546
		x"b0",	--2547
		x"18",	--2548
		x"92",	--2549
		x"0f",	--2550
		x"0e",	--2551
		x"1f",	--2552
		x"18",	--2553
		x"df",	--2554
		x"85",	--2555
		x"ee",	--2556
		x"1f",	--2557
		x"18",	--2558
		x"3f",	--2559
		x"3f",	--2560
		x"13",	--2561
		x"92",	--2562
		x"18",	--2563
		x"1e",	--2564
		x"18",	--2565
		x"1f",	--2566
		x"1a",	--2567
		x"0e",	--2568
		x"02",	--2569
		x"92",	--2570
		x"1a",	--2571
		x"f2",	--2572
		x"10",	--2573
		x"81",	--2574
		x"3e",	--2575
		x"3f",	--2576
		x"b1",	--2577
		x"f0",	--2578
		x"00",	--2579
		x"00",	--2580
		x"82",	--2581
		x"18",	--2582
		x"ec",	--2583
		x"0c",	--2584
		x"0d",	--2585
		x"3e",	--2586
		x"00",	--2587
		x"3f",	--2588
		x"6e",	--2589
		x"b0",	--2590
		x"d4",	--2591
		x"3e",	--2592
		x"82",	--2593
		x"82",	--2594
		x"f2",	--2595
		x"11",	--2596
		x"80",	--2597
		x"30",	--2598
		x"1e",	--2599
		x"18",	--2600
		x"1f",	--2601
		x"1a",	--2602
		x"0e",	--2603
		x"05",	--2604
		x"1f",	--2605
		x"18",	--2606
		x"1f",	--2607
		x"1a",	--2608
		x"30",	--2609
		x"1d",	--2610
		x"18",	--2611
		x"1e",	--2612
		x"1a",	--2613
		x"3f",	--2614
		x"40",	--2615
		x"0f",	--2616
		x"0f",	--2617
		x"30",	--2618
		x"1f",	--2619
		x"1a",	--2620
		x"5f",	--2621
		x"ee",	--2622
		x"1d",	--2623
		x"1a",	--2624
		x"1e",	--2625
		x"18",	--2626
		x"0d",	--2627
		x"0b",	--2628
		x"1e",	--2629
		x"1a",	--2630
		x"3e",	--2631
		x"3f",	--2632
		x"03",	--2633
		x"82",	--2634
		x"1a",	--2635
		x"30",	--2636
		x"92",	--2637
		x"1a",	--2638
		x"30",	--2639
		x"4f",	--2640
		x"30",	--2641
		x"0b",	--2642
		x"0a",	--2643
		x"0a",	--2644
		x"0b",	--2645
		x"0c",	--2646
		x"3d",	--2647
		x"00",	--2648
		x"b0",	--2649
		x"d8",	--2650
		x"0f",	--2651
		x"07",	--2652
		x"0e",	--2653
		x"0f",	--2654
		x"b0",	--2655
		x"1e",	--2656
		x"3a",	--2657
		x"3b",	--2658
		x"30",	--2659
		x"0c",	--2660
		x"3d",	--2661
		x"00",	--2662
		x"0e",	--2663
		x"0f",	--2664
		x"b0",	--2665
		x"c4",	--2666
		x"b0",	--2667
		x"1e",	--2668
		x"0e",	--2669
		x"3f",	--2670
		x"00",	--2671
		x"3a",	--2672
		x"3b",	--2673
		x"30",	--2674
		x"0b",	--2675
		x"0a",	--2676
		x"09",	--2677
		x"08",	--2678
		x"07",	--2679
		x"06",	--2680
		x"05",	--2681
		x"04",	--2682
		x"31",	--2683
		x"fa",	--2684
		x"08",	--2685
		x"6b",	--2686
		x"6b",	--2687
		x"67",	--2688
		x"6c",	--2689
		x"6c",	--2690
		x"e9",	--2691
		x"6b",	--2692
		x"02",	--2693
		x"30",	--2694
		x"66",	--2695
		x"6c",	--2696
		x"e3",	--2697
		x"6c",	--2698
		x"bb",	--2699
		x"6b",	--2700
		x"df",	--2701
		x"91",	--2702
		x"02",	--2703
		x"00",	--2704
		x"1b",	--2705
		x"02",	--2706
		x"14",	--2707
		x"04",	--2708
		x"15",	--2709
		x"06",	--2710
		x"16",	--2711
		x"04",	--2712
		x"17",	--2713
		x"06",	--2714
		x"2c",	--2715
		x"0c",	--2716
		x"09",	--2717
		x"0c",	--2718
		x"bf",	--2719
		x"39",	--2720
		x"20",	--2721
		x"50",	--2722
		x"1c",	--2723
		x"d7",	--2724
		x"81",	--2725
		x"02",	--2726
		x"81",	--2727
		x"04",	--2728
		x"4c",	--2729
		x"7c",	--2730
		x"1f",	--2731
		x"0b",	--2732
		x"0a",	--2733
		x"0b",	--2734
		x"12",	--2735
		x"0b",	--2736
		x"0a",	--2737
		x"7c",	--2738
		x"fb",	--2739
		x"81",	--2740
		x"02",	--2741
		x"81",	--2742
		x"04",	--2743
		x"1c",	--2744
		x"0d",	--2745
		x"79",	--2746
		x"1f",	--2747
		x"04",	--2748
		x"0c",	--2749
		x"0d",	--2750
		x"79",	--2751
		x"fc",	--2752
		x"3c",	--2753
		x"3d",	--2754
		x"0c",	--2755
		x"0d",	--2756
		x"1a",	--2757
		x"0b",	--2758
		x"0c",	--2759
		x"02",	--2760
		x"0d",	--2761
		x"e5",	--2762
		x"16",	--2763
		x"02",	--2764
		x"17",	--2765
		x"04",	--2766
		x"06",	--2767
		x"07",	--2768
		x"5f",	--2769
		x"01",	--2770
		x"5f",	--2771
		x"01",	--2772
		x"28",	--2773
		x"c8",	--2774
		x"01",	--2775
		x"a8",	--2776
		x"02",	--2777
		x"0e",	--2778
		x"0f",	--2779
		x"0e",	--2780
		x"0f",	--2781
		x"88",	--2782
		x"04",	--2783
		x"88",	--2784
		x"06",	--2785
		x"f8",	--2786
		x"03",	--2787
		x"00",	--2788
		x"0f",	--2789
		x"4d",	--2790
		x"0f",	--2791
		x"31",	--2792
		x"06",	--2793
		x"34",	--2794
		x"35",	--2795
		x"36",	--2796
		x"37",	--2797
		x"38",	--2798
		x"39",	--2799
		x"3a",	--2800
		x"3b",	--2801
		x"30",	--2802
		x"2b",	--2803
		x"67",	--2804
		x"81",	--2805
		x"00",	--2806
		x"04",	--2807
		x"05",	--2808
		x"5f",	--2809
		x"01",	--2810
		x"5f",	--2811
		x"01",	--2812
		x"d8",	--2813
		x"4f",	--2814
		x"68",	--2815
		x"0e",	--2816
		x"0f",	--2817
		x"0e",	--2818
		x"0f",	--2819
		x"0f",	--2820
		x"69",	--2821
		x"c8",	--2822
		x"01",	--2823
		x"a8",	--2824
		x"02",	--2825
		x"88",	--2826
		x"04",	--2827
		x"88",	--2828
		x"06",	--2829
		x"0c",	--2830
		x"0d",	--2831
		x"3c",	--2832
		x"3d",	--2833
		x"3d",	--2834
		x"ff",	--2835
		x"05",	--2836
		x"3d",	--2837
		x"00",	--2838
		x"17",	--2839
		x"3c",	--2840
		x"15",	--2841
		x"1b",	--2842
		x"02",	--2843
		x"3b",	--2844
		x"0e",	--2845
		x"0f",	--2846
		x"0a",	--2847
		x"3b",	--2848
		x"0c",	--2849
		x"0d",	--2850
		x"3c",	--2851
		x"3d",	--2852
		x"3d",	--2853
		x"ff",	--2854
		x"f5",	--2855
		x"3c",	--2856
		x"88",	--2857
		x"04",	--2858
		x"88",	--2859
		x"06",	--2860
		x"88",	--2861
		x"02",	--2862
		x"f8",	--2863
		x"03",	--2864
		x"00",	--2865
		x"0f",	--2866
		x"b3",	--2867
		x"0c",	--2868
		x"0d",	--2869
		x"1c",	--2870
		x"0d",	--2871
		x"12",	--2872
		x"0f",	--2873
		x"0e",	--2874
		x"0a",	--2875
		x"0b",	--2876
		x"0a",	--2877
		x"0b",	--2878
		x"88",	--2879
		x"04",	--2880
		x"88",	--2881
		x"06",	--2882
		x"98",	--2883
		x"02",	--2884
		x"0f",	--2885
		x"a1",	--2886
		x"6b",	--2887
		x"9f",	--2888
		x"ad",	--2889
		x"00",	--2890
		x"9d",	--2891
		x"02",	--2892
		x"02",	--2893
		x"9d",	--2894
		x"04",	--2895
		x"04",	--2896
		x"9d",	--2897
		x"06",	--2898
		x"06",	--2899
		x"5e",	--2900
		x"01",	--2901
		x"5e",	--2902
		x"01",	--2903
		x"cd",	--2904
		x"01",	--2905
		x"0f",	--2906
		x"8c",	--2907
		x"06",	--2908
		x"07",	--2909
		x"9a",	--2910
		x"39",	--2911
		x"19",	--2912
		x"39",	--2913
		x"20",	--2914
		x"8f",	--2915
		x"3e",	--2916
		x"3c",	--2917
		x"b6",	--2918
		x"c1",	--2919
		x"0e",	--2920
		x"0f",	--2921
		x"0e",	--2922
		x"0f",	--2923
		x"97",	--2924
		x"0f",	--2925
		x"79",	--2926
		x"d8",	--2927
		x"01",	--2928
		x"a8",	--2929
		x"02",	--2930
		x"3e",	--2931
		x"3f",	--2932
		x"1e",	--2933
		x"0f",	--2934
		x"88",	--2935
		x"04",	--2936
		x"88",	--2937
		x"06",	--2938
		x"92",	--2939
		x"0c",	--2940
		x"7b",	--2941
		x"81",	--2942
		x"00",	--2943
		x"81",	--2944
		x"02",	--2945
		x"81",	--2946
		x"04",	--2947
		x"4d",	--2948
		x"7d",	--2949
		x"1f",	--2950
		x"0c",	--2951
		x"4b",	--2952
		x"0c",	--2953
		x"0d",	--2954
		x"12",	--2955
		x"0d",	--2956
		x"0c",	--2957
		x"7b",	--2958
		x"fb",	--2959
		x"81",	--2960
		x"02",	--2961
		x"81",	--2962
		x"04",	--2963
		x"1c",	--2964
		x"0d",	--2965
		x"79",	--2966
		x"1f",	--2967
		x"04",	--2968
		x"0c",	--2969
		x"0d",	--2970
		x"79",	--2971
		x"fc",	--2972
		x"3c",	--2973
		x"3d",	--2974
		x"0c",	--2975
		x"0d",	--2976
		x"1a",	--2977
		x"0b",	--2978
		x"0c",	--2979
		x"04",	--2980
		x"0d",	--2981
		x"02",	--2982
		x"0a",	--2983
		x"0b",	--2984
		x"14",	--2985
		x"02",	--2986
		x"15",	--2987
		x"04",	--2988
		x"04",	--2989
		x"05",	--2990
		x"49",	--2991
		x"0a",	--2992
		x"0b",	--2993
		x"18",	--2994
		x"6c",	--2995
		x"33",	--2996
		x"df",	--2997
		x"01",	--2998
		x"01",	--2999
		x"2f",	--3000
		x"3f",	--3001
		x"76",	--3002
		x"2c",	--3003
		x"31",	--3004
		x"e0",	--3005
		x"81",	--3006
		x"04",	--3007
		x"81",	--3008
		x"06",	--3009
		x"81",	--3010
		x"00",	--3011
		x"81",	--3012
		x"02",	--3013
		x"0e",	--3014
		x"3e",	--3015
		x"18",	--3016
		x"0f",	--3017
		x"2f",	--3018
		x"b0",	--3019
		x"e0",	--3020
		x"0e",	--3021
		x"3e",	--3022
		x"10",	--3023
		x"0f",	--3024
		x"b0",	--3025
		x"e0",	--3026
		x"0d",	--3027
		x"3d",	--3028
		x"0e",	--3029
		x"3e",	--3030
		x"10",	--3031
		x"0f",	--3032
		x"3f",	--3033
		x"18",	--3034
		x"b0",	--3035
		x"e6",	--3036
		x"b0",	--3037
		x"02",	--3038
		x"31",	--3039
		x"20",	--3040
		x"30",	--3041
		x"31",	--3042
		x"e0",	--3043
		x"81",	--3044
		x"04",	--3045
		x"81",	--3046
		x"06",	--3047
		x"81",	--3048
		x"00",	--3049
		x"81",	--3050
		x"02",	--3051
		x"0e",	--3052
		x"3e",	--3053
		x"18",	--3054
		x"0f",	--3055
		x"2f",	--3056
		x"b0",	--3057
		x"e0",	--3058
		x"0e",	--3059
		x"3e",	--3060
		x"10",	--3061
		x"0f",	--3062
		x"b0",	--3063
		x"e0",	--3064
		x"d1",	--3065
		x"11",	--3066
		x"0d",	--3067
		x"3d",	--3068
		x"0e",	--3069
		x"3e",	--3070
		x"10",	--3071
		x"0f",	--3072
		x"3f",	--3073
		x"18",	--3074
		x"b0",	--3075
		x"e6",	--3076
		x"b0",	--3077
		x"02",	--3078
		x"31",	--3079
		x"20",	--3080
		x"30",	--3081
		x"0b",	--3082
		x"0a",	--3083
		x"09",	--3084
		x"08",	--3085
		x"07",	--3086
		x"06",	--3087
		x"05",	--3088
		x"04",	--3089
		x"31",	--3090
		x"dc",	--3091
		x"81",	--3092
		x"04",	--3093
		x"81",	--3094
		x"06",	--3095
		x"81",	--3096
		x"00",	--3097
		x"81",	--3098
		x"02",	--3099
		x"0e",	--3100
		x"3e",	--3101
		x"18",	--3102
		x"0f",	--3103
		x"2f",	--3104
		x"b0",	--3105
		x"e0",	--3106
		x"0e",	--3107
		x"3e",	--3108
		x"10",	--3109
		x"0f",	--3110
		x"b0",	--3111
		x"e0",	--3112
		x"5f",	--3113
		x"18",	--3114
		x"6f",	--3115
		x"b6",	--3116
		x"5e",	--3117
		x"10",	--3118
		x"6e",	--3119
		x"d9",	--3120
		x"6f",	--3121
		x"ae",	--3122
		x"6e",	--3123
		x"e2",	--3124
		x"6f",	--3125
		x"ac",	--3126
		x"6e",	--3127
		x"d1",	--3128
		x"14",	--3129
		x"1c",	--3130
		x"15",	--3131
		x"1e",	--3132
		x"18",	--3133
		x"14",	--3134
		x"19",	--3135
		x"16",	--3136
		x"3c",	--3137
		x"20",	--3138
		x"0e",	--3139
		x"0f",	--3140
		x"06",	--3141
		x"07",	--3142
		x"81",	--3143
		x"20",	--3144
		x"81",	--3145
		x"22",	--3146
		x"0a",	--3147
		x"0b",	--3148
		x"81",	--3149
		x"20",	--3150
		x"08",	--3151
		x"08",	--3152
		x"09",	--3153
		x"12",	--3154
		x"05",	--3155
		x"04",	--3156
		x"b1",	--3157
		x"20",	--3158
		x"19",	--3159
		x"14",	--3160
		x"0d",	--3161
		x"0a",	--3162
		x"0b",	--3163
		x"0e",	--3164
		x"0f",	--3165
		x"1c",	--3166
		x"0d",	--3167
		x"0b",	--3168
		x"03",	--3169
		x"0b",	--3170
		x"0c",	--3171
		x"0d",	--3172
		x"0e",	--3173
		x"0f",	--3174
		x"06",	--3175
		x"07",	--3176
		x"09",	--3177
		x"e5",	--3178
		x"16",	--3179
		x"07",	--3180
		x"e2",	--3181
		x"0a",	--3182
		x"f5",	--3183
		x"f2",	--3184
		x"81",	--3185
		x"20",	--3186
		x"81",	--3187
		x"22",	--3188
		x"0c",	--3189
		x"1a",	--3190
		x"1a",	--3191
		x"1a",	--3192
		x"12",	--3193
		x"06",	--3194
		x"26",	--3195
		x"81",	--3196
		x"0a",	--3197
		x"5d",	--3198
		x"d1",	--3199
		x"11",	--3200
		x"19",	--3201
		x"83",	--3202
		x"c1",	--3203
		x"09",	--3204
		x"0c",	--3205
		x"3c",	--3206
		x"3f",	--3207
		x"00",	--3208
		x"18",	--3209
		x"1d",	--3210
		x"0a",	--3211
		x"3d",	--3212
		x"1a",	--3213
		x"20",	--3214
		x"1b",	--3215
		x"22",	--3216
		x"0c",	--3217
		x"0e",	--3218
		x"0f",	--3219
		x"0b",	--3220
		x"2a",	--3221
		x"0a",	--3222
		x"0b",	--3223
		x"3d",	--3224
		x"3f",	--3225
		x"00",	--3226
		x"f5",	--3227
		x"81",	--3228
		x"20",	--3229
		x"81",	--3230
		x"22",	--3231
		x"81",	--3232
		x"0a",	--3233
		x"0c",	--3234
		x"0d",	--3235
		x"3c",	--3236
		x"7f",	--3237
		x"0d",	--3238
		x"3c",	--3239
		x"40",	--3240
		x"44",	--3241
		x"81",	--3242
		x"0c",	--3243
		x"81",	--3244
		x"0e",	--3245
		x"f1",	--3246
		x"03",	--3247
		x"08",	--3248
		x"0f",	--3249
		x"3f",	--3250
		x"b0",	--3251
		x"02",	--3252
		x"31",	--3253
		x"24",	--3254
		x"34",	--3255
		x"35",	--3256
		x"36",	--3257
		x"37",	--3258
		x"38",	--3259
		x"39",	--3260
		x"3a",	--3261
		x"3b",	--3262
		x"30",	--3263
		x"1e",	--3264
		x"0f",	--3265
		x"d3",	--3266
		x"3a",	--3267
		x"03",	--3268
		x"08",	--3269
		x"1e",	--3270
		x"10",	--3271
		x"1c",	--3272
		x"20",	--3273
		x"1d",	--3274
		x"22",	--3275
		x"12",	--3276
		x"0d",	--3277
		x"0c",	--3278
		x"06",	--3279
		x"07",	--3280
		x"06",	--3281
		x"37",	--3282
		x"00",	--3283
		x"81",	--3284
		x"20",	--3285
		x"81",	--3286
		x"22",	--3287
		x"12",	--3288
		x"0f",	--3289
		x"0e",	--3290
		x"1a",	--3291
		x"0f",	--3292
		x"e7",	--3293
		x"81",	--3294
		x"0a",	--3295
		x"a6",	--3296
		x"6e",	--3297
		x"36",	--3298
		x"5f",	--3299
		x"d1",	--3300
		x"11",	--3301
		x"19",	--3302
		x"20",	--3303
		x"c1",	--3304
		x"19",	--3305
		x"0f",	--3306
		x"3f",	--3307
		x"18",	--3308
		x"c5",	--3309
		x"0d",	--3310
		x"ba",	--3311
		x"0c",	--3312
		x"0d",	--3313
		x"3c",	--3314
		x"80",	--3315
		x"0d",	--3316
		x"0c",	--3317
		x"b3",	--3318
		x"0d",	--3319
		x"b1",	--3320
		x"81",	--3321
		x"20",	--3322
		x"03",	--3323
		x"81",	--3324
		x"22",	--3325
		x"ab",	--3326
		x"3e",	--3327
		x"40",	--3328
		x"0f",	--3329
		x"3e",	--3330
		x"80",	--3331
		x"3f",	--3332
		x"a4",	--3333
		x"4d",	--3334
		x"7b",	--3335
		x"4f",	--3336
		x"de",	--3337
		x"5f",	--3338
		x"d1",	--3339
		x"11",	--3340
		x"19",	--3341
		x"06",	--3342
		x"c1",	--3343
		x"11",	--3344
		x"0f",	--3345
		x"3f",	--3346
		x"10",	--3347
		x"9e",	--3348
		x"4f",	--3349
		x"f8",	--3350
		x"6f",	--3351
		x"f1",	--3352
		x"3f",	--3353
		x"76",	--3354
		x"97",	--3355
		x"0b",	--3356
		x"0a",	--3357
		x"09",	--3358
		x"08",	--3359
		x"07",	--3360
		x"31",	--3361
		x"e8",	--3362
		x"81",	--3363
		x"04",	--3364
		x"81",	--3365
		x"06",	--3366
		x"81",	--3367
		x"00",	--3368
		x"81",	--3369
		x"02",	--3370
		x"0e",	--3371
		x"3e",	--3372
		x"10",	--3373
		x"0f",	--3374
		x"2f",	--3375
		x"b0",	--3376
		x"e0",	--3377
		x"0e",	--3378
		x"3e",	--3379
		x"0f",	--3380
		x"b0",	--3381
		x"e0",	--3382
		x"5f",	--3383
		x"10",	--3384
		x"6f",	--3385
		x"5d",	--3386
		x"5e",	--3387
		x"08",	--3388
		x"6e",	--3389
		x"82",	--3390
		x"d1",	--3391
		x"09",	--3392
		x"11",	--3393
		x"6f",	--3394
		x"58",	--3395
		x"6f",	--3396
		x"56",	--3397
		x"6e",	--3398
		x"6f",	--3399
		x"6e",	--3400
		x"4c",	--3401
		x"1d",	--3402
		x"12",	--3403
		x"1d",	--3404
		x"0a",	--3405
		x"81",	--3406
		x"12",	--3407
		x"1e",	--3408
		x"14",	--3409
		x"1f",	--3410
		x"16",	--3411
		x"18",	--3412
		x"0c",	--3413
		x"19",	--3414
		x"0e",	--3415
		x"0f",	--3416
		x"1e",	--3417
		x"0e",	--3418
		x"0f",	--3419
		x"3d",	--3420
		x"81",	--3421
		x"12",	--3422
		x"37",	--3423
		x"1f",	--3424
		x"0c",	--3425
		x"3d",	--3426
		x"00",	--3427
		x"0a",	--3428
		x"0b",	--3429
		x"0b",	--3430
		x"0a",	--3431
		x"0b",	--3432
		x"0e",	--3433
		x"0f",	--3434
		x"12",	--3435
		x"0d",	--3436
		x"0c",	--3437
		x"0e",	--3438
		x"0f",	--3439
		x"37",	--3440
		x"0b",	--3441
		x"0f",	--3442
		x"f7",	--3443
		x"f2",	--3444
		x"0e",	--3445
		x"f4",	--3446
		x"ef",	--3447
		x"09",	--3448
		x"e5",	--3449
		x"0e",	--3450
		x"e3",	--3451
		x"dd",	--3452
		x"0c",	--3453
		x"0d",	--3454
		x"3c",	--3455
		x"7f",	--3456
		x"0d",	--3457
		x"3c",	--3458
		x"40",	--3459
		x"1c",	--3460
		x"81",	--3461
		x"14",	--3462
		x"81",	--3463
		x"16",	--3464
		x"0f",	--3465
		x"3f",	--3466
		x"10",	--3467
		x"b0",	--3468
		x"02",	--3469
		x"31",	--3470
		x"18",	--3471
		x"37",	--3472
		x"38",	--3473
		x"39",	--3474
		x"3a",	--3475
		x"3b",	--3476
		x"30",	--3477
		x"e1",	--3478
		x"10",	--3479
		x"0f",	--3480
		x"3f",	--3481
		x"10",	--3482
		x"f0",	--3483
		x"4f",	--3484
		x"fa",	--3485
		x"3f",	--3486
		x"76",	--3487
		x"eb",	--3488
		x"0d",	--3489
		x"e2",	--3490
		x"0c",	--3491
		x"0d",	--3492
		x"3c",	--3493
		x"80",	--3494
		x"0d",	--3495
		x"0c",	--3496
		x"db",	--3497
		x"0d",	--3498
		x"d9",	--3499
		x"0e",	--3500
		x"02",	--3501
		x"0f",	--3502
		x"d5",	--3503
		x"3a",	--3504
		x"40",	--3505
		x"0b",	--3506
		x"3a",	--3507
		x"80",	--3508
		x"3b",	--3509
		x"ce",	--3510
		x"81",	--3511
		x"14",	--3512
		x"81",	--3513
		x"16",	--3514
		x"81",	--3515
		x"12",	--3516
		x"0f",	--3517
		x"3f",	--3518
		x"10",	--3519
		x"cb",	--3520
		x"0f",	--3521
		x"3f",	--3522
		x"c8",	--3523
		x"31",	--3524
		x"e8",	--3525
		x"81",	--3526
		x"04",	--3527
		x"81",	--3528
		x"06",	--3529
		x"81",	--3530
		x"00",	--3531
		x"81",	--3532
		x"02",	--3533
		x"0e",	--3534
		x"3e",	--3535
		x"10",	--3536
		x"0f",	--3537
		x"2f",	--3538
		x"b0",	--3539
		x"e0",	--3540
		x"0e",	--3541
		x"3e",	--3542
		x"0f",	--3543
		x"b0",	--3544
		x"e0",	--3545
		x"e1",	--3546
		x"10",	--3547
		x"0d",	--3548
		x"e1",	--3549
		x"08",	--3550
		x"0a",	--3551
		x"0e",	--3552
		x"3e",	--3553
		x"0f",	--3554
		x"3f",	--3555
		x"10",	--3556
		x"b0",	--3557
		x"04",	--3558
		x"31",	--3559
		x"18",	--3560
		x"30",	--3561
		x"3f",	--3562
		x"fb",	--3563
		x"31",	--3564
		x"e8",	--3565
		x"81",	--3566
		x"04",	--3567
		x"81",	--3568
		x"06",	--3569
		x"81",	--3570
		x"00",	--3571
		x"81",	--3572
		x"02",	--3573
		x"0e",	--3574
		x"3e",	--3575
		x"10",	--3576
		x"0f",	--3577
		x"2f",	--3578
		x"b0",	--3579
		x"e0",	--3580
		x"0e",	--3581
		x"3e",	--3582
		x"0f",	--3583
		x"b0",	--3584
		x"e0",	--3585
		x"e1",	--3586
		x"10",	--3587
		x"0d",	--3588
		x"e1",	--3589
		x"08",	--3590
		x"0a",	--3591
		x"0e",	--3592
		x"3e",	--3593
		x"0f",	--3594
		x"3f",	--3595
		x"10",	--3596
		x"b0",	--3597
		x"04",	--3598
		x"31",	--3599
		x"18",	--3600
		x"30",	--3601
		x"3f",	--3602
		x"fb",	--3603
		x"31",	--3604
		x"e8",	--3605
		x"81",	--3606
		x"04",	--3607
		x"81",	--3608
		x"06",	--3609
		x"81",	--3610
		x"00",	--3611
		x"81",	--3612
		x"02",	--3613
		x"0e",	--3614
		x"3e",	--3615
		x"10",	--3616
		x"0f",	--3617
		x"2f",	--3618
		x"b0",	--3619
		x"e0",	--3620
		x"0e",	--3621
		x"3e",	--3622
		x"0f",	--3623
		x"b0",	--3624
		x"e0",	--3625
		x"e1",	--3626
		x"10",	--3627
		x"0d",	--3628
		x"e1",	--3629
		x"08",	--3630
		x"0a",	--3631
		x"0e",	--3632
		x"3e",	--3633
		x"0f",	--3634
		x"3f",	--3635
		x"10",	--3636
		x"b0",	--3637
		x"04",	--3638
		x"31",	--3639
		x"18",	--3640
		x"30",	--3641
		x"1f",	--3642
		x"fb",	--3643
		x"0b",	--3644
		x"0a",	--3645
		x"31",	--3646
		x"f1",	--3647
		x"03",	--3648
		x"00",	--3649
		x"0d",	--3650
		x"0d",	--3651
		x"0d",	--3652
		x"0d",	--3653
		x"4c",	--3654
		x"c1",	--3655
		x"01",	--3656
		x"0e",	--3657
		x"0b",	--3658
		x"0f",	--3659
		x"09",	--3660
		x"e1",	--3661
		x"00",	--3662
		x"0f",	--3663
		x"b0",	--3664
		x"02",	--3665
		x"31",	--3666
		x"3a",	--3667
		x"3b",	--3668
		x"30",	--3669
		x"b1",	--3670
		x"1e",	--3671
		x"02",	--3672
		x"4c",	--3673
		x"1b",	--3674
		x"0a",	--3675
		x"0b",	--3676
		x"81",	--3677
		x"04",	--3678
		x"81",	--3679
		x"06",	--3680
		x"0e",	--3681
		x"0f",	--3682
		x"b0",	--3683
		x"90",	--3684
		x"3f",	--3685
		x"1f",	--3686
		x"e7",	--3687
		x"81",	--3688
		x"04",	--3689
		x"81",	--3690
		x"06",	--3691
		x"4e",	--3692
		x"7e",	--3693
		x"1f",	--3694
		x"0f",	--3695
		x"3e",	--3696
		x"1e",	--3697
		x"0e",	--3698
		x"81",	--3699
		x"02",	--3700
		x"d9",	--3701
		x"0e",	--3702
		x"10",	--3703
		x"0a",	--3704
		x"0b",	--3705
		x"3a",	--3706
		x"3b",	--3707
		x"1a",	--3708
		x"0b",	--3709
		x"de",	--3710
		x"91",	--3711
		x"04",	--3712
		x"04",	--3713
		x"91",	--3714
		x"06",	--3715
		x"06",	--3716
		x"7e",	--3717
		x"f8",	--3718
		x"e8",	--3719
		x"3f",	--3720
		x"00",	--3721
		x"ed",	--3722
		x"0e",	--3723
		x"3f",	--3724
		x"00",	--3725
		x"c3",	--3726
		x"31",	--3727
		x"f4",	--3728
		x"81",	--3729
		x"00",	--3730
		x"81",	--3731
		x"02",	--3732
		x"0e",	--3733
		x"2e",	--3734
		x"0f",	--3735
		x"b0",	--3736
		x"e0",	--3737
		x"5f",	--3738
		x"04",	--3739
		x"6f",	--3740
		x"28",	--3741
		x"27",	--3742
		x"6f",	--3743
		x"07",	--3744
		x"1d",	--3745
		x"06",	--3746
		x"0d",	--3747
		x"21",	--3748
		x"3d",	--3749
		x"1f",	--3750
		x"09",	--3751
		x"c1",	--3752
		x"05",	--3753
		x"26",	--3754
		x"3e",	--3755
		x"3f",	--3756
		x"ff",	--3757
		x"31",	--3758
		x"0c",	--3759
		x"30",	--3760
		x"1e",	--3761
		x"08",	--3762
		x"1f",	--3763
		x"0a",	--3764
		x"3c",	--3765
		x"1e",	--3766
		x"4c",	--3767
		x"4d",	--3768
		x"7d",	--3769
		x"1f",	--3770
		x"0f",	--3771
		x"c1",	--3772
		x"05",	--3773
		x"ef",	--3774
		x"3e",	--3775
		x"3f",	--3776
		x"1e",	--3777
		x"0f",	--3778
		x"31",	--3779
		x"0c",	--3780
		x"30",	--3781
		x"0e",	--3782
		x"0f",	--3783
		x"31",	--3784
		x"0c",	--3785
		x"30",	--3786
		x"12",	--3787
		x"0f",	--3788
		x"0e",	--3789
		x"7d",	--3790
		x"fb",	--3791
		x"eb",	--3792
		x"0e",	--3793
		x"3f",	--3794
		x"00",	--3795
		x"31",	--3796
		x"0c",	--3797
		x"30",	--3798
		x"0b",	--3799
		x"0a",	--3800
		x"09",	--3801
		x"08",	--3802
		x"31",	--3803
		x"0a",	--3804
		x"0b",	--3805
		x"c1",	--3806
		x"01",	--3807
		x"0e",	--3808
		x"0d",	--3809
		x"0b",	--3810
		x"0b",	--3811
		x"e1",	--3812
		x"00",	--3813
		x"0f",	--3814
		x"b0",	--3815
		x"02",	--3816
		x"31",	--3817
		x"38",	--3818
		x"39",	--3819
		x"3a",	--3820
		x"3b",	--3821
		x"30",	--3822
		x"f1",	--3823
		x"03",	--3824
		x"00",	--3825
		x"b1",	--3826
		x"1e",	--3827
		x"02",	--3828
		x"81",	--3829
		x"04",	--3830
		x"81",	--3831
		x"06",	--3832
		x"0e",	--3833
		x"0f",	--3834
		x"b0",	--3835
		x"90",	--3836
		x"3f",	--3837
		x"0f",	--3838
		x"18",	--3839
		x"e5",	--3840
		x"81",	--3841
		x"04",	--3842
		x"81",	--3843
		x"06",	--3844
		x"4e",	--3845
		x"7e",	--3846
		x"1f",	--3847
		x"06",	--3848
		x"3e",	--3849
		x"1e",	--3850
		x"0e",	--3851
		x"81",	--3852
		x"02",	--3853
		x"d7",	--3854
		x"91",	--3855
		x"04",	--3856
		x"04",	--3857
		x"91",	--3858
		x"06",	--3859
		x"06",	--3860
		x"7e",	--3861
		x"f8",	--3862
		x"f1",	--3863
		x"0e",	--3864
		x"3e",	--3865
		x"1e",	--3866
		x"1c",	--3867
		x"0d",	--3868
		x"48",	--3869
		x"78",	--3870
		x"1f",	--3871
		x"04",	--3872
		x"0c",	--3873
		x"0d",	--3874
		x"78",	--3875
		x"fc",	--3876
		x"3c",	--3877
		x"3d",	--3878
		x"0c",	--3879
		x"0d",	--3880
		x"18",	--3881
		x"09",	--3882
		x"0c",	--3883
		x"04",	--3884
		x"0d",	--3885
		x"02",	--3886
		x"08",	--3887
		x"09",	--3888
		x"7e",	--3889
		x"1f",	--3890
		x"0e",	--3891
		x"0d",	--3892
		x"0e",	--3893
		x"0d",	--3894
		x"0e",	--3895
		x"81",	--3896
		x"04",	--3897
		x"81",	--3898
		x"06",	--3899
		x"3e",	--3900
		x"1e",	--3901
		x"0e",	--3902
		x"81",	--3903
		x"02",	--3904
		x"a4",	--3905
		x"12",	--3906
		x"0b",	--3907
		x"0a",	--3908
		x"7e",	--3909
		x"fb",	--3910
		x"ec",	--3911
		x"0b",	--3912
		x"0a",	--3913
		x"09",	--3914
		x"1f",	--3915
		x"17",	--3916
		x"3e",	--3917
		x"00",	--3918
		x"2c",	--3919
		x"3a",	--3920
		x"18",	--3921
		x"0b",	--3922
		x"39",	--3923
		x"0c",	--3924
		x"0d",	--3925
		x"4f",	--3926
		x"4f",	--3927
		x"17",	--3928
		x"3c",	--3929
		x"7e",	--3930
		x"6e",	--3931
		x"0f",	--3932
		x"0a",	--3933
		x"0b",	--3934
		x"0f",	--3935
		x"39",	--3936
		x"3a",	--3937
		x"3b",	--3938
		x"30",	--3939
		x"3f",	--3940
		x"00",	--3941
		x"0f",	--3942
		x"3a",	--3943
		x"0b",	--3944
		x"39",	--3945
		x"18",	--3946
		x"0c",	--3947
		x"0d",	--3948
		x"4f",	--3949
		x"4f",	--3950
		x"e9",	--3951
		x"12",	--3952
		x"0d",	--3953
		x"0c",	--3954
		x"7f",	--3955
		x"fb",	--3956
		x"e3",	--3957
		x"3a",	--3958
		x"10",	--3959
		x"0b",	--3960
		x"39",	--3961
		x"10",	--3962
		x"ef",	--3963
		x"3a",	--3964
		x"20",	--3965
		x"0b",	--3966
		x"09",	--3967
		x"ea",	--3968
		x"0b",	--3969
		x"0a",	--3970
		x"09",	--3971
		x"08",	--3972
		x"07",	--3973
		x"0d",	--3974
		x"1e",	--3975
		x"04",	--3976
		x"1f",	--3977
		x"06",	--3978
		x"5a",	--3979
		x"01",	--3980
		x"6c",	--3981
		x"6c",	--3982
		x"70",	--3983
		x"6c",	--3984
		x"6a",	--3985
		x"6c",	--3986
		x"36",	--3987
		x"0e",	--3988
		x"32",	--3989
		x"1b",	--3990
		x"02",	--3991
		x"3b",	--3992
		x"82",	--3993
		x"6d",	--3994
		x"3b",	--3995
		x"80",	--3996
		x"5e",	--3997
		x"0c",	--3998
		x"0d",	--3999
		x"3c",	--4000
		x"7f",	--4001
		x"0d",	--4002
		x"3c",	--4003
		x"40",	--4004
		x"40",	--4005
		x"3e",	--4006
		x"3f",	--4007
		x"0f",	--4008
		x"0f",	--4009
		x"4a",	--4010
		x"0d",	--4011
		x"3d",	--4012
		x"7f",	--4013
		x"12",	--4014
		x"0f",	--4015
		x"0e",	--4016
		x"12",	--4017
		x"0f",	--4018
		x"0e",	--4019
		x"12",	--4020
		x"0f",	--4021
		x"0e",	--4022
		x"12",	--4023
		x"0f",	--4024
		x"0e",	--4025
		x"12",	--4026
		x"0f",	--4027
		x"0e",	--4028
		x"12",	--4029
		x"0f",	--4030
		x"0e",	--4031
		x"12",	--4032
		x"0f",	--4033
		x"0e",	--4034
		x"3e",	--4035
		x"3f",	--4036
		x"7f",	--4037
		x"4d",	--4038
		x"05",	--4039
		x"0f",	--4040
		x"cc",	--4041
		x"4d",	--4042
		x"0e",	--4043
		x"0f",	--4044
		x"4d",	--4045
		x"0d",	--4046
		x"0d",	--4047
		x"0d",	--4048
		x"0d",	--4049
		x"0d",	--4050
		x"0d",	--4051
		x"0d",	--4052
		x"0c",	--4053
		x"3c",	--4054
		x"7f",	--4055
		x"0c",	--4056
		x"4f",	--4057
		x"0f",	--4058
		x"0f",	--4059
		x"0f",	--4060
		x"0d",	--4061
		x"0d",	--4062
		x"0f",	--4063
		x"37",	--4064
		x"38",	--4065
		x"39",	--4066
		x"3a",	--4067
		x"3b",	--4068
		x"30",	--4069
		x"0d",	--4070
		x"be",	--4071
		x"0c",	--4072
		x"0d",	--4073
		x"3c",	--4074
		x"80",	--4075
		x"0d",	--4076
		x"0c",	--4077
		x"02",	--4078
		x"0d",	--4079
		x"b8",	--4080
		x"3e",	--4081
		x"40",	--4082
		x"0f",	--4083
		x"b4",	--4084
		x"12",	--4085
		x"0f",	--4086
		x"0e",	--4087
		x"0d",	--4088
		x"3d",	--4089
		x"80",	--4090
		x"b2",	--4091
		x"7d",	--4092
		x"0e",	--4093
		x"0f",	--4094
		x"cd",	--4095
		x"0e",	--4096
		x"3f",	--4097
		x"10",	--4098
		x"3e",	--4099
		x"3f",	--4100
		x"7f",	--4101
		x"7d",	--4102
		x"c5",	--4103
		x"37",	--4104
		x"82",	--4105
		x"07",	--4106
		x"37",	--4107
		x"1a",	--4108
		x"4f",	--4109
		x"0c",	--4110
		x"0d",	--4111
		x"4b",	--4112
		x"7b",	--4113
		x"1f",	--4114
		x"05",	--4115
		x"12",	--4116
		x"0d",	--4117
		x"0c",	--4118
		x"7b",	--4119
		x"fb",	--4120
		x"18",	--4121
		x"09",	--4122
		x"77",	--4123
		x"1f",	--4124
		x"04",	--4125
		x"08",	--4126
		x"09",	--4127
		x"77",	--4128
		x"fc",	--4129
		x"38",	--4130
		x"39",	--4131
		x"08",	--4132
		x"09",	--4133
		x"1e",	--4134
		x"0f",	--4135
		x"08",	--4136
		x"04",	--4137
		x"09",	--4138
		x"02",	--4139
		x"0e",	--4140
		x"0f",	--4141
		x"08",	--4142
		x"09",	--4143
		x"08",	--4144
		x"09",	--4145
		x"0e",	--4146
		x"0f",	--4147
		x"3e",	--4148
		x"7f",	--4149
		x"0f",	--4150
		x"3e",	--4151
		x"40",	--4152
		x"26",	--4153
		x"38",	--4154
		x"3f",	--4155
		x"09",	--4156
		x"0e",	--4157
		x"0f",	--4158
		x"12",	--4159
		x"0f",	--4160
		x"0e",	--4161
		x"12",	--4162
		x"0f",	--4163
		x"0e",	--4164
		x"12",	--4165
		x"0f",	--4166
		x"0e",	--4167
		x"12",	--4168
		x"0f",	--4169
		x"0e",	--4170
		x"12",	--4171
		x"0f",	--4172
		x"0e",	--4173
		x"12",	--4174
		x"0f",	--4175
		x"0e",	--4176
		x"12",	--4177
		x"0f",	--4178
		x"0e",	--4179
		x"3e",	--4180
		x"3f",	--4181
		x"7f",	--4182
		x"5d",	--4183
		x"39",	--4184
		x"00",	--4185
		x"72",	--4186
		x"4d",	--4187
		x"70",	--4188
		x"08",	--4189
		x"09",	--4190
		x"da",	--4191
		x"0f",	--4192
		x"d8",	--4193
		x"0e",	--4194
		x"0f",	--4195
		x"3e",	--4196
		x"80",	--4197
		x"0f",	--4198
		x"0e",	--4199
		x"04",	--4200
		x"38",	--4201
		x"40",	--4202
		x"09",	--4203
		x"d0",	--4204
		x"0f",	--4205
		x"ce",	--4206
		x"f9",	--4207
		x"0b",	--4208
		x"0a",	--4209
		x"2a",	--4210
		x"5b",	--4211
		x"02",	--4212
		x"3b",	--4213
		x"7f",	--4214
		x"1d",	--4215
		x"02",	--4216
		x"12",	--4217
		x"0d",	--4218
		x"12",	--4219
		x"0d",	--4220
		x"12",	--4221
		x"0d",	--4222
		x"12",	--4223
		x"0d",	--4224
		x"12",	--4225
		x"0d",	--4226
		x"12",	--4227
		x"0d",	--4228
		x"12",	--4229
		x"0d",	--4230
		x"4d",	--4231
		x"5f",	--4232
		x"03",	--4233
		x"3f",	--4234
		x"80",	--4235
		x"0f",	--4236
		x"0f",	--4237
		x"ce",	--4238
		x"01",	--4239
		x"0d",	--4240
		x"2d",	--4241
		x"0a",	--4242
		x"51",	--4243
		x"be",	--4244
		x"82",	--4245
		x"02",	--4246
		x"0c",	--4247
		x"0d",	--4248
		x"0c",	--4249
		x"0d",	--4250
		x"0c",	--4251
		x"0d",	--4252
		x"0c",	--4253
		x"0d",	--4254
		x"0c",	--4255
		x"0d",	--4256
		x"0c",	--4257
		x"0d",	--4258
		x"0c",	--4259
		x"0d",	--4260
		x"0c",	--4261
		x"0d",	--4262
		x"fe",	--4263
		x"03",	--4264
		x"00",	--4265
		x"3d",	--4266
		x"00",	--4267
		x"0b",	--4268
		x"3f",	--4269
		x"81",	--4270
		x"0c",	--4271
		x"0d",	--4272
		x"0a",	--4273
		x"3f",	--4274
		x"3d",	--4275
		x"00",	--4276
		x"f9",	--4277
		x"8e",	--4278
		x"02",	--4279
		x"8e",	--4280
		x"04",	--4281
		x"8e",	--4282
		x"06",	--4283
		x"3a",	--4284
		x"3b",	--4285
		x"30",	--4286
		x"3d",	--4287
		x"ff",	--4288
		x"2a",	--4289
		x"3d",	--4290
		x"81",	--4291
		x"8e",	--4292
		x"02",	--4293
		x"fe",	--4294
		x"03",	--4295
		x"00",	--4296
		x"0c",	--4297
		x"0d",	--4298
		x"0c",	--4299
		x"0d",	--4300
		x"0c",	--4301
		x"0d",	--4302
		x"0c",	--4303
		x"0d",	--4304
		x"0c",	--4305
		x"0d",	--4306
		x"0c",	--4307
		x"0d",	--4308
		x"0c",	--4309
		x"0d",	--4310
		x"0c",	--4311
		x"0d",	--4312
		x"0a",	--4313
		x"0b",	--4314
		x"0a",	--4315
		x"3b",	--4316
		x"00",	--4317
		x"8e",	--4318
		x"04",	--4319
		x"8e",	--4320
		x"06",	--4321
		x"3a",	--4322
		x"3b",	--4323
		x"30",	--4324
		x"0b",	--4325
		x"ad",	--4326
		x"ee",	--4327
		x"00",	--4328
		x"3a",	--4329
		x"3b",	--4330
		x"30",	--4331
		x"0a",	--4332
		x"0c",	--4333
		x"0c",	--4334
		x"0d",	--4335
		x"0c",	--4336
		x"3d",	--4337
		x"10",	--4338
		x"0c",	--4339
		x"02",	--4340
		x"0d",	--4341
		x"08",	--4342
		x"de",	--4343
		x"00",	--4344
		x"e4",	--4345
		x"0b",	--4346
		x"f2",	--4347
		x"ee",	--4348
		x"00",	--4349
		x"e3",	--4350
		x"ce",	--4351
		x"00",	--4352
		x"dc",	--4353
		x"0b",	--4354
		x"6d",	--4355
		x"6d",	--4356
		x"12",	--4357
		x"6c",	--4358
		x"6c",	--4359
		x"0f",	--4360
		x"6d",	--4361
		x"41",	--4362
		x"6c",	--4363
		x"11",	--4364
		x"6d",	--4365
		x"0d",	--4366
		x"6c",	--4367
		x"14",	--4368
		x"5d",	--4369
		x"01",	--4370
		x"5d",	--4371
		x"01",	--4372
		x"14",	--4373
		x"4d",	--4374
		x"09",	--4375
		x"1e",	--4376
		x"0f",	--4377
		x"3b",	--4378
		x"30",	--4379
		x"6c",	--4380
		x"28",	--4381
		x"ce",	--4382
		x"01",	--4383
		x"f7",	--4384
		x"3e",	--4385
		x"0f",	--4386
		x"3b",	--4387
		x"30",	--4388
		x"cf",	--4389
		x"01",	--4390
		x"f0",	--4391
		x"3e",	--4392
		x"f8",	--4393
		x"1b",	--4394
		x"02",	--4395
		x"1c",	--4396
		x"02",	--4397
		x"0c",	--4398
		x"e6",	--4399
		x"0b",	--4400
		x"16",	--4401
		x"1b",	--4402
		x"04",	--4403
		x"1f",	--4404
		x"06",	--4405
		x"1c",	--4406
		x"04",	--4407
		x"1e",	--4408
		x"06",	--4409
		x"0e",	--4410
		x"da",	--4411
		x"0f",	--4412
		x"02",	--4413
		x"0c",	--4414
		x"d6",	--4415
		x"0f",	--4416
		x"06",	--4417
		x"0e",	--4418
		x"02",	--4419
		x"0b",	--4420
		x"02",	--4421
		x"0e",	--4422
		x"d1",	--4423
		x"4d",	--4424
		x"ce",	--4425
		x"3e",	--4426
		x"d6",	--4427
		x"6c",	--4428
		x"d7",	--4429
		x"5e",	--4430
		x"01",	--4431
		x"5f",	--4432
		x"01",	--4433
		x"0e",	--4434
		x"c5",	--4435
		x"1e",	--4436
		x"1e",	--4437
		x"1e",	--4438
		x"0b",	--4439
		x"1d",	--4440
		x"1c",	--4441
		x"cd",	--4442
		x"00",	--4443
		x"1d",	--4444
		x"82",	--4445
		x"1c",	--4446
		x"3e",	--4447
		x"82",	--4448
		x"1e",	--4449
		x"30",	--4450
		x"3f",	--4451
		x"30",	--4452
		x"0b",	--4453
		x"0a",	--4454
		x"21",	--4455
		x"81",	--4456
		x"00",	--4457
		x"1a",	--4458
		x"1c",	--4459
		x"1b",	--4460
		x"1e",	--4461
		x"0d",	--4462
		x"0e",	--4463
		x"3f",	--4464
		x"a8",	--4465
		x"b0",	--4466
		x"fc",	--4467
		x"0f",	--4468
		x"05",	--4469
		x"0e",	--4470
		x"0e",	--4471
		x"ce",	--4472
		x"ff",	--4473
		x"04",	--4474
		x"1e",	--4475
		x"1c",	--4476
		x"ce",	--4477
		x"00",	--4478
		x"21",	--4479
		x"3a",	--4480
		x"3b",	--4481
		x"30",	--4482
		x"92",	--4483
		x"02",	--4484
		x"1c",	--4485
		x"b2",	--4486
		x"ff",	--4487
		x"1e",	--4488
		x"0e",	--4489
		x"3e",	--4490
		x"06",	--4491
		x"1f",	--4492
		x"04",	--4493
		x"b0",	--4494
		x"ca",	--4495
		x"30",	--4496
		x"92",	--4497
		x"02",	--4498
		x"1c",	--4499
		x"92",	--4500
		x"04",	--4501
		x"1e",	--4502
		x"0e",	--4503
		x"3e",	--4504
		x"1f",	--4505
		x"06",	--4506
		x"b0",	--4507
		x"ca",	--4508
		x"30",	--4509
		x"0c",	--4510
		x"82",	--4511
		x"1c",	--4512
		x"b2",	--4513
		x"ff",	--4514
		x"1e",	--4515
		x"0e",	--4516
		x"0f",	--4517
		x"b0",	--4518
		x"ca",	--4519
		x"30",	--4520
		x"82",	--4521
		x"1c",	--4522
		x"82",	--4523
		x"1e",	--4524
		x"0e",	--4525
		x"0f",	--4526
		x"b0",	--4527
		x"ca",	--4528
		x"30",	--4529
		x"0b",	--4530
		x"0a",	--4531
		x"09",	--4532
		x"08",	--4533
		x"07",	--4534
		x"06",	--4535
		x"05",	--4536
		x"04",	--4537
		x"31",	--4538
		x"08",	--4539
		x"81",	--4540
		x"04",	--4541
		x"09",	--4542
		x"1f",	--4543
		x"1a",	--4544
		x"1d",	--4545
		x"1c",	--4546
		x"4c",	--4547
		x"04",	--4548
		x"84",	--4549
		x"45",	--4550
		x"4e",	--4551
		x"7e",	--4552
		x"40",	--4553
		x"11",	--4554
		x"f1",	--4555
		x"30",	--4556
		x"00",	--4557
		x"0e",	--4558
		x"8e",	--4559
		x"5e",	--4560
		x"03",	--4561
		x"7e",	--4562
		x"58",	--4563
		x"02",	--4564
		x"7e",	--4565
		x"78",	--4566
		x"c1",	--4567
		x"01",	--4568
		x"0c",	--4569
		x"2c",	--4570
		x"0f",	--4571
		x"7e",	--4572
		x"20",	--4573
		x"04",	--4574
		x"f1",	--4575
		x"30",	--4576
		x"00",	--4577
		x"04",	--4578
		x"4c",	--4579
		x"05",	--4580
		x"c1",	--4581
		x"00",	--4582
		x"0c",	--4583
		x"1c",	--4584
		x"01",	--4585
		x"0c",	--4586
		x"0a",	--4587
		x"8c",	--4588
		x"8c",	--4589
		x"8c",	--4590
		x"8c",	--4591
		x"0b",	--4592
		x"06",	--4593
		x"0c",	--4594
		x"8c",	--4595
		x"8c",	--4596
		x"8c",	--4597
		x"8c",	--4598
		x"07",	--4599
		x"0a",	--4600
		x"0b",	--4601
		x"0e",	--4602
		x"8e",	--4603
		x"c1",	--4604
		x"02",	--4605
		x"6e",	--4606
		x"02",	--4607
		x"07",	--4608
		x"01",	--4609
		x"37",	--4610
		x"4f",	--4611
		x"7f",	--4612
		x"10",	--4613
		x"3c",	--4614
		x"1d",	--4615
		x"04",	--4616
		x"3d",	--4617
		x"1d",	--4618
		x"cd",	--4619
		x"00",	--4620
		x"fc",	--4621
		x"1d",	--4622
		x"04",	--4623
		x"09",	--4624
		x"02",	--4625
		x"09",	--4626
		x"01",	--4627
		x"09",	--4628
		x"e1",	--4629
		x"02",	--4630
		x"05",	--4631
		x"09",	--4632
		x"02",	--4633
		x"09",	--4634
		x"01",	--4635
		x"09",	--4636
		x"05",	--4637
		x"07",	--4638
		x"01",	--4639
		x"05",	--4640
		x"4f",	--4641
		x"0d",	--4642
		x"f1",	--4643
		x"20",	--4644
		x"06",	--4645
		x"06",	--4646
		x"0b",	--4647
		x"0e",	--4648
		x"0f",	--4649
		x"0f",	--4650
		x"6f",	--4651
		x"8f",	--4652
		x"16",	--4653
		x"88",	--4654
		x"01",	--4655
		x"06",	--4656
		x"06",	--4657
		x"f6",	--4658
		x"0b",	--4659
		x"f1",	--4660
		x"30",	--4661
		x"06",	--4662
		x"05",	--4663
		x"05",	--4664
		x"5f",	--4665
		x"06",	--4666
		x"8f",	--4667
		x"88",	--4668
		x"1b",	--4669
		x"0f",	--4670
		x"0f",	--4671
		x"0f",	--4672
		x"f7",	--4673
		x"0a",	--4674
		x"06",	--4675
		x"0b",	--4676
		x"07",	--4677
		x"1b",	--4678
		x"0f",	--4679
		x"0f",	--4680
		x"6f",	--4681
		x"8f",	--4682
		x"16",	--4683
		x"88",	--4684
		x"06",	--4685
		x"f7",	--4686
		x"e1",	--4687
		x"02",	--4688
		x"02",	--4689
		x"4a",	--4690
		x"08",	--4691
		x"1a",	--4692
		x"04",	--4693
		x"0a",	--4694
		x"0d",	--4695
		x"3f",	--4696
		x"30",	--4697
		x"88",	--4698
		x"7a",	--4699
		x"4a",	--4700
		x"fa",	--4701
		x"44",	--4702
		x"0b",	--4703
		x"f3",	--4704
		x"37",	--4705
		x"8f",	--4706
		x"88",	--4707
		x"1b",	--4708
		x"0f",	--4709
		x"0f",	--4710
		x"6f",	--4711
		x"4f",	--4712
		x"07",	--4713
		x"07",	--4714
		x"f5",	--4715
		x"04",	--4716
		x"3f",	--4717
		x"20",	--4718
		x"88",	--4719
		x"1b",	--4720
		x"0b",	--4721
		x"fa",	--4722
		x"0f",	--4723
		x"31",	--4724
		x"34",	--4725
		x"35",	--4726
		x"36",	--4727
		x"37",	--4728
		x"38",	--4729
		x"39",	--4730
		x"3a",	--4731
		x"3b",	--4732
		x"30",	--4733
		x"0b",	--4734
		x"0a",	--4735
		x"09",	--4736
		x"08",	--4737
		x"07",	--4738
		x"06",	--4739
		x"05",	--4740
		x"04",	--4741
		x"31",	--4742
		x"b6",	--4743
		x"81",	--4744
		x"3a",	--4745
		x"06",	--4746
		x"05",	--4747
		x"81",	--4748
		x"3e",	--4749
		x"c1",	--4750
		x"2f",	--4751
		x"c1",	--4752
		x"2b",	--4753
		x"c1",	--4754
		x"2e",	--4755
		x"c1",	--4756
		x"2a",	--4757
		x"81",	--4758
		x"30",	--4759
		x"81",	--4760
		x"26",	--4761
		x"07",	--4762
		x"81",	--4763
		x"2c",	--4764
		x"0e",	--4765
		x"3e",	--4766
		x"1c",	--4767
		x"81",	--4768
		x"1c",	--4769
		x"30",	--4770
		x"76",	--4771
		x"0f",	--4772
		x"1f",	--4773
		x"81",	--4774
		x"40",	--4775
		x"07",	--4776
		x"1e",	--4777
		x"7e",	--4778
		x"25",	--4779
		x"13",	--4780
		x"81",	--4781
		x"00",	--4782
		x"81",	--4783
		x"02",	--4784
		x"81",	--4785
		x"3e",	--4786
		x"c1",	--4787
		x"2f",	--4788
		x"c1",	--4789
		x"2b",	--4790
		x"c1",	--4791
		x"2e",	--4792
		x"c1",	--4793
		x"2a",	--4794
		x"81",	--4795
		x"30",	--4796
		x"30",	--4797
		x"6c",	--4798
		x"05",	--4799
		x"8e",	--4800
		x"0f",	--4801
		x"91",	--4802
		x"3c",	--4803
		x"91",	--4804
		x"2c",	--4805
		x"30",	--4806
		x"52",	--4807
		x"7e",	--4808
		x"63",	--4809
		x"c5",	--4810
		x"7e",	--4811
		x"64",	--4812
		x"27",	--4813
		x"7e",	--4814
		x"30",	--4815
		x"94",	--4816
		x"7e",	--4817
		x"31",	--4818
		x"1a",	--4819
		x"7e",	--4820
		x"2a",	--4821
		x"77",	--4822
		x"7e",	--4823
		x"2b",	--4824
		x"0a",	--4825
		x"7e",	--4826
		x"23",	--4827
		x"42",	--4828
		x"7e",	--4829
		x"25",	--4830
		x"e0",	--4831
		x"7e",	--4832
		x"20",	--4833
		x"32",	--4834
		x"56",	--4835
		x"7e",	--4836
		x"2d",	--4837
		x"49",	--4838
		x"7e",	--4839
		x"2e",	--4840
		x"5b",	--4841
		x"7e",	--4842
		x"2b",	--4843
		x"28",	--4844
		x"47",	--4845
		x"7e",	--4846
		x"3a",	--4847
		x"8c",	--4848
		x"7e",	--4849
		x"58",	--4850
		x"21",	--4851
		x"e9",	--4852
		x"7e",	--4853
		x"6f",	--4854
		x"24",	--4855
		x"7e",	--4856
		x"70",	--4857
		x"0a",	--4858
		x"7e",	--4859
		x"69",	--4860
		x"e3",	--4861
		x"7e",	--4862
		x"6c",	--4863
		x"22",	--4864
		x"7e",	--4865
		x"64",	--4866
		x"11",	--4867
		x"dc",	--4868
		x"7e",	--4869
		x"73",	--4870
		x"98",	--4871
		x"7e",	--4872
		x"74",	--4873
		x"04",	--4874
		x"7e",	--4875
		x"70",	--4876
		x"07",	--4877
		x"b8",	--4878
		x"7e",	--4879
		x"75",	--4880
		x"d1",	--4881
		x"7e",	--4882
		x"78",	--4883
		x"d2",	--4884
		x"19",	--4885
		x"3e",	--4886
		x"18",	--4887
		x"2c",	--4888
		x"08",	--4889
		x"30",	--4890
		x"40",	--4891
		x"b1",	--4892
		x"28",	--4893
		x"cb",	--4894
		x"f1",	--4895
		x"00",	--4896
		x"30",	--4897
		x"70",	--4898
		x"69",	--4899
		x"59",	--4900
		x"6e",	--4901
		x"04",	--4902
		x"7e",	--4903
		x"fe",	--4904
		x"6e",	--4905
		x"01",	--4906
		x"5e",	--4907
		x"c1",	--4908
		x"00",	--4909
		x"30",	--4910
		x"70",	--4911
		x"f1",	--4912
		x"10",	--4913
		x"00",	--4914
		x"30",	--4915
		x"70",	--4916
		x"f1",	--4917
		x"2b",	--4918
		x"02",	--4919
		x"30",	--4920
		x"70",	--4921
		x"f1",	--4922
		x"2b",	--4923
		x"02",	--4924
		x"02",	--4925
		x"30",	--4926
		x"70",	--4927
		x"f1",	--4928
		x"20",	--4929
		x"02",	--4930
		x"30",	--4931
		x"70",	--4932
		x"c1",	--4933
		x"2a",	--4934
		x"02",	--4935
		x"30",	--4936
		x"56",	--4937
		x"d1",	--4938
		x"2e",	--4939
		x"30",	--4940
		x"70",	--4941
		x"0e",	--4942
		x"2e",	--4943
		x"2a",	--4944
		x"0a",	--4945
		x"03",	--4946
		x"81",	--4947
		x"26",	--4948
		x"0d",	--4949
		x"c1",	--4950
		x"2e",	--4951
		x"02",	--4952
		x"30",	--4953
		x"66",	--4954
		x"f1",	--4955
		x"10",	--4956
		x"00",	--4957
		x"3a",	--4958
		x"81",	--4959
		x"26",	--4960
		x"91",	--4961
		x"26",	--4962
		x"05",	--4963
		x"27",	--4964
		x"81",	--4965
		x"26",	--4966
		x"15",	--4967
		x"c1",	--4968
		x"2e",	--4969
		x"12",	--4970
		x"69",	--4971
		x"79",	--4972
		x"10",	--4973
		x"5e",	--4974
		x"01",	--4975
		x"4e",	--4976
		x"4e",	--4977
		x"0e",	--4978
		x"0e",	--4979
		x"4e",	--4980
		x"6a",	--4981
		x"7a",	--4982
		x"7f",	--4983
		x"4a",	--4984
		x"c1",	--4985
		x"00",	--4986
		x"30",	--4987
		x"70",	--4988
		x"1a",	--4989
		x"26",	--4990
		x"0a",	--4991
		x"0c",	--4992
		x"0c",	--4993
		x"0c",	--4994
		x"0a",	--4995
		x"81",	--4996
		x"26",	--4997
		x"b1",	--4998
		x"d0",	--4999
		x"26",	--5000
		x"8e",	--5001
		x"81",	--5002
		x"26",	--5003
		x"d1",	--5004
		x"2a",	--5005
		x"30",	--5006
		x"70",	--5007
		x"07",	--5008
		x"27",	--5009
		x"6e",	--5010
		x"c1",	--5011
		x"2e",	--5012
		x"03",	--5013
		x"c1",	--5014
		x"2a",	--5015
		x"26",	--5016
		x"c1",	--5017
		x"04",	--5018
		x"c1",	--5019
		x"05",	--5020
		x"0e",	--5021
		x"2e",	--5022
		x"03",	--5023
		x"07",	--5024
		x"27",	--5025
		x"2e",	--5026
		x"c1",	--5027
		x"2e",	--5028
		x"07",	--5029
		x"e1",	--5030
		x"01",	--5031
		x"1f",	--5032
		x"26",	--5033
		x"c1",	--5034
		x"03",	--5035
		x"06",	--5036
		x"c1",	--5037
		x"2a",	--5038
		x"03",	--5039
		x"91",	--5040
		x"26",	--5041
		x"30",	--5042
		x"0e",	--5043
		x"02",	--5044
		x"3e",	--5045
		x"7e",	--5046
		x"11",	--5047
		x"04",	--5048
		x"11",	--5049
		x"04",	--5050
		x"1d",	--5051
		x"34",	--5052
		x"1f",	--5053
		x"3e",	--5054
		x"b0",	--5055
		x"64",	--5056
		x"21",	--5057
		x"81",	--5058
		x"2c",	--5059
		x"05",	--5060
		x"30",	--5061
		x"52",	--5062
		x"07",	--5063
		x"27",	--5064
		x"29",	--5065
		x"81",	--5066
		x"1e",	--5067
		x"5e",	--5068
		x"09",	--5069
		x"01",	--5070
		x"4e",	--5071
		x"4e",	--5072
		x"4e",	--5073
		x"4e",	--5074
		x"6a",	--5075
		x"7a",	--5076
		x"f7",	--5077
		x"4a",	--5078
		x"c1",	--5079
		x"00",	--5080
		x"05",	--5081
		x"b1",	--5082
		x"10",	--5083
		x"28",	--5084
		x"53",	--5085
		x"d1",	--5086
		x"01",	--5087
		x"06",	--5088
		x"e1",	--5089
		x"00",	--5090
		x"b1",	--5091
		x"0a",	--5092
		x"28",	--5093
		x"03",	--5094
		x"b1",	--5095
		x"10",	--5096
		x"28",	--5097
		x"6b",	--5098
		x"6b",	--5099
		x"24",	--5100
		x"0c",	--5101
		x"3c",	--5102
		x"28",	--5103
		x"17",	--5104
		x"02",	--5105
		x"16",	--5106
		x"04",	--5107
		x"1b",	--5108
		x"06",	--5109
		x"81",	--5110
		x"1e",	--5111
		x"81",	--5112
		x"20",	--5113
		x"81",	--5114
		x"22",	--5115
		x"81",	--5116
		x"24",	--5117
		x"d1",	--5118
		x"2b",	--5119
		x"08",	--5120
		x"06",	--5121
		x"07",	--5122
		x"04",	--5123
		x"06",	--5124
		x"02",	--5125
		x"0b",	--5126
		x"02",	--5127
		x"c1",	--5128
		x"2b",	--5129
		x"0b",	--5130
		x"0b",	--5131
		x"0b",	--5132
		x"c1",	--5133
		x"2f",	--5134
		x"05",	--5135
		x"20",	--5136
		x"5b",	--5137
		x"07",	--5138
		x"0d",	--5139
		x"27",	--5140
		x"28",	--5141
		x"1b",	--5142
		x"02",	--5143
		x"81",	--5144
		x"1e",	--5145
		x"81",	--5146
		x"20",	--5147
		x"d1",	--5148
		x"2b",	--5149
		x"08",	--5150
		x"09",	--5151
		x"06",	--5152
		x"27",	--5153
		x"2b",	--5154
		x"81",	--5155
		x"1e",	--5156
		x"d1",	--5157
		x"2b",	--5158
		x"0b",	--5159
		x"02",	--5160
		x"c1",	--5161
		x"2b",	--5162
		x"0b",	--5163
		x"0b",	--5164
		x"0b",	--5165
		x"c1",	--5166
		x"2f",	--5167
		x"05",	--5168
		x"f1",	--5169
		x"00",	--5170
		x"12",	--5171
		x"c1",	--5172
		x"2b",	--5173
		x"0f",	--5174
		x"68",	--5175
		x"b1",	--5176
		x"10",	--5177
		x"28",	--5178
		x"03",	--5179
		x"78",	--5180
		x"40",	--5181
		x"05",	--5182
		x"b1",	--5183
		x"28",	--5184
		x"04",	--5185
		x"78",	--5186
		x"20",	--5187
		x"c1",	--5188
		x"00",	--5189
		x"68",	--5190
		x"68",	--5191
		x"30",	--5192
		x"c1",	--5193
		x"2f",	--5194
		x"2d",	--5195
		x"f1",	--5196
		x"2d",	--5197
		x"02",	--5198
		x"68",	--5199
		x"11",	--5200
		x"b1",	--5201
		x"1e",	--5202
		x"b1",	--5203
		x"20",	--5204
		x"b1",	--5205
		x"22",	--5206
		x"b1",	--5207
		x"24",	--5208
		x"91",	--5209
		x"1e",	--5210
		x"81",	--5211
		x"20",	--5212
		x"81",	--5213
		x"22",	--5214
		x"81",	--5215
		x"24",	--5216
		x"17",	--5217
		x"58",	--5218
		x"0f",	--5219
		x"1a",	--5220
		x"1e",	--5221
		x"1b",	--5222
		x"20",	--5223
		x"3a",	--5224
		x"3b",	--5225
		x"0e",	--5226
		x"0f",	--5227
		x"1e",	--5228
		x"0f",	--5229
		x"81",	--5230
		x"1e",	--5231
		x"81",	--5232
		x"20",	--5233
		x"06",	--5234
		x"1a",	--5235
		x"1e",	--5236
		x"3a",	--5237
		x"1a",	--5238
		x"81",	--5239
		x"1e",	--5240
		x"c1",	--5241
		x"1b",	--5242
		x"68",	--5243
		x"6a",	--5244
		x"16",	--5245
		x"1e",	--5246
		x"91",	--5247
		x"20",	--5248
		x"3c",	--5249
		x"18",	--5250
		x"22",	--5251
		x"14",	--5252
		x"24",	--5253
		x"07",	--5254
		x"37",	--5255
		x"1a",	--5256
		x"09",	--5257
		x"91",	--5258
		x"28",	--5259
		x"32",	--5260
		x"1b",	--5261
		x"28",	--5262
		x"8b",	--5263
		x"8b",	--5264
		x"8b",	--5265
		x"8b",	--5266
		x"81",	--5267
		x"34",	--5268
		x"81",	--5269
		x"36",	--5270
		x"81",	--5271
		x"38",	--5272
		x"11",	--5273
		x"3a",	--5274
		x"11",	--5275
		x"3a",	--5276
		x"11",	--5277
		x"3a",	--5278
		x"11",	--5279
		x"3a",	--5280
		x"0c",	--5281
		x"1d",	--5282
		x"44",	--5283
		x"0e",	--5284
		x"0f",	--5285
		x"b0",	--5286
		x"06",	--5287
		x"31",	--5288
		x"0b",	--5289
		x"3c",	--5290
		x"0a",	--5291
		x"05",	--5292
		x"7b",	--5293
		x"30",	--5294
		x"c7",	--5295
		x"00",	--5296
		x"0c",	--5297
		x"4b",	--5298
		x"d1",	--5299
		x"01",	--5300
		x"03",	--5301
		x"7a",	--5302
		x"37",	--5303
		x"02",	--5304
		x"7a",	--5305
		x"57",	--5306
		x"4a",	--5307
		x"c7",	--5308
		x"00",	--5309
		x"06",	--5310
		x"36",	--5311
		x"11",	--5312
		x"3a",	--5313
		x"11",	--5314
		x"3a",	--5315
		x"11",	--5316
		x"3a",	--5317
		x"11",	--5318
		x"3a",	--5319
		x"0c",	--5320
		x"1d",	--5321
		x"44",	--5322
		x"0e",	--5323
		x"0f",	--5324
		x"b0",	--5325
		x"e0",	--5326
		x"31",	--5327
		x"09",	--5328
		x"81",	--5329
		x"3c",	--5330
		x"08",	--5331
		x"04",	--5332
		x"37",	--5333
		x"0c",	--5334
		x"b2",	--5335
		x"0d",	--5336
		x"b0",	--5337
		x"0e",	--5338
		x"ae",	--5339
		x"0f",	--5340
		x"ac",	--5341
		x"81",	--5342
		x"1e",	--5343
		x"81",	--5344
		x"20",	--5345
		x"81",	--5346
		x"22",	--5347
		x"81",	--5348
		x"24",	--5349
		x"6c",	--5350
		x"58",	--5351
		x"3e",	--5352
		x"14",	--5353
		x"1e",	--5354
		x"17",	--5355
		x"20",	--5356
		x"08",	--5357
		x"38",	--5358
		x"1a",	--5359
		x"19",	--5360
		x"28",	--5361
		x"89",	--5362
		x"89",	--5363
		x"89",	--5364
		x"89",	--5365
		x"1c",	--5366
		x"28",	--5367
		x"0d",	--5368
		x"0e",	--5369
		x"0f",	--5370
		x"b0",	--5371
		x"0a",	--5372
		x"0b",	--5373
		x"3e",	--5374
		x"0a",	--5375
		x"05",	--5376
		x"7b",	--5377
		x"30",	--5378
		x"c8",	--5379
		x"00",	--5380
		x"0c",	--5381
		x"4b",	--5382
		x"d1",	--5383
		x"01",	--5384
		x"03",	--5385
		x"7a",	--5386
		x"37",	--5387
		x"02",	--5388
		x"7a",	--5389
		x"57",	--5390
		x"4a",	--5391
		x"c8",	--5392
		x"00",	--5393
		x"06",	--5394
		x"36",	--5395
		x"1c",	--5396
		x"28",	--5397
		x"0d",	--5398
		x"0e",	--5399
		x"0f",	--5400
		x"b0",	--5401
		x"d4",	--5402
		x"04",	--5403
		x"07",	--5404
		x"38",	--5405
		x"0e",	--5406
		x"d0",	--5407
		x"0f",	--5408
		x"ce",	--5409
		x"81",	--5410
		x"1e",	--5411
		x"81",	--5412
		x"20",	--5413
		x"2c",	--5414
		x"17",	--5415
		x"1e",	--5416
		x"08",	--5417
		x"38",	--5418
		x"1a",	--5419
		x"1e",	--5420
		x"28",	--5421
		x"0f",	--5422
		x"b0",	--5423
		x"7a",	--5424
		x"0d",	--5425
		x"3f",	--5426
		x"0a",	--5427
		x"05",	--5428
		x"7d",	--5429
		x"30",	--5430
		x"c8",	--5431
		x"00",	--5432
		x"0c",	--5433
		x"4d",	--5434
		x"d1",	--5435
		x"01",	--5436
		x"03",	--5437
		x"7c",	--5438
		x"37",	--5439
		x"02",	--5440
		x"7c",	--5441
		x"57",	--5442
		x"4c",	--5443
		x"c8",	--5444
		x"00",	--5445
		x"06",	--5446
		x"36",	--5447
		x"1e",	--5448
		x"28",	--5449
		x"0f",	--5450
		x"b0",	--5451
		x"60",	--5452
		x"07",	--5453
		x"38",	--5454
		x"0f",	--5455
		x"db",	--5456
		x"81",	--5457
		x"1e",	--5458
		x"b1",	--5459
		x"0a",	--5460
		x"28",	--5461
		x"02",	--5462
		x"c1",	--5463
		x"02",	--5464
		x"c1",	--5465
		x"2e",	--5466
		x"2a",	--5467
		x"0f",	--5468
		x"3f",	--5469
		x"1c",	--5470
		x"81",	--5471
		x"42",	--5472
		x"1a",	--5473
		x"1c",	--5474
		x"8a",	--5475
		x"8a",	--5476
		x"8a",	--5477
		x"8a",	--5478
		x"81",	--5479
		x"44",	--5480
		x"81",	--5481
		x"46",	--5482
		x"0a",	--5483
		x"8a",	--5484
		x"8a",	--5485
		x"8a",	--5486
		x"8a",	--5487
		x"81",	--5488
		x"48",	--5489
		x"1c",	--5490
		x"42",	--5491
		x"1d",	--5492
		x"44",	--5493
		x"1c",	--5494
		x"46",	--5495
		x"1d",	--5496
		x"48",	--5497
		x"2c",	--5498
		x"1c",	--5499
		x"26",	--5500
		x"0e",	--5501
		x"e1",	--5502
		x"01",	--5503
		x"5e",	--5504
		x"26",	--5505
		x"4e",	--5506
		x"c1",	--5507
		x"03",	--5508
		x"06",	--5509
		x"c1",	--5510
		x"2a",	--5511
		x"03",	--5512
		x"91",	--5513
		x"26",	--5514
		x"30",	--5515
		x"11",	--5516
		x"04",	--5517
		x"11",	--5518
		x"04",	--5519
		x"1d",	--5520
		x"34",	--5521
		x"0e",	--5522
		x"1e",	--5523
		x"1f",	--5524
		x"3e",	--5525
		x"b0",	--5526
		x"64",	--5527
		x"21",	--5528
		x"81",	--5529
		x"2c",	--5530
		x"0d",	--5531
		x"7f",	--5532
		x"8f",	--5533
		x"91",	--5534
		x"3c",	--5535
		x"0e",	--5536
		x"0e",	--5537
		x"19",	--5538
		x"40",	--5539
		x"f7",	--5540
		x"81",	--5541
		x"3e",	--5542
		x"81",	--5543
		x"2c",	--5544
		x"07",	--5545
		x"0e",	--5546
		x"91",	--5547
		x"26",	--5548
		x"30",	--5549
		x"d1",	--5550
		x"2e",	--5551
		x"c1",	--5552
		x"2a",	--5553
		x"03",	--5554
		x"05",	--5555
		x"d1",	--5556
		x"2a",	--5557
		x"81",	--5558
		x"26",	--5559
		x"17",	--5560
		x"16",	--5561
		x"40",	--5562
		x"6e",	--5563
		x"4e",	--5564
		x"02",	--5565
		x"30",	--5566
		x"48",	--5567
		x"1f",	--5568
		x"2c",	--5569
		x"31",	--5570
		x"4a",	--5571
		x"34",	--5572
		x"35",	--5573
		x"36",	--5574
		x"37",	--5575
		x"38",	--5576
		x"39",	--5577
		x"3a",	--5578
		x"3b",	--5579
		x"30",	--5580
		x"0d",	--5581
		x"0f",	--5582
		x"04",	--5583
		x"3d",	--5584
		x"03",	--5585
		x"3f",	--5586
		x"1f",	--5587
		x"0e",	--5588
		x"03",	--5589
		x"5d",	--5590
		x"3e",	--5591
		x"1e",	--5592
		x"0d",	--5593
		x"b0",	--5594
		x"60",	--5595
		x"3d",	--5596
		x"6d",	--5597
		x"02",	--5598
		x"3e",	--5599
		x"1e",	--5600
		x"5d",	--5601
		x"02",	--5602
		x"3f",	--5603
		x"1f",	--5604
		x"30",	--5605
		x"b0",	--5606
		x"9a",	--5607
		x"0f",	--5608
		x"30",	--5609
		x"0b",	--5610
		x"0a",	--5611
		x"09",	--5612
		x"79",	--5613
		x"20",	--5614
		x"0a",	--5615
		x"0b",	--5616
		x"0c",	--5617
		x"0d",	--5618
		x"0e",	--5619
		x"0f",	--5620
		x"0c",	--5621
		x"0d",	--5622
		x"0d",	--5623
		x"06",	--5624
		x"02",	--5625
		x"0c",	--5626
		x"03",	--5627
		x"0c",	--5628
		x"0d",	--5629
		x"1e",	--5630
		x"19",	--5631
		x"f2",	--5632
		x"39",	--5633
		x"3a",	--5634
		x"3b",	--5635
		x"30",	--5636
		x"b0",	--5637
		x"d4",	--5638
		x"0e",	--5639
		x"0f",	--5640
		x"30",	--5641
		x"0b",	--5642
		x"0b",	--5643
		x"0f",	--5644
		x"06",	--5645
		x"3b",	--5646
		x"03",	--5647
		x"3e",	--5648
		x"3f",	--5649
		x"1e",	--5650
		x"0f",	--5651
		x"0d",	--5652
		x"05",	--5653
		x"5b",	--5654
		x"3c",	--5655
		x"3d",	--5656
		x"1c",	--5657
		x"0d",	--5658
		x"b0",	--5659
		x"d4",	--5660
		x"6b",	--5661
		x"04",	--5662
		x"3c",	--5663
		x"3d",	--5664
		x"1c",	--5665
		x"0d",	--5666
		x"5b",	--5667
		x"04",	--5668
		x"3e",	--5669
		x"3f",	--5670
		x"1e",	--5671
		x"0f",	--5672
		x"3b",	--5673
		x"30",	--5674
		x"b0",	--5675
		x"14",	--5676
		x"0e",	--5677
		x"0f",	--5678
		x"30",	--5679
		x"7c",	--5680
		x"10",	--5681
		x"0d",	--5682
		x"0e",	--5683
		x"0f",	--5684
		x"0e",	--5685
		x"0e",	--5686
		x"02",	--5687
		x"0e",	--5688
		x"1f",	--5689
		x"1c",	--5690
		x"f8",	--5691
		x"30",	--5692
		x"b0",	--5693
		x"60",	--5694
		x"0f",	--5695
		x"30",	--5696
		x"07",	--5697
		x"06",	--5698
		x"05",	--5699
		x"04",	--5700
		x"30",	--5701
		x"40",	--5702
		x"04",	--5703
		x"05",	--5704
		x"06",	--5705
		x"07",	--5706
		x"08",	--5707
		x"09",	--5708
		x"0a",	--5709
		x"0b",	--5710
		x"0c",	--5711
		x"0d",	--5712
		x"0e",	--5713
		x"0f",	--5714
		x"08",	--5715
		x"09",	--5716
		x"0a",	--5717
		x"0b",	--5718
		x"0b",	--5719
		x"0e",	--5720
		x"08",	--5721
		x"0a",	--5722
		x"0b",	--5723
		x"05",	--5724
		x"09",	--5725
		x"08",	--5726
		x"02",	--5727
		x"08",	--5728
		x"05",	--5729
		x"08",	--5730
		x"09",	--5731
		x"0a",	--5732
		x"0b",	--5733
		x"1c",	--5734
		x"91",	--5735
		x"00",	--5736
		x"e5",	--5737
		x"21",	--5738
		x"34",	--5739
		x"35",	--5740
		x"36",	--5741
		x"37",	--5742
		x"30",	--5743
		x"0b",	--5744
		x"0a",	--5745
		x"09",	--5746
		x"08",	--5747
		x"18",	--5748
		x"0a",	--5749
		x"19",	--5750
		x"0c",	--5751
		x"1a",	--5752
		x"0e",	--5753
		x"1b",	--5754
		x"10",	--5755
		x"b0",	--5756
		x"82",	--5757
		x"38",	--5758
		x"39",	--5759
		x"3a",	--5760
		x"3b",	--5761
		x"30",	--5762
		x"0b",	--5763
		x"0a",	--5764
		x"09",	--5765
		x"08",	--5766
		x"18",	--5767
		x"0a",	--5768
		x"19",	--5769
		x"0c",	--5770
		x"1a",	--5771
		x"0e",	--5772
		x"1b",	--5773
		x"10",	--5774
		x"b0",	--5775
		x"82",	--5776
		x"0c",	--5777
		x"0d",	--5778
		x"0e",	--5779
		x"0f",	--5780
		x"38",	--5781
		x"39",	--5782
		x"3a",	--5783
		x"3b",	--5784
		x"30",	--5785
		x"0b",	--5786
		x"0a",	--5787
		x"09",	--5788
		x"08",	--5789
		x"07",	--5790
		x"18",	--5791
		x"0c",	--5792
		x"19",	--5793
		x"0e",	--5794
		x"1a",	--5795
		x"10",	--5796
		x"1b",	--5797
		x"12",	--5798
		x"b0",	--5799
		x"82",	--5800
		x"17",	--5801
		x"14",	--5802
		x"87",	--5803
		x"00",	--5804
		x"87",	--5805
		x"02",	--5806
		x"87",	--5807
		x"04",	--5808
		x"87",	--5809
		x"06",	--5810
		x"37",	--5811
		x"38",	--5812
		x"39",	--5813
		x"3a",	--5814
		x"3b",	--5815
		x"30",	--5816
		x"00",	--5817
		x"32",	--5818
		x"f0",	--5819
		x"fd",	--5820
		x"53",	--5821
		x"6f",	--5822
		x"0d",	--5823
		x"00",	--5824
		x"6f",	--5825
		x"72",	--5826
		x"63",	--5827
		x"20",	--5828
		x"73",	--5829
		x"67",	--5830
		x"3a",	--5831
		x"0a",	--5832
		x"09",	--5833
		x"63",	--5834
		x"4c",	--5835
		x"46",	--5836
		x"20",	--5837
		x"49",	--5838
		x"48",	--5839
		x"20",	--5840
		x"54",	--5841
		x"4d",	--5842
		x"4f",	--5843
		x"54",	--5844
		x"0d",	--5845
		x"00",	--5846
		x"64",	--5847
		x"25",	--5848
		x"0d",	--5849
		x"00",	--5850
		x"6f",	--5851
		x"20",	--5852
		x"6d",	--5853
		x"6c",	--5854
		x"6d",	--5855
		x"6e",	--5856
		x"65",	--5857
		x"20",	--5858
		x"65",	--5859
		x"0d",	--5860
		x"00",	--5861
		x"61",	--5862
		x"74",	--5863
		x"6e",	--5864
		x"20",	--5865
		x"6f",	--5866
		x"20",	--5867
		x"20",	--5868
		x"65",	--5869
		x"20",	--5870
		x"62",	--5871
		x"6e",	--5872
		x"66",	--5873
		x"6c",	--5874
		x"0d",	--5875
		x"00",	--5876
		x"65",	--5877
		x"73",	--5878
		x"6f",	--5879
		x"6c",	--5880
		x"20",	--5881
		x"6f",	--5882
		x"20",	--5883
		x"65",	--5884
		x"20",	--5885
		x"68",	--5886
		x"74",	--5887
		x"0a",	--5888
		x"53",	--5889
		x"6f",	--5890
		x"0d",	--5891
		x"00",	--5892
		x"72",	--5893
		x"6f",	--5894
		x"3a",	--5895
		x"6d",	--5896
		x"73",	--5897
		x"69",	--5898
		x"67",	--5899
		x"61",	--5900
		x"67",	--5901
		x"6d",	--5902
		x"6e",	--5903
		x"0d",	--5904
		x"00",	--5905
		x"6f",	--5906
		x"72",	--5907
		x"63",	--5908
		x"20",	--5909
		x"73",	--5910
		x"67",	--5911
		x"3a",	--5912
		x"0a",	--5913
		x"09",	--5914
		x"73",	--5915
		x"4c",	--5916
		x"46",	--5917
		x"20",	--5918
		x"49",	--5919
		x"48",	--5920
		x"20",	--5921
		x"54",	--5922
		x"4d",	--5923
		x"4f",	--5924
		x"54",	--5925
		x"0d",	--5926
		x"00",	--5927
		x"64",	--5928
		x"25",	--5929
		x"0d",	--5930
		x"00",	--5931
		x"6c",	--5932
		x"20",	--5933
		x"6c",	--5934
		x"00",	--5935
		x"73",	--5936
		x"0a",	--5937
		x"25",	--5938
		x"20",	--5939
		x"64",	--5940
		x"0a",	--5941
		x"5c",	--5942
		x"84",	--5943
		x"8a",	--5944
		x"92",	--5945
		x"9a",	--5946
		x"a2",	--5947
		x"74",	--5948
		x"7c",	--5949
		x"0d",	--5950
		x"3d",	--5951
		x"3d",	--5952
		x"3d",	--5953
		x"20",	--5954
		x"61",	--5955
		x"63",	--5956
		x"6c",	--5957
		x"4d",	--5958
		x"55",	--5959
		x"3d",	--5960
		x"3d",	--5961
		x"3d",	--5962
		x"0d",	--5963
		x"00",	--5964
		x"6e",	--5965
		x"65",	--5966
		x"61",	--5967
		x"74",	--5968
		x"76",	--5969
		x"20",	--5970
		x"6f",	--5971
		x"65",	--5972
		x"77",	--5973
		x"69",	--5974
		x"65",	--5975
		x"72",	--5976
		x"61",	--5977
		x"00",	--5978
		x"75",	--5979
		x"7a",	--5980
		x"72",	--5981
		x"70",	--5982
		x"6d",	--5983
		x"65",	--5984
		x"63",	--5985
		x"64",	--5986
		x"72",	--5987
		x"73",	--5988
		x"65",	--5989
		x"64",	--5990
		x"63",	--5991
		x"6e",	--5992
		x"72",	--5993
		x"6c",	--5994
		x"65",	--5995
		x"00",	--5996
		x"70",	--5997
		x"65",	--5998
		x"20",	--5999
		x"6f",	--6000
		x"66",	--6001
		x"67",	--6002
		x"72",	--6003
		x"74",	--6004
		x"6f",	--6005
		x"00",	--6006
		x"6f",	--6007
		x"74",	--6008
		x"6f",	--6009
		x"64",	--6010
		x"72",	--6011
		x"0d",	--6012
		x"00",	--6013
		x"20",	--6014
		x"00",	--6015
		x"63",	--6016
		x"55",	--6017
		x"0d",	--6018
		x"00",	--6019
		x"4f",	--6020
		x"4e",	--6021
		x"0a",	--6022
		x"52",	--6023
		x"47",	--6024
		x"54",	--6025
		x"0a",	--6026
		x"4c",	--6027
		x"46",	--6028
		x"0d",	--6029
		x"00",	--6030
		x"77",	--6031
		x"69",	--6032
		x"65",	--6033
		x"0d",	--6034
		x"65",	--6035
		x"72",	--6036
		x"72",	--6037
		x"20",	--6038
		x"69",	--6039
		x"73",	--6040
		x"6e",	--6041
		x"20",	--6042
		x"72",	--6043
		x"75",	--6044
		x"65",	--6045
		x"74",	--6046
		x"0a",	--6047
		x"63",	--6048
		x"72",	--6049
		x"65",	--6050
		x"74",	--6051
		x"75",	--6052
		x"61",	--6053
		x"65",	--6054
		x"0d",	--6055
		x"00",	--6056
		x"25",	--6057
		x"20",	--6058
		x"45",	--6059
		x"49",	--6060
		x"54",	--6061
		x"52",	--6062
		x"56",	--6063
		x"4c",	--6064
		x"45",	--6065
		x"0a",	--6066
		x"72",	--6067
		x"25",	--6068
		x"20",	--6069
		x"3d",	--6070
		x"64",	--6071
		x"0a",	--6072
		x"09",	--6073
		x"73",	--6074
		x"52",	--6075
		x"47",	--6076
		x"53",	--6077
		x"45",	--6078
		x"0d",	--6079
		x"00",	--6080
		x"65",	--6081
		x"64",	--6082
		x"0d",	--6083
		x"25",	--6084
		x"20",	--6085
		x"73",	--6086
		x"6e",	--6087
		x"74",	--6088
		x"61",	--6089
		x"6e",	--6090
		x"6d",	--6091
		x"65",	--6092
		x"0d",	--6093
		x"00",	--6094
		x"63",	--6095
		x"25",	--6096
		x"0d",	--6097
		x"00",	--6098
		x"63",	--6099
		x"20",	--6100
		x"6f",	--6101
		x"73",	--6102
		x"63",	--6103
		x"20",	--6104
		x"6f",	--6105
		x"6d",	--6106
		x"6e",	--6107
		x"0d",	--6108
		x"00",	--6109
		x"e2",	--6110
		x"10",	--6111
		x"10",	--6112
		x"10",	--6113
		x"10",	--6114
		x"10",	--6115
		x"10",	--6116
		x"10",	--6117
		x"10",	--6118
		x"10",	--6119
		x"10",	--6120
		x"10",	--6121
		x"10",	--6122
		x"10",	--6123
		x"10",	--6124
		x"10",	--6125
		x"10",	--6126
		x"10",	--6127
		x"10",	--6128
		x"10",	--6129
		x"10",	--6130
		x"10",	--6131
		x"10",	--6132
		x"10",	--6133
		x"10",	--6134
		x"10",	--6135
		x"10",	--6136
		x"10",	--6137
		x"10",	--6138
		x"d4",	--6139
		x"10",	--6140
		x"10",	--6141
		x"10",	--6142
		x"10",	--6143
		x"10",	--6144
		x"10",	--6145
		x"10",	--6146
		x"10",	--6147
		x"10",	--6148
		x"10",	--6149
		x"10",	--6150
		x"10",	--6151
		x"10",	--6152
		x"10",	--6153
		x"10",	--6154
		x"10",	--6155
		x"10",	--6156
		x"10",	--6157
		x"10",	--6158
		x"10",	--6159
		x"10",	--6160
		x"10",	--6161
		x"10",	--6162
		x"10",	--6163
		x"10",	--6164
		x"10",	--6165
		x"10",	--6166
		x"10",	--6167
		x"10",	--6168
		x"10",	--6169
		x"10",	--6170
		x"c6",	--6171
		x"b8",	--6172
		x"aa",	--6173
		x"10",	--6174
		x"10",	--6175
		x"10",	--6176
		x"10",	--6177
		x"10",	--6178
		x"10",	--6179
		x"10",	--6180
		x"92",	--6181
		x"10",	--6182
		x"80",	--6183
		x"10",	--6184
		x"10",	--6185
		x"10",	--6186
		x"10",	--6187
		x"64",	--6188
		x"10",	--6189
		x"10",	--6190
		x"10",	--6191
		x"56",	--6192
		x"44",	--6193
		x"30",	--6194
		x"32",	--6195
		x"34",	--6196
		x"36",	--6197
		x"38",	--6198
		x"61",	--6199
		x"63",	--6200
		x"65",	--6201
		x"00",	--6202
		x"00",	--6203
		x"00",	--6204
		x"00",	--6205
		x"00",	--6206
		x"00",	--6207
		x"02",	--6208
		x"03",	--6209
		x"03",	--6210
		x"04",	--6211
		x"04",	--6212
		x"04",	--6213
		x"04",	--6214
		x"05",	--6215
		x"05",	--6216
		x"05",	--6217
		x"05",	--6218
		x"05",	--6219
		x"05",	--6220
		x"05",	--6221
		x"05",	--6222
		x"06",	--6223
		x"06",	--6224
		x"06",	--6225
		x"06",	--6226
		x"06",	--6227
		x"06",	--6228
		x"06",	--6229
		x"06",	--6230
		x"06",	--6231
		x"06",	--6232
		x"06",	--6233
		x"06",	--6234
		x"06",	--6235
		x"06",	--6236
		x"06",	--6237
		x"06",	--6238
		x"07",	--6239
		x"07",	--6240
		x"07",	--6241
		x"07",	--6242
		x"07",	--6243
		x"07",	--6244
		x"07",	--6245
		x"07",	--6246
		x"07",	--6247
		x"07",	--6248
		x"07",	--6249
		x"07",	--6250
		x"07",	--6251
		x"07",	--6252
		x"07",	--6253
		x"07",	--6254
		x"07",	--6255
		x"07",	--6256
		x"07",	--6257
		x"07",	--6258
		x"07",	--6259
		x"07",	--6260
		x"07",	--6261
		x"07",	--6262
		x"07",	--6263
		x"07",	--6264
		x"07",	--6265
		x"07",	--6266
		x"07",	--6267
		x"07",	--6268
		x"07",	--6269
		x"07",	--6270
		x"08",	--6271
		x"08",	--6272
		x"08",	--6273
		x"08",	--6274
		x"08",	--6275
		x"08",	--6276
		x"08",	--6277
		x"08",	--6278
		x"08",	--6279
		x"08",	--6280
		x"08",	--6281
		x"08",	--6282
		x"08",	--6283
		x"08",	--6284
		x"08",	--6285
		x"08",	--6286
		x"08",	--6287
		x"08",	--6288
		x"08",	--6289
		x"08",	--6290
		x"08",	--6291
		x"08",	--6292
		x"08",	--6293
		x"08",	--6294
		x"08",	--6295
		x"08",	--6296
		x"08",	--6297
		x"08",	--6298
		x"08",	--6299
		x"08",	--6300
		x"08",	--6301
		x"08",	--6302
		x"08",	--6303
		x"08",	--6304
		x"08",	--6305
		x"08",	--6306
		x"08",	--6307
		x"08",	--6308
		x"08",	--6309
		x"08",	--6310
		x"08",	--6311
		x"08",	--6312
		x"08",	--6313
		x"08",	--6314
		x"08",	--6315
		x"08",	--6316
		x"08",	--6317
		x"08",	--6318
		x"08",	--6319
		x"08",	--6320
		x"08",	--6321
		x"08",	--6322
		x"08",	--6323
		x"08",	--6324
		x"08",	--6325
		x"08",	--6326
		x"08",	--6327
		x"08",	--6328
		x"08",	--6329
		x"08",	--6330
		x"08",	--6331
		x"08",	--6332
		x"08",	--6333
		x"08",	--6334
		x"28",	--6335
		x"75",	--6336
		x"6c",	--6337
		x"00",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"68",	--6342
		x"6c",	--6343
		x"00",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"48",	--8176
		x"48",	--8177
		x"48",	--8178
		x"48",	--8179
		x"48",	--8180
		x"48",	--8181
		x"48",	--8182
		x"ec",	--8183
		x"3e",	--8184
		x"48",	--8185
		x"48",	--8186
		x"48",	--8187
		x"48",	--8188
		x"48",	--8189
		x"48",	--8190
		x"00");	--8191
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"f1",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"d4",	--44
		x"12",	--45
		x"ce",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"ee",	--50
		x"12",	--51
		x"d2",	--52
		x"53",	--53
		x"40",	--54
		x"ee",	--55
		x"40",	--56
		x"c9",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"ce",	--61
		x"40",	--62
		x"ee",	--63
		x"40",	--64
		x"cb",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"ce",	--69
		x"40",	--70
		x"ee",	--71
		x"40",	--72
		x"cb",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"ce",	--77
		x"40",	--78
		x"ee",	--79
		x"40",	--80
		x"c3",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"ce",	--85
		x"40",	--86
		x"ee",	--87
		x"40",	--88
		x"c6",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"ce",	--93
		x"40",	--94
		x"ee",	--95
		x"40",	--96
		x"c8",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"ce",	--101
		x"40",	--102
		x"ee",	--103
		x"40",	--104
		x"c3",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"ce",	--109
		x"40",	--110
		x"ee",	--111
		x"40",	--112
		x"c5",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"ce",	--117
		x"40",	--118
		x"ee",	--119
		x"40",	--120
		x"c5",	--121
		x"40",	--122
		x"00",	--123
		x"12",	--124
		x"ce",	--125
		x"43",	--126
		x"43",	--127
		x"12",	--128
		x"ce",	--129
		x"43",	--130
		x"40",	--131
		x"4e",	--132
		x"40",	--133
		x"01",	--134
		x"41",	--135
		x"50",	--136
		x"00",	--137
		x"12",	--138
		x"cd",	--139
		x"41",	--140
		x"50",	--141
		x"00",	--142
		x"12",	--143
		x"cd",	--144
		x"43",	--145
		x"40",	--146
		x"4e",	--147
		x"40",	--148
		x"01",	--149
		x"41",	--150
		x"50",	--151
		x"00",	--152
		x"12",	--153
		x"cd",	--154
		x"41",	--155
		x"50",	--156
		x"00",	--157
		x"12",	--158
		x"cd",	--159
		x"41",	--160
		x"50",	--161
		x"00",	--162
		x"41",	--163
		x"50",	--164
		x"00",	--165
		x"12",	--166
		x"c6",	--167
		x"40",	--168
		x"01",	--169
		x"41",	--170
		x"52",	--171
		x"12",	--172
		x"d0",	--173
		x"40",	--174
		x"01",	--175
		x"41",	--176
		x"53",	--177
		x"12",	--178
		x"d0",	--179
		x"41",	--180
		x"53",	--181
		x"41",	--182
		x"52",	--183
		x"12",	--184
		x"c8",	--185
		x"41",	--186
		x"50",	--187
		x"00",	--188
		x"41",	--189
		x"50",	--190
		x"00",	--191
		x"12",	--192
		x"c8",	--193
		x"12",	--194
		x"cf",	--195
		x"40",	--196
		x"01",	--197
		x"41",	--198
		x"12",	--199
		x"d0",	--200
		x"41",	--201
		x"12",	--202
		x"c3",	--203
		x"40",	--204
		x"00",	--205
		x"40",	--206
		x"11",	--207
		x"41",	--208
		x"12",	--209
		x"d1",	--210
		x"12",	--211
		x"41",	--212
		x"12",	--213
		x"12",	--214
		x"12",	--215
		x"12",	--216
		x"39",	--217
		x"12",	--218
		x"b7",	--219
		x"12",	--220
		x"3a",	--221
		x"12",	--222
		x"49",	--223
		x"40",	--224
		x"00",	--225
		x"41",	--226
		x"50",	--227
		x"00",	--228
		x"41",	--229
		x"50",	--230
		x"00",	--231
		x"41",	--232
		x"50",	--233
		x"00",	--234
		x"12",	--235
		x"c5",	--236
		x"50",	--237
		x"00",	--238
		x"12",	--239
		x"41",	--240
		x"12",	--241
		x"12",	--242
		x"12",	--243
		x"12",	--244
		x"39",	--245
		x"12",	--246
		x"b7",	--247
		x"12",	--248
		x"3a",	--249
		x"12",	--250
		x"49",	--251
		x"40",	--252
		x"00",	--253
		x"41",	--254
		x"50",	--255
		x"00",	--256
		x"41",	--257
		x"50",	--258
		x"00",	--259
		x"41",	--260
		x"50",	--261
		x"00",	--262
		x"12",	--263
		x"c5",	--264
		x"50",	--265
		x"00",	--266
		x"41",	--267
		x"50",	--268
		x"00",	--269
		x"41",	--270
		x"50",	--271
		x"00",	--272
		x"12",	--273
		x"c3",	--274
		x"12",	--275
		x"c3",	--276
		x"40",	--277
		x"ff",	--278
		x"00",	--279
		x"d2",	--280
		x"43",	--281
		x"43",	--282
		x"3c",	--283
		x"43",	--284
		x"3c",	--285
		x"43",	--286
		x"3c",	--287
		x"43",	--288
		x"12",	--289
		x"d4",	--290
		x"93",	--291
		x"27",	--292
		x"12",	--293
		x"d4",	--294
		x"93",	--295
		x"20",	--296
		x"90",	--297
		x"00",	--298
		x"24",	--299
		x"90",	--300
		x"00",	--301
		x"27",	--302
		x"92",	--303
		x"20",	--304
		x"3c",	--305
		x"12",	--306
		x"ee",	--307
		x"12",	--308
		x"d2",	--309
		x"53",	--310
		x"40",	--311
		x"00",	--312
		x"51",	--313
		x"5f",	--314
		x"43",	--315
		x"00",	--316
		x"4f",	--317
		x"41",	--318
		x"00",	--319
		x"12",	--320
		x"cf",	--321
		x"43",	--322
		x"3f",	--323
		x"93",	--324
		x"27",	--325
		x"53",	--326
		x"12",	--327
		x"ee",	--328
		x"12",	--329
		x"d2",	--330
		x"53",	--331
		x"3f",	--332
		x"90",	--333
		x"00",	--334
		x"2f",	--335
		x"93",	--336
		x"02",	--337
		x"24",	--338
		x"4f",	--339
		x"11",	--340
		x"12",	--341
		x"12",	--342
		x"ee",	--343
		x"4f",	--344
		x"00",	--345
		x"12",	--346
		x"d2",	--347
		x"52",	--348
		x"41",	--349
		x"00",	--350
		x"40",	--351
		x"00",	--352
		x"51",	--353
		x"5a",	--354
		x"4f",	--355
		x"00",	--356
		x"53",	--357
		x"3f",	--358
		x"93",	--359
		x"20",	--360
		x"90",	--361
		x"00",	--362
		x"23",	--363
		x"3f",	--364
		x"93",	--365
		x"23",	--366
		x"90",	--367
		x"00",	--368
		x"24",	--369
		x"90",	--370
		x"00",	--371
		x"34",	--372
		x"90",	--373
		x"00",	--374
		x"23",	--375
		x"3c",	--376
		x"90",	--377
		x"00",	--378
		x"24",	--379
		x"90",	--380
		x"00",	--381
		x"23",	--382
		x"3c",	--383
		x"12",	--384
		x"ef",	--385
		x"12",	--386
		x"d2",	--387
		x"53",	--388
		x"12",	--389
		x"c4",	--390
		x"43",	--391
		x"3f",	--392
		x"12",	--393
		x"ef",	--394
		x"12",	--395
		x"d2",	--396
		x"53",	--397
		x"12",	--398
		x"c4",	--399
		x"43",	--400
		x"3f",	--401
		x"12",	--402
		x"ef",	--403
		x"12",	--404
		x"d2",	--405
		x"53",	--406
		x"12",	--407
		x"c4",	--408
		x"43",	--409
		x"3f",	--410
		x"12",	--411
		x"ef",	--412
		x"12",	--413
		x"d2",	--414
		x"53",	--415
		x"12",	--416
		x"c4",	--417
		x"43",	--418
		x"3f",	--419
		x"40",	--420
		x"ed",	--421
		x"4f",	--422
		x"02",	--423
		x"41",	--424
		x"12",	--425
		x"12",	--426
		x"82",	--427
		x"4f",	--428
		x"4e",	--429
		x"93",	--430
		x"38",	--431
		x"41",	--432
		x"4b",	--433
		x"00",	--434
		x"12",	--435
		x"cc",	--436
		x"4f",	--437
		x"93",	--438
		x"24",	--439
		x"41",	--440
		x"4b",	--441
		x"00",	--442
		x"4d",	--443
		x"00",	--444
		x"12",	--445
		x"cc",	--446
		x"4f",	--447
		x"41",	--448
		x"00",	--449
		x"42",	--450
		x"02",	--451
		x"12",	--452
		x"d1",	--453
		x"43",	--454
		x"52",	--455
		x"41",	--456
		x"41",	--457
		x"41",	--458
		x"40",	--459
		x"00",	--460
		x"40",	--461
		x"11",	--462
		x"3f",	--463
		x"40",	--464
		x"11",	--465
		x"3f",	--466
		x"43",	--467
		x"42",	--468
		x"02",	--469
		x"12",	--470
		x"c6",	--471
		x"43",	--472
		x"42",	--473
		x"02",	--474
		x"12",	--475
		x"c6",	--476
		x"12",	--477
		x"ed",	--478
		x"12",	--479
		x"d2",	--480
		x"53",	--481
		x"41",	--482
		x"93",	--483
		x"02",	--484
		x"24",	--485
		x"42",	--486
		x"02",	--487
		x"12",	--488
		x"c6",	--489
		x"42",	--490
		x"02",	--491
		x"12",	--492
		x"c6",	--493
		x"41",	--494
		x"43",	--495
		x"40",	--496
		x"c3",	--497
		x"12",	--498
		x"cf",	--499
		x"4f",	--500
		x"02",	--501
		x"3f",	--502
		x"4f",	--503
		x"02",	--504
		x"4e",	--505
		x"02",	--506
		x"41",	--507
		x"12",	--508
		x"12",	--509
		x"83",	--510
		x"4e",	--511
		x"90",	--512
		x"00",	--513
		x"38",	--514
		x"20",	--515
		x"41",	--516
		x"4b",	--517
		x"00",	--518
		x"12",	--519
		x"cd",	--520
		x"4f",	--521
		x"41",	--522
		x"4b",	--523
		x"00",	--524
		x"12",	--525
		x"cd",	--526
		x"4f",	--527
		x"12",	--528
		x"12",	--529
		x"12",	--530
		x"ed",	--531
		x"12",	--532
		x"d2",	--533
		x"50",	--534
		x"00",	--535
		x"4a",	--536
		x"42",	--537
		x"02",	--538
		x"12",	--539
		x"c6",	--540
		x"4b",	--541
		x"42",	--542
		x"02",	--543
		x"12",	--544
		x"c6",	--545
		x"43",	--546
		x"53",	--547
		x"41",	--548
		x"41",	--549
		x"41",	--550
		x"41",	--551
		x"4b",	--552
		x"00",	--553
		x"12",	--554
		x"cc",	--555
		x"43",	--556
		x"4f",	--557
		x"42",	--558
		x"02",	--559
		x"12",	--560
		x"d0",	--561
		x"3f",	--562
		x"12",	--563
		x"ed",	--564
		x"12",	--565
		x"d2",	--566
		x"4b",	--567
		x"00",	--568
		x"12",	--569
		x"ed",	--570
		x"12",	--571
		x"d2",	--572
		x"52",	--573
		x"43",	--574
		x"3f",	--575
		x"40",	--576
		x"ff",	--577
		x"42",	--578
		x"02",	--579
		x"12",	--580
		x"c6",	--581
		x"40",	--582
		x"00",	--583
		x"42",	--584
		x"02",	--585
		x"12",	--586
		x"c6",	--587
		x"43",	--588
		x"40",	--589
		x"00",	--590
		x"42",	--591
		x"02",	--592
		x"12",	--593
		x"d0",	--594
		x"41",	--595
		x"40",	--596
		x"00",	--597
		x"42",	--598
		x"02",	--599
		x"12",	--600
		x"c6",	--601
		x"40",	--602
		x"ff",	--603
		x"42",	--604
		x"02",	--605
		x"12",	--606
		x"c6",	--607
		x"43",	--608
		x"40",	--609
		x"00",	--610
		x"42",	--611
		x"02",	--612
		x"12",	--613
		x"d0",	--614
		x"41",	--615
		x"40",	--616
		x"ff",	--617
		x"42",	--618
		x"02",	--619
		x"12",	--620
		x"c6",	--621
		x"40",	--622
		x"ff",	--623
		x"42",	--624
		x"02",	--625
		x"12",	--626
		x"c6",	--627
		x"43",	--628
		x"40",	--629
		x"00",	--630
		x"42",	--631
		x"02",	--632
		x"12",	--633
		x"d0",	--634
		x"41",	--635
		x"40",	--636
		x"00",	--637
		x"42",	--638
		x"02",	--639
		x"12",	--640
		x"c6",	--641
		x"40",	--642
		x"00",	--643
		x"42",	--644
		x"02",	--645
		x"12",	--646
		x"c6",	--647
		x"43",	--648
		x"40",	--649
		x"00",	--650
		x"42",	--651
		x"02",	--652
		x"12",	--653
		x"d0",	--654
		x"41",	--655
		x"12",	--656
		x"ed",	--657
		x"12",	--658
		x"d2",	--659
		x"53",	--660
		x"43",	--661
		x"41",	--662
		x"40",	--663
		x"c0",	--664
		x"01",	--665
		x"40",	--666
		x"00",	--667
		x"01",	--668
		x"40",	--669
		x"02",	--670
		x"01",	--671
		x"12",	--672
		x"ed",	--673
		x"12",	--674
		x"d2",	--675
		x"43",	--676
		x"01",	--677
		x"40",	--678
		x"ed",	--679
		x"00",	--680
		x"12",	--681
		x"d2",	--682
		x"53",	--683
		x"43",	--684
		x"41",	--685
		x"12",	--686
		x"12",	--687
		x"12",	--688
		x"4f",	--689
		x"4f",	--690
		x"00",	--691
		x"12",	--692
		x"d0",	--693
		x"4e",	--694
		x"4f",	--695
		x"89",	--696
		x"00",	--697
		x"79",	--698
		x"00",	--699
		x"12",	--700
		x"dc",	--701
		x"4a",	--702
		x"00",	--703
		x"4b",	--704
		x"00",	--705
		x"4e",	--706
		x"4f",	--707
		x"49",	--708
		x"12",	--709
		x"ca",	--710
		x"43",	--711
		x"40",	--712
		x"3f",	--713
		x"12",	--714
		x"d7",	--715
		x"4e",	--716
		x"4f",	--717
		x"40",	--718
		x"66",	--719
		x"40",	--720
		x"3f",	--721
		x"12",	--722
		x"db",	--723
		x"93",	--724
		x"24",	--725
		x"34",	--726
		x"40",	--727
		x"cc",	--728
		x"40",	--729
		x"3d",	--730
		x"4a",	--731
		x"4b",	--732
		x"12",	--733
		x"dc",	--734
		x"93",	--735
		x"34",	--736
		x"40",	--737
		x"cc",	--738
		x"40",	--739
		x"3d",	--740
		x"4a",	--741
		x"4b",	--742
		x"49",	--743
		x"00",	--744
		x"12",	--745
		x"ce",	--746
		x"41",	--747
		x"41",	--748
		x"41",	--749
		x"41",	--750
		x"40",	--751
		x"66",	--752
		x"40",	--753
		x"3f",	--754
		x"3f",	--755
		x"12",	--756
		x"12",	--757
		x"4f",	--758
		x"4c",	--759
		x"4e",	--760
		x"00",	--761
		x"4d",	--762
		x"00",	--763
		x"12",	--764
		x"00",	--765
		x"12",	--766
		x"00",	--767
		x"12",	--768
		x"00",	--769
		x"12",	--770
		x"00",	--771
		x"12",	--772
		x"00",	--773
		x"12",	--774
		x"00",	--775
		x"41",	--776
		x"00",	--777
		x"41",	--778
		x"00",	--779
		x"12",	--780
		x"c9",	--781
		x"50",	--782
		x"00",	--783
		x"4a",	--784
		x"00",	--785
		x"4b",	--786
		x"40",	--787
		x"c5",	--788
		x"12",	--789
		x"cf",	--790
		x"4f",	--791
		x"00",	--792
		x"41",	--793
		x"41",	--794
		x"41",	--795
		x"12",	--796
		x"4f",	--797
		x"4f",	--798
		x"00",	--799
		x"12",	--800
		x"d0",	--801
		x"4e",	--802
		x"00",	--803
		x"4f",	--804
		x"00",	--805
		x"43",	--806
		x"4b",	--807
		x"00",	--808
		x"4b",	--809
		x"00",	--810
		x"12",	--811
		x"d0",	--812
		x"41",	--813
		x"41",	--814
		x"12",	--815
		x"4f",	--816
		x"43",	--817
		x"40",	--818
		x"3f",	--819
		x"4f",	--820
		x"00",	--821
		x"12",	--822
		x"ce",	--823
		x"4b",	--824
		x"00",	--825
		x"12",	--826
		x"d0",	--827
		x"41",	--828
		x"41",	--829
		x"12",	--830
		x"4f",	--831
		x"4e",	--832
		x"10",	--833
		x"11",	--834
		x"10",	--835
		x"11",	--836
		x"4d",	--837
		x"12",	--838
		x"dc",	--839
		x"4e",	--840
		x"4f",	--841
		x"4b",	--842
		x"12",	--843
		x"ca",	--844
		x"41",	--845
		x"41",	--846
		x"12",	--847
		x"12",	--848
		x"43",	--849
		x"40",	--850
		x"3f",	--851
		x"4a",	--852
		x"4b",	--853
		x"42",	--854
		x"02",	--855
		x"12",	--856
		x"ce",	--857
		x"4a",	--858
		x"4b",	--859
		x"42",	--860
		x"02",	--861
		x"12",	--862
		x"ce",	--863
		x"12",	--864
		x"ee",	--865
		x"12",	--866
		x"d2",	--867
		x"53",	--868
		x"41",	--869
		x"41",	--870
		x"41",	--871
		x"4f",	--872
		x"02",	--873
		x"4e",	--874
		x"02",	--875
		x"41",	--876
		x"12",	--877
		x"12",	--878
		x"83",	--879
		x"4f",	--880
		x"4e",	--881
		x"93",	--882
		x"02",	--883
		x"24",	--884
		x"90",	--885
		x"00",	--886
		x"38",	--887
		x"20",	--888
		x"41",	--889
		x"4b",	--890
		x"00",	--891
		x"12",	--892
		x"cc",	--893
		x"4f",	--894
		x"41",	--895
		x"4b",	--896
		x"00",	--897
		x"12",	--898
		x"cc",	--899
		x"4f",	--900
		x"12",	--901
		x"12",	--902
		x"12",	--903
		x"ee",	--904
		x"12",	--905
		x"d2",	--906
		x"50",	--907
		x"00",	--908
		x"4a",	--909
		x"43",	--910
		x"12",	--911
		x"dd",	--912
		x"43",	--913
		x"40",	--914
		x"42",	--915
		x"12",	--916
		x"da",	--917
		x"4e",	--918
		x"4f",	--919
		x"43",	--920
		x"40",	--921
		x"3f",	--922
		x"12",	--923
		x"d7",	--924
		x"4e",	--925
		x"4f",	--926
		x"42",	--927
		x"02",	--928
		x"12",	--929
		x"ce",	--930
		x"4b",	--931
		x"43",	--932
		x"12",	--933
		x"dd",	--934
		x"43",	--935
		x"40",	--936
		x"42",	--937
		x"12",	--938
		x"da",	--939
		x"4e",	--940
		x"4f",	--941
		x"42",	--942
		x"02",	--943
		x"12",	--944
		x"ce",	--945
		x"43",	--946
		x"53",	--947
		x"41",	--948
		x"41",	--949
		x"41",	--950
		x"41",	--951
		x"4b",	--952
		x"00",	--953
		x"12",	--954
		x"cc",	--955
		x"43",	--956
		x"4f",	--957
		x"42",	--958
		x"02",	--959
		x"12",	--960
		x"d0",	--961
		x"3f",	--962
		x"43",	--963
		x"40",	--964
		x"c6",	--965
		x"12",	--966
		x"cf",	--967
		x"4f",	--968
		x"02",	--969
		x"3f",	--970
		x"12",	--971
		x"ee",	--972
		x"12",	--973
		x"d2",	--974
		x"40",	--975
		x"ee",	--976
		x"00",	--977
		x"12",	--978
		x"d2",	--979
		x"4b",	--980
		x"00",	--981
		x"12",	--982
		x"ee",	--983
		x"12",	--984
		x"d2",	--985
		x"52",	--986
		x"43",	--987
		x"3f",	--988
		x"12",	--989
		x"12",	--990
		x"42",	--991
		x"02",	--992
		x"12",	--993
		x"d0",	--994
		x"4e",	--995
		x"4f",	--996
		x"42",	--997
		x"02",	--998
		x"12",	--999
		x"d0",	--1000
		x"12",	--1001
		x"12",	--1002
		x"e3",	--1003
		x"e3",	--1004
		x"53",	--1005
		x"63",	--1006
		x"12",	--1007
		x"12",	--1008
		x"12",	--1009
		x"ee",	--1010
		x"12",	--1011
		x"02",	--1012
		x"12",	--1013
		x"e3",	--1014
		x"50",	--1015
		x"00",	--1016
		x"12",	--1017
		x"02",	--1018
		x"12",	--1019
		x"ee",	--1020
		x"12",	--1021
		x"d2",	--1022
		x"52",	--1023
		x"41",	--1024
		x"41",	--1025
		x"41",	--1026
		x"4f",	--1027
		x"02",	--1028
		x"4e",	--1029
		x"02",	--1030
		x"41",	--1031
		x"4f",	--1032
		x"02",	--1033
		x"4e",	--1034
		x"02",	--1035
		x"41",	--1036
		x"12",	--1037
		x"12",	--1038
		x"12",	--1039
		x"12",	--1040
		x"83",	--1041
		x"4f",	--1042
		x"4e",	--1043
		x"43",	--1044
		x"00",	--1045
		x"93",	--1046
		x"24",	--1047
		x"93",	--1048
		x"02",	--1049
		x"24",	--1050
		x"43",	--1051
		x"02",	--1052
		x"41",	--1053
		x"4b",	--1054
		x"00",	--1055
		x"12",	--1056
		x"cc",	--1057
		x"4f",	--1058
		x"90",	--1059
		x"00",	--1060
		x"34",	--1061
		x"43",	--1062
		x"49",	--1063
		x"48",	--1064
		x"42",	--1065
		x"02",	--1066
		x"12",	--1067
		x"d0",	--1068
		x"43",	--1069
		x"53",	--1070
		x"41",	--1071
		x"41",	--1072
		x"41",	--1073
		x"41",	--1074
		x"41",	--1075
		x"93",	--1076
		x"02",	--1077
		x"24",	--1078
		x"43",	--1079
		x"02",	--1080
		x"42",	--1081
		x"02",	--1082
		x"12",	--1083
		x"d0",	--1084
		x"43",	--1085
		x"53",	--1086
		x"41",	--1087
		x"41",	--1088
		x"41",	--1089
		x"41",	--1090
		x"41",	--1091
		x"41",	--1092
		x"4b",	--1093
		x"00",	--1094
		x"12",	--1095
		x"cc",	--1096
		x"4f",	--1097
		x"90",	--1098
		x"00",	--1099
		x"3b",	--1100
		x"41",	--1101
		x"4b",	--1102
		x"00",	--1103
		x"12",	--1104
		x"cc",	--1105
		x"4f",	--1106
		x"41",	--1107
		x"4b",	--1108
		x"00",	--1109
		x"12",	--1110
		x"cc",	--1111
		x"4f",	--1112
		x"12",	--1113
		x"12",	--1114
		x"12",	--1115
		x"ee",	--1116
		x"12",	--1117
		x"d2",	--1118
		x"50",	--1119
		x"00",	--1120
		x"4a",	--1121
		x"43",	--1122
		x"12",	--1123
		x"dd",	--1124
		x"43",	--1125
		x"40",	--1126
		x"42",	--1127
		x"12",	--1128
		x"da",	--1129
		x"4e",	--1130
		x"4f",	--1131
		x"42",	--1132
		x"02",	--1133
		x"12",	--1134
		x"ce",	--1135
		x"4b",	--1136
		x"43",	--1137
		x"12",	--1138
		x"dd",	--1139
		x"43",	--1140
		x"40",	--1141
		x"42",	--1142
		x"12",	--1143
		x"da",	--1144
		x"4e",	--1145
		x"4f",	--1146
		x"42",	--1147
		x"02",	--1148
		x"12",	--1149
		x"ce",	--1150
		x"3f",	--1151
		x"43",	--1152
		x"12",	--1153
		x"c7",	--1154
		x"43",	--1155
		x"53",	--1156
		x"41",	--1157
		x"41",	--1158
		x"41",	--1159
		x"41",	--1160
		x"41",	--1161
		x"43",	--1162
		x"40",	--1163
		x"c7",	--1164
		x"12",	--1165
		x"cf",	--1166
		x"4f",	--1167
		x"02",	--1168
		x"3f",	--1169
		x"43",	--1170
		x"93",	--1171
		x"02",	--1172
		x"24",	--1173
		x"43",	--1174
		x"4f",	--1175
		x"02",	--1176
		x"43",	--1177
		x"41",	--1178
		x"42",	--1179
		x"00",	--1180
		x"4e",	--1181
		x"be",	--1182
		x"20",	--1183
		x"df",	--1184
		x"00",	--1185
		x"41",	--1186
		x"cf",	--1187
		x"00",	--1188
		x"41",	--1189
		x"42",	--1190
		x"02",	--1191
		x"92",	--1192
		x"2c",	--1193
		x"4e",	--1194
		x"5f",	--1195
		x"4f",	--1196
		x"ee",	--1197
		x"43",	--1198
		x"00",	--1199
		x"90",	--1200
		x"00",	--1201
		x"38",	--1202
		x"43",	--1203
		x"02",	--1204
		x"41",	--1205
		x"53",	--1206
		x"4e",	--1207
		x"02",	--1208
		x"41",	--1209
		x"40",	--1210
		x"00",	--1211
		x"00",	--1212
		x"3f",	--1213
		x"40",	--1214
		x"00",	--1215
		x"00",	--1216
		x"3f",	--1217
		x"42",	--1218
		x"00",	--1219
		x"3f",	--1220
		x"40",	--1221
		x"00",	--1222
		x"00",	--1223
		x"3f",	--1224
		x"40",	--1225
		x"00",	--1226
		x"00",	--1227
		x"3f",	--1228
		x"40",	--1229
		x"00",	--1230
		x"00",	--1231
		x"3f",	--1232
		x"40",	--1233
		x"00",	--1234
		x"00",	--1235
		x"3f",	--1236
		x"4d",	--1237
		x"00",	--1238
		x"4e",	--1239
		x"00",	--1240
		x"41",	--1241
		x"00",	--1242
		x"00",	--1243
		x"41",	--1244
		x"00",	--1245
		x"00",	--1246
		x"41",	--1247
		x"00",	--1248
		x"00",	--1249
		x"41",	--1250
		x"00",	--1251
		x"00",	--1252
		x"41",	--1253
		x"00",	--1254
		x"00",	--1255
		x"41",	--1256
		x"00",	--1257
		x"00",	--1258
		x"43",	--1259
		x"00",	--1260
		x"43",	--1261
		x"00",	--1262
		x"43",	--1263
		x"00",	--1264
		x"43",	--1265
		x"00",	--1266
		x"43",	--1267
		x"00",	--1268
		x"43",	--1269
		x"00",	--1270
		x"43",	--1271
		x"00",	--1272
		x"43",	--1273
		x"00",	--1274
		x"41",	--1275
		x"43",	--1276
		x"00",	--1277
		x"43",	--1278
		x"00",	--1279
		x"43",	--1280
		x"00",	--1281
		x"43",	--1282
		x"00",	--1283
		x"43",	--1284
		x"00",	--1285
		x"43",	--1286
		x"00",	--1287
		x"41",	--1288
		x"4d",	--1289
		x"00",	--1290
		x"4e",	--1291
		x"00",	--1292
		x"41",	--1293
		x"4d",	--1294
		x"00",	--1295
		x"4e",	--1296
		x"00",	--1297
		x"41",	--1298
		x"4d",	--1299
		x"00",	--1300
		x"4e",	--1301
		x"00",	--1302
		x"41",	--1303
		x"4d",	--1304
		x"00",	--1305
		x"4e",	--1306
		x"00",	--1307
		x"41",	--1308
		x"4d",	--1309
		x"00",	--1310
		x"4e",	--1311
		x"00",	--1312
		x"41",	--1313
		x"12",	--1314
		x"12",	--1315
		x"12",	--1316
		x"12",	--1317
		x"12",	--1318
		x"12",	--1319
		x"12",	--1320
		x"4f",	--1321
		x"4d",	--1322
		x"4e",	--1323
		x"4f",	--1324
		x"00",	--1325
		x"4f",	--1326
		x"00",	--1327
		x"4f",	--1328
		x"00",	--1329
		x"4f",	--1330
		x"00",	--1331
		x"4a",	--1332
		x"4b",	--1333
		x"46",	--1334
		x"47",	--1335
		x"12",	--1336
		x"dc",	--1337
		x"49",	--1338
		x"00",	--1339
		x"49",	--1340
		x"00",	--1341
		x"93",	--1342
		x"34",	--1343
		x"46",	--1344
		x"47",	--1345
		x"12",	--1346
		x"d7",	--1347
		x"4e",	--1348
		x"4f",	--1349
		x"4e",	--1350
		x"00",	--1351
		x"4f",	--1352
		x"00",	--1353
		x"4e",	--1354
		x"4f",	--1355
		x"4a",	--1356
		x"4b",	--1357
		x"12",	--1358
		x"dc",	--1359
		x"93",	--1360
		x"34",	--1361
		x"4a",	--1362
		x"00",	--1363
		x"4b",	--1364
		x"00",	--1365
		x"44",	--1366
		x"45",	--1367
		x"4a",	--1368
		x"4b",	--1369
		x"12",	--1370
		x"d7",	--1371
		x"4e",	--1372
		x"4f",	--1373
		x"49",	--1374
		x"00",	--1375
		x"49",	--1376
		x"00",	--1377
		x"12",	--1378
		x"d7",	--1379
		x"4e",	--1380
		x"4f",	--1381
		x"4e",	--1382
		x"00",	--1383
		x"4f",	--1384
		x"00",	--1385
		x"49",	--1386
		x"49",	--1387
		x"00",	--1388
		x"4a",	--1389
		x"4b",	--1390
		x"12",	--1391
		x"d8",	--1392
		x"4e",	--1393
		x"4f",	--1394
		x"49",	--1395
		x"00",	--1396
		x"49",	--1397
		x"00",	--1398
		x"46",	--1399
		x"47",	--1400
		x"12",	--1401
		x"d8",	--1402
		x"44",	--1403
		x"45",	--1404
		x"12",	--1405
		x"d7",	--1406
		x"4e",	--1407
		x"4f",	--1408
		x"49",	--1409
		x"00",	--1410
		x"49",	--1411
		x"00",	--1412
		x"4a",	--1413
		x"4b",	--1414
		x"12",	--1415
		x"d7",	--1416
		x"49",	--1417
		x"00",	--1418
		x"49",	--1419
		x"00",	--1420
		x"12",	--1421
		x"d8",	--1422
		x"46",	--1423
		x"47",	--1424
		x"12",	--1425
		x"d7",	--1426
		x"41",	--1427
		x"41",	--1428
		x"41",	--1429
		x"41",	--1430
		x"41",	--1431
		x"41",	--1432
		x"41",	--1433
		x"41",	--1434
		x"46",	--1435
		x"47",	--1436
		x"12",	--1437
		x"d7",	--1438
		x"4e",	--1439
		x"4f",	--1440
		x"4e",	--1441
		x"00",	--1442
		x"4f",	--1443
		x"00",	--1444
		x"4e",	--1445
		x"4f",	--1446
		x"4a",	--1447
		x"4b",	--1448
		x"12",	--1449
		x"db",	--1450
		x"93",	--1451
		x"24",	--1452
		x"37",	--1453
		x"46",	--1454
		x"47",	--1455
		x"3f",	--1456
		x"12",	--1457
		x"12",	--1458
		x"83",	--1459
		x"4f",	--1460
		x"4e",	--1461
		x"12",	--1462
		x"ef",	--1463
		x"12",	--1464
		x"d2",	--1465
		x"53",	--1466
		x"90",	--1467
		x"00",	--1468
		x"38",	--1469
		x"41",	--1470
		x"4b",	--1471
		x"00",	--1472
		x"12",	--1473
		x"cc",	--1474
		x"4f",	--1475
		x"41",	--1476
		x"4b",	--1477
		x"00",	--1478
		x"12",	--1479
		x"cc",	--1480
		x"4f",	--1481
		x"12",	--1482
		x"12",	--1483
		x"12",	--1484
		x"ef",	--1485
		x"12",	--1486
		x"d2",	--1487
		x"50",	--1488
		x"00",	--1489
		x"4b",	--1490
		x"00",	--1491
		x"43",	--1492
		x"53",	--1493
		x"41",	--1494
		x"41",	--1495
		x"41",	--1496
		x"12",	--1497
		x"ef",	--1498
		x"12",	--1499
		x"d2",	--1500
		x"40",	--1501
		x"ef",	--1502
		x"00",	--1503
		x"12",	--1504
		x"d2",	--1505
		x"4b",	--1506
		x"00",	--1507
		x"12",	--1508
		x"ef",	--1509
		x"12",	--1510
		x"d2",	--1511
		x"52",	--1512
		x"43",	--1513
		x"3f",	--1514
		x"12",	--1515
		x"83",	--1516
		x"4e",	--1517
		x"93",	--1518
		x"24",	--1519
		x"38",	--1520
		x"12",	--1521
		x"ef",	--1522
		x"12",	--1523
		x"d2",	--1524
		x"53",	--1525
		x"41",	--1526
		x"4b",	--1527
		x"00",	--1528
		x"12",	--1529
		x"cc",	--1530
		x"12",	--1531
		x"12",	--1532
		x"12",	--1533
		x"ef",	--1534
		x"12",	--1535
		x"d2",	--1536
		x"50",	--1537
		x"00",	--1538
		x"43",	--1539
		x"53",	--1540
		x"41",	--1541
		x"41",	--1542
		x"12",	--1543
		x"ef",	--1544
		x"12",	--1545
		x"d2",	--1546
		x"40",	--1547
		x"ef",	--1548
		x"00",	--1549
		x"12",	--1550
		x"d2",	--1551
		x"4b",	--1552
		x"00",	--1553
		x"12",	--1554
		x"ef",	--1555
		x"12",	--1556
		x"d2",	--1557
		x"52",	--1558
		x"43",	--1559
		x"3f",	--1560
		x"12",	--1561
		x"12",	--1562
		x"43",	--1563
		x"00",	--1564
		x"4f",	--1565
		x"93",	--1566
		x"24",	--1567
		x"53",	--1568
		x"43",	--1569
		x"43",	--1570
		x"3c",	--1571
		x"90",	--1572
		x"00",	--1573
		x"2c",	--1574
		x"5c",	--1575
		x"5c",	--1576
		x"5c",	--1577
		x"5c",	--1578
		x"11",	--1579
		x"5d",	--1580
		x"50",	--1581
		x"ff",	--1582
		x"43",	--1583
		x"4f",	--1584
		x"93",	--1585
		x"24",	--1586
		x"90",	--1587
		x"00",	--1588
		x"24",	--1589
		x"4d",	--1590
		x"50",	--1591
		x"ff",	--1592
		x"93",	--1593
		x"23",	--1594
		x"90",	--1595
		x"00",	--1596
		x"2c",	--1597
		x"5c",	--1598
		x"4c",	--1599
		x"5b",	--1600
		x"5b",	--1601
		x"5b",	--1602
		x"11",	--1603
		x"5d",	--1604
		x"50",	--1605
		x"ff",	--1606
		x"4f",	--1607
		x"93",	--1608
		x"23",	--1609
		x"43",	--1610
		x"00",	--1611
		x"4c",	--1612
		x"41",	--1613
		x"41",	--1614
		x"41",	--1615
		x"43",	--1616
		x"3f",	--1617
		x"4d",	--1618
		x"50",	--1619
		x"ff",	--1620
		x"90",	--1621
		x"00",	--1622
		x"2c",	--1623
		x"5c",	--1624
		x"5c",	--1625
		x"5c",	--1626
		x"5c",	--1627
		x"11",	--1628
		x"5d",	--1629
		x"50",	--1630
		x"ff",	--1631
		x"43",	--1632
		x"3f",	--1633
		x"4d",	--1634
		x"50",	--1635
		x"ff",	--1636
		x"90",	--1637
		x"00",	--1638
		x"2c",	--1639
		x"5c",	--1640
		x"5c",	--1641
		x"5c",	--1642
		x"5c",	--1643
		x"11",	--1644
		x"5d",	--1645
		x"50",	--1646
		x"ff",	--1647
		x"43",	--1648
		x"3f",	--1649
		x"11",	--1650
		x"12",	--1651
		x"12",	--1652
		x"ef",	--1653
		x"12",	--1654
		x"d2",	--1655
		x"52",	--1656
		x"43",	--1657
		x"4c",	--1658
		x"41",	--1659
		x"41",	--1660
		x"41",	--1661
		x"43",	--1662
		x"3f",	--1663
		x"12",	--1664
		x"12",	--1665
		x"43",	--1666
		x"00",	--1667
		x"4f",	--1668
		x"93",	--1669
		x"24",	--1670
		x"53",	--1671
		x"43",	--1672
		x"43",	--1673
		x"3c",	--1674
		x"4b",	--1675
		x"50",	--1676
		x"ff",	--1677
		x"90",	--1678
		x"00",	--1679
		x"2c",	--1680
		x"5c",	--1681
		x"4c",	--1682
		x"5d",	--1683
		x"5d",	--1684
		x"5d",	--1685
		x"11",	--1686
		x"5b",	--1687
		x"50",	--1688
		x"ff",	--1689
		x"4f",	--1690
		x"93",	--1691
		x"24",	--1692
		x"90",	--1693
		x"00",	--1694
		x"23",	--1695
		x"43",	--1696
		x"4f",	--1697
		x"93",	--1698
		x"23",	--1699
		x"12",	--1700
		x"c2",	--1701
		x"43",	--1702
		x"4a",	--1703
		x"01",	--1704
		x"4c",	--1705
		x"01",	--1706
		x"42",	--1707
		x"01",	--1708
		x"41",	--1709
		x"43",	--1710
		x"00",	--1711
		x"41",	--1712
		x"41",	--1713
		x"41",	--1714
		x"11",	--1715
		x"12",	--1716
		x"12",	--1717
		x"ef",	--1718
		x"12",	--1719
		x"d2",	--1720
		x"52",	--1721
		x"43",	--1722
		x"41",	--1723
		x"41",	--1724
		x"41",	--1725
		x"43",	--1726
		x"3f",	--1727
		x"12",	--1728
		x"12",	--1729
		x"4e",	--1730
		x"4c",	--1731
		x"4e",	--1732
		x"00",	--1733
		x"4d",	--1734
		x"00",	--1735
		x"4c",	--1736
		x"00",	--1737
		x"4d",	--1738
		x"43",	--1739
		x"40",	--1740
		x"36",	--1741
		x"40",	--1742
		x"01",	--1743
		x"12",	--1744
		x"ec",	--1745
		x"4e",	--1746
		x"00",	--1747
		x"12",	--1748
		x"c2",	--1749
		x"43",	--1750
		x"4a",	--1751
		x"01",	--1752
		x"40",	--1753
		x"00",	--1754
		x"01",	--1755
		x"42",	--1756
		x"01",	--1757
		x"00",	--1758
		x"41",	--1759
		x"43",	--1760
		x"41",	--1761
		x"41",	--1762
		x"41",	--1763
		x"12",	--1764
		x"12",	--1765
		x"12",	--1766
		x"43",	--1767
		x"00",	--1768
		x"40",	--1769
		x"3f",	--1770
		x"00",	--1771
		x"4f",	--1772
		x"4b",	--1773
		x"00",	--1774
		x"43",	--1775
		x"12",	--1776
		x"dd",	--1777
		x"43",	--1778
		x"40",	--1779
		x"3f",	--1780
		x"12",	--1781
		x"d8",	--1782
		x"4e",	--1783
		x"4f",	--1784
		x"4b",	--1785
		x"00",	--1786
		x"43",	--1787
		x"12",	--1788
		x"dd",	--1789
		x"4e",	--1790
		x"4f",	--1791
		x"48",	--1792
		x"49",	--1793
		x"12",	--1794
		x"d7",	--1795
		x"12",	--1796
		x"d4",	--1797
		x"4e",	--1798
		x"00",	--1799
		x"43",	--1800
		x"00",	--1801
		x"41",	--1802
		x"41",	--1803
		x"41",	--1804
		x"41",	--1805
		x"12",	--1806
		x"12",	--1807
		x"12",	--1808
		x"4d",	--1809
		x"4e",	--1810
		x"4d",	--1811
		x"00",	--1812
		x"4e",	--1813
		x"00",	--1814
		x"4f",	--1815
		x"49",	--1816
		x"00",	--1817
		x"43",	--1818
		x"12",	--1819
		x"dd",	--1820
		x"4e",	--1821
		x"4f",	--1822
		x"4a",	--1823
		x"4b",	--1824
		x"12",	--1825
		x"d8",	--1826
		x"4e",	--1827
		x"4f",	--1828
		x"49",	--1829
		x"00",	--1830
		x"43",	--1831
		x"12",	--1832
		x"dd",	--1833
		x"4e",	--1834
		x"4f",	--1835
		x"4a",	--1836
		x"4b",	--1837
		x"12",	--1838
		x"d7",	--1839
		x"12",	--1840
		x"d4",	--1841
		x"4e",	--1842
		x"00",	--1843
		x"41",	--1844
		x"41",	--1845
		x"41",	--1846
		x"41",	--1847
		x"4f",	--1848
		x"4e",	--1849
		x"00",	--1850
		x"41",	--1851
		x"12",	--1852
		x"12",	--1853
		x"93",	--1854
		x"02",	--1855
		x"38",	--1856
		x"40",	--1857
		x"02",	--1858
		x"43",	--1859
		x"12",	--1860
		x"4b",	--1861
		x"ff",	--1862
		x"11",	--1863
		x"12",	--1864
		x"12",	--1865
		x"ef",	--1866
		x"12",	--1867
		x"d2",	--1868
		x"50",	--1869
		x"00",	--1870
		x"53",	--1871
		x"50",	--1872
		x"00",	--1873
		x"92",	--1874
		x"02",	--1875
		x"3b",	--1876
		x"43",	--1877
		x"41",	--1878
		x"41",	--1879
		x"41",	--1880
		x"42",	--1881
		x"02",	--1882
		x"90",	--1883
		x"00",	--1884
		x"34",	--1885
		x"4e",	--1886
		x"5f",	--1887
		x"5e",	--1888
		x"5f",	--1889
		x"50",	--1890
		x"02",	--1891
		x"40",	--1892
		x"00",	--1893
		x"00",	--1894
		x"40",	--1895
		x"ce",	--1896
		x"00",	--1897
		x"40",	--1898
		x"02",	--1899
		x"00",	--1900
		x"53",	--1901
		x"4e",	--1902
		x"02",	--1903
		x"41",	--1904
		x"12",	--1905
		x"42",	--1906
		x"02",	--1907
		x"90",	--1908
		x"00",	--1909
		x"34",	--1910
		x"4b",	--1911
		x"5c",	--1912
		x"5b",	--1913
		x"5c",	--1914
		x"50",	--1915
		x"02",	--1916
		x"4f",	--1917
		x"00",	--1918
		x"4e",	--1919
		x"00",	--1920
		x"4d",	--1921
		x"00",	--1922
		x"53",	--1923
		x"4b",	--1924
		x"02",	--1925
		x"43",	--1926
		x"41",	--1927
		x"41",	--1928
		x"43",	--1929
		x"3f",	--1930
		x"12",	--1931
		x"50",	--1932
		x"ff",	--1933
		x"42",	--1934
		x"02",	--1935
		x"93",	--1936
		x"38",	--1937
		x"92",	--1938
		x"02",	--1939
		x"24",	--1940
		x"40",	--1941
		x"02",	--1942
		x"43",	--1943
		x"3c",	--1944
		x"50",	--1945
		x"00",	--1946
		x"9f",	--1947
		x"ff",	--1948
		x"24",	--1949
		x"53",	--1950
		x"9b",	--1951
		x"23",	--1952
		x"12",	--1953
		x"ef",	--1954
		x"12",	--1955
		x"d2",	--1956
		x"53",	--1957
		x"43",	--1958
		x"50",	--1959
		x"00",	--1960
		x"41",	--1961
		x"41",	--1962
		x"43",	--1963
		x"4e",	--1964
		x"00",	--1965
		x"4e",	--1966
		x"93",	--1967
		x"24",	--1968
		x"53",	--1969
		x"43",	--1970
		x"3c",	--1971
		x"4e",	--1972
		x"93",	--1973
		x"24",	--1974
		x"53",	--1975
		x"92",	--1976
		x"34",	--1977
		x"90",	--1978
		x"00",	--1979
		x"23",	--1980
		x"43",	--1981
		x"ff",	--1982
		x"4f",	--1983
		x"5d",	--1984
		x"51",	--1985
		x"4e",	--1986
		x"00",	--1987
		x"53",	--1988
		x"4e",	--1989
		x"93",	--1990
		x"23",	--1991
		x"4c",	--1992
		x"5e",	--1993
		x"5e",	--1994
		x"5c",	--1995
		x"50",	--1996
		x"02",	--1997
		x"41",	--1998
		x"12",	--1999
		x"00",	--2000
		x"50",	--2001
		x"00",	--2002
		x"41",	--2003
		x"41",	--2004
		x"43",	--2005
		x"3f",	--2006
		x"d0",	--2007
		x"02",	--2008
		x"01",	--2009
		x"40",	--2010
		x"0b",	--2011
		x"01",	--2012
		x"43",	--2013
		x"41",	--2014
		x"12",	--2015
		x"4f",	--2016
		x"42",	--2017
		x"02",	--2018
		x"90",	--2019
		x"00",	--2020
		x"34",	--2021
		x"4f",	--2022
		x"5c",	--2023
		x"4c",	--2024
		x"5d",	--2025
		x"5d",	--2026
		x"5d",	--2027
		x"8c",	--2028
		x"50",	--2029
		x"03",	--2030
		x"43",	--2031
		x"00",	--2032
		x"43",	--2033
		x"00",	--2034
		x"43",	--2035
		x"00",	--2036
		x"4b",	--2037
		x"00",	--2038
		x"4e",	--2039
		x"00",	--2040
		x"4f",	--2041
		x"53",	--2042
		x"4e",	--2043
		x"02",	--2044
		x"41",	--2045
		x"41",	--2046
		x"43",	--2047
		x"3f",	--2048
		x"5f",	--2049
		x"4f",	--2050
		x"5c",	--2051
		x"5c",	--2052
		x"5c",	--2053
		x"8f",	--2054
		x"50",	--2055
		x"03",	--2056
		x"43",	--2057
		x"00",	--2058
		x"4e",	--2059
		x"00",	--2060
		x"43",	--2061
		x"00",	--2062
		x"4d",	--2063
		x"00",	--2064
		x"43",	--2065
		x"00",	--2066
		x"43",	--2067
		x"41",	--2068
		x"5f",	--2069
		x"4f",	--2070
		x"5e",	--2071
		x"5e",	--2072
		x"5e",	--2073
		x"8f",	--2074
		x"43",	--2075
		x"03",	--2076
		x"43",	--2077
		x"41",	--2078
		x"12",	--2079
		x"12",	--2080
		x"12",	--2081
		x"12",	--2082
		x"12",	--2083
		x"12",	--2084
		x"12",	--2085
		x"12",	--2086
		x"12",	--2087
		x"93",	--2088
		x"02",	--2089
		x"38",	--2090
		x"40",	--2091
		x"03",	--2092
		x"4a",	--2093
		x"53",	--2094
		x"4a",	--2095
		x"52",	--2096
		x"4a",	--2097
		x"50",	--2098
		x"00",	--2099
		x"43",	--2100
		x"3c",	--2101
		x"53",	--2102
		x"4f",	--2103
		x"00",	--2104
		x"53",	--2105
		x"50",	--2106
		x"00",	--2107
		x"50",	--2108
		x"00",	--2109
		x"50",	--2110
		x"00",	--2111
		x"50",	--2112
		x"00",	--2113
		x"92",	--2114
		x"02",	--2115
		x"34",	--2116
		x"93",	--2117
		x"00",	--2118
		x"27",	--2119
		x"4b",	--2120
		x"9b",	--2121
		x"00",	--2122
		x"2b",	--2123
		x"43",	--2124
		x"00",	--2125
		x"4b",	--2126
		x"00",	--2127
		x"12",	--2128
		x"00",	--2129
		x"93",	--2130
		x"00",	--2131
		x"27",	--2132
		x"47",	--2133
		x"53",	--2134
		x"4f",	--2135
		x"00",	--2136
		x"98",	--2137
		x"2b",	--2138
		x"43",	--2139
		x"00",	--2140
		x"3f",	--2141
		x"f0",	--2142
		x"ff",	--2143
		x"01",	--2144
		x"41",	--2145
		x"41",	--2146
		x"41",	--2147
		x"41",	--2148
		x"41",	--2149
		x"41",	--2150
		x"41",	--2151
		x"41",	--2152
		x"41",	--2153
		x"13",	--2154
		x"4e",	--2155
		x"00",	--2156
		x"43",	--2157
		x"41",	--2158
		x"4f",	--2159
		x"4f",	--2160
		x"4f",	--2161
		x"00",	--2162
		x"41",	--2163
		x"43",	--2164
		x"00",	--2165
		x"41",	--2166
		x"4e",	--2167
		x"00",	--2168
		x"40",	--2169
		x"d0",	--2170
		x"12",	--2171
		x"cf",	--2172
		x"4f",	--2173
		x"02",	--2174
		x"43",	--2175
		x"41",	--2176
		x"4d",	--2177
		x"4f",	--2178
		x"4e",	--2179
		x"00",	--2180
		x"43",	--2181
		x"4c",	--2182
		x"42",	--2183
		x"02",	--2184
		x"12",	--2185
		x"d0",	--2186
		x"41",	--2187
		x"42",	--2188
		x"00",	--2189
		x"f2",	--2190
		x"23",	--2191
		x"4f",	--2192
		x"00",	--2193
		x"43",	--2194
		x"41",	--2195
		x"f0",	--2196
		x"00",	--2197
		x"4f",	--2198
		x"f0",	--2199
		x"11",	--2200
		x"12",	--2201
		x"d1",	--2202
		x"41",	--2203
		x"12",	--2204
		x"4f",	--2205
		x"4f",	--2206
		x"11",	--2207
		x"11",	--2208
		x"11",	--2209
		x"11",	--2210
		x"4e",	--2211
		x"12",	--2212
		x"d1",	--2213
		x"4b",	--2214
		x"12",	--2215
		x"d1",	--2216
		x"41",	--2217
		x"41",	--2218
		x"12",	--2219
		x"12",	--2220
		x"4f",	--2221
		x"40",	--2222
		x"00",	--2223
		x"4a",	--2224
		x"4b",	--2225
		x"f0",	--2226
		x"00",	--2227
		x"24",	--2228
		x"11",	--2229
		x"53",	--2230
		x"23",	--2231
		x"f3",	--2232
		x"24",	--2233
		x"40",	--2234
		x"00",	--2235
		x"12",	--2236
		x"d1",	--2237
		x"53",	--2238
		x"93",	--2239
		x"23",	--2240
		x"41",	--2241
		x"41",	--2242
		x"41",	--2243
		x"40",	--2244
		x"00",	--2245
		x"3f",	--2246
		x"12",	--2247
		x"4f",	--2248
		x"4f",	--2249
		x"10",	--2250
		x"11",	--2251
		x"4e",	--2252
		x"12",	--2253
		x"d1",	--2254
		x"4b",	--2255
		x"12",	--2256
		x"d1",	--2257
		x"41",	--2258
		x"41",	--2259
		x"12",	--2260
		x"12",	--2261
		x"4e",	--2262
		x"4f",	--2263
		x"4f",	--2264
		x"10",	--2265
		x"11",	--2266
		x"4d",	--2267
		x"12",	--2268
		x"d1",	--2269
		x"4b",	--2270
		x"12",	--2271
		x"d1",	--2272
		x"4b",	--2273
		x"4a",	--2274
		x"10",	--2275
		x"10",	--2276
		x"ec",	--2277
		x"ec",	--2278
		x"4d",	--2279
		x"12",	--2280
		x"d1",	--2281
		x"4a",	--2282
		x"12",	--2283
		x"d1",	--2284
		x"41",	--2285
		x"41",	--2286
		x"41",	--2287
		x"12",	--2288
		x"12",	--2289
		x"12",	--2290
		x"4f",	--2291
		x"93",	--2292
		x"24",	--2293
		x"4e",	--2294
		x"53",	--2295
		x"43",	--2296
		x"4a",	--2297
		x"5b",	--2298
		x"4d",	--2299
		x"11",	--2300
		x"12",	--2301
		x"d1",	--2302
		x"99",	--2303
		x"24",	--2304
		x"53",	--2305
		x"b0",	--2306
		x"00",	--2307
		x"20",	--2308
		x"40",	--2309
		x"00",	--2310
		x"12",	--2311
		x"d1",	--2312
		x"3f",	--2313
		x"40",	--2314
		x"00",	--2315
		x"12",	--2316
		x"d1",	--2317
		x"3f",	--2318
		x"41",	--2319
		x"41",	--2320
		x"41",	--2321
		x"41",	--2322
		x"12",	--2323
		x"12",	--2324
		x"12",	--2325
		x"4f",	--2326
		x"93",	--2327
		x"24",	--2328
		x"4e",	--2329
		x"53",	--2330
		x"43",	--2331
		x"4a",	--2332
		x"11",	--2333
		x"12",	--2334
		x"d1",	--2335
		x"99",	--2336
		x"24",	--2337
		x"53",	--2338
		x"b0",	--2339
		x"00",	--2340
		x"23",	--2341
		x"40",	--2342
		x"00",	--2343
		x"12",	--2344
		x"d1",	--2345
		x"4a",	--2346
		x"11",	--2347
		x"12",	--2348
		x"d1",	--2349
		x"99",	--2350
		x"23",	--2351
		x"41",	--2352
		x"41",	--2353
		x"41",	--2354
		x"41",	--2355
		x"12",	--2356
		x"12",	--2357
		x"12",	--2358
		x"50",	--2359
		x"ff",	--2360
		x"4f",	--2361
		x"93",	--2362
		x"38",	--2363
		x"90",	--2364
		x"00",	--2365
		x"38",	--2366
		x"43",	--2367
		x"41",	--2368
		x"59",	--2369
		x"40",	--2370
		x"00",	--2371
		x"4b",	--2372
		x"12",	--2373
		x"eb",	--2374
		x"50",	--2375
		x"00",	--2376
		x"4f",	--2377
		x"00",	--2378
		x"53",	--2379
		x"40",	--2380
		x"00",	--2381
		x"4b",	--2382
		x"12",	--2383
		x"eb",	--2384
		x"4f",	--2385
		x"90",	--2386
		x"00",	--2387
		x"37",	--2388
		x"49",	--2389
		x"53",	--2390
		x"51",	--2391
		x"40",	--2392
		x"00",	--2393
		x"4b",	--2394
		x"12",	--2395
		x"eb",	--2396
		x"50",	--2397
		x"00",	--2398
		x"4f",	--2399
		x"00",	--2400
		x"53",	--2401
		x"41",	--2402
		x"5a",	--2403
		x"4f",	--2404
		x"11",	--2405
		x"12",	--2406
		x"d1",	--2407
		x"93",	--2408
		x"23",	--2409
		x"50",	--2410
		x"00",	--2411
		x"41",	--2412
		x"41",	--2413
		x"41",	--2414
		x"41",	--2415
		x"40",	--2416
		x"00",	--2417
		x"12",	--2418
		x"d1",	--2419
		x"e3",	--2420
		x"53",	--2421
		x"3f",	--2422
		x"43",	--2423
		x"43",	--2424
		x"3f",	--2425
		x"12",	--2426
		x"12",	--2427
		x"12",	--2428
		x"41",	--2429
		x"52",	--2430
		x"4b",	--2431
		x"49",	--2432
		x"93",	--2433
		x"20",	--2434
		x"3c",	--2435
		x"11",	--2436
		x"12",	--2437
		x"d1",	--2438
		x"49",	--2439
		x"4a",	--2440
		x"53",	--2441
		x"4a",	--2442
		x"00",	--2443
		x"93",	--2444
		x"24",	--2445
		x"90",	--2446
		x"00",	--2447
		x"23",	--2448
		x"49",	--2449
		x"53",	--2450
		x"49",	--2451
		x"00",	--2452
		x"50",	--2453
		x"ff",	--2454
		x"90",	--2455
		x"00",	--2456
		x"2f",	--2457
		x"4f",	--2458
		x"5f",	--2459
		x"4f",	--2460
		x"ef",	--2461
		x"41",	--2462
		x"41",	--2463
		x"41",	--2464
		x"41",	--2465
		x"4b",	--2466
		x"52",	--2467
		x"4b",	--2468
		x"00",	--2469
		x"4b",	--2470
		x"12",	--2471
		x"d1",	--2472
		x"49",	--2473
		x"3f",	--2474
		x"4b",	--2475
		x"53",	--2476
		x"4b",	--2477
		x"12",	--2478
		x"d1",	--2479
		x"49",	--2480
		x"3f",	--2481
		x"4b",	--2482
		x"53",	--2483
		x"4f",	--2484
		x"49",	--2485
		x"93",	--2486
		x"27",	--2487
		x"53",	--2488
		x"11",	--2489
		x"12",	--2490
		x"d1",	--2491
		x"49",	--2492
		x"93",	--2493
		x"23",	--2494
		x"3f",	--2495
		x"4b",	--2496
		x"52",	--2497
		x"4b",	--2498
		x"00",	--2499
		x"4b",	--2500
		x"12",	--2501
		x"d2",	--2502
		x"49",	--2503
		x"3f",	--2504
		x"4b",	--2505
		x"53",	--2506
		x"4b",	--2507
		x"4e",	--2508
		x"10",	--2509
		x"11",	--2510
		x"10",	--2511
		x"11",	--2512
		x"12",	--2513
		x"d1",	--2514
		x"49",	--2515
		x"3f",	--2516
		x"4b",	--2517
		x"53",	--2518
		x"4b",	--2519
		x"12",	--2520
		x"d2",	--2521
		x"49",	--2522
		x"3f",	--2523
		x"4b",	--2524
		x"53",	--2525
		x"4b",	--2526
		x"12",	--2527
		x"d1",	--2528
		x"49",	--2529
		x"3f",	--2530
		x"4b",	--2531
		x"53",	--2532
		x"4b",	--2533
		x"12",	--2534
		x"d1",	--2535
		x"49",	--2536
		x"3f",	--2537
		x"4b",	--2538
		x"53",	--2539
		x"4b",	--2540
		x"12",	--2541
		x"d1",	--2542
		x"49",	--2543
		x"3f",	--2544
		x"40",	--2545
		x"00",	--2546
		x"12",	--2547
		x"d1",	--2548
		x"3f",	--2549
		x"12",	--2550
		x"12",	--2551
		x"42",	--2552
		x"02",	--2553
		x"42",	--2554
		x"00",	--2555
		x"04",	--2556
		x"42",	--2557
		x"02",	--2558
		x"90",	--2559
		x"00",	--2560
		x"34",	--2561
		x"53",	--2562
		x"02",	--2563
		x"42",	--2564
		x"02",	--2565
		x"42",	--2566
		x"02",	--2567
		x"9f",	--2568
		x"20",	--2569
		x"53",	--2570
		x"02",	--2571
		x"40",	--2572
		x"00",	--2573
		x"00",	--2574
		x"41",	--2575
		x"41",	--2576
		x"c0",	--2577
		x"00",	--2578
		x"00",	--2579
		x"13",	--2580
		x"43",	--2581
		x"02",	--2582
		x"3f",	--2583
		x"4e",	--2584
		x"4f",	--2585
		x"40",	--2586
		x"36",	--2587
		x"40",	--2588
		x"01",	--2589
		x"12",	--2590
		x"eb",	--2591
		x"53",	--2592
		x"4e",	--2593
		x"00",	--2594
		x"40",	--2595
		x"00",	--2596
		x"00",	--2597
		x"41",	--2598
		x"42",	--2599
		x"02",	--2600
		x"42",	--2601
		x"02",	--2602
		x"9f",	--2603
		x"38",	--2604
		x"42",	--2605
		x"02",	--2606
		x"82",	--2607
		x"02",	--2608
		x"41",	--2609
		x"42",	--2610
		x"02",	--2611
		x"42",	--2612
		x"02",	--2613
		x"40",	--2614
		x"00",	--2615
		x"8d",	--2616
		x"8e",	--2617
		x"41",	--2618
		x"42",	--2619
		x"02",	--2620
		x"4f",	--2621
		x"04",	--2622
		x"42",	--2623
		x"02",	--2624
		x"42",	--2625
		x"02",	--2626
		x"9e",	--2627
		x"24",	--2628
		x"42",	--2629
		x"02",	--2630
		x"90",	--2631
		x"00",	--2632
		x"38",	--2633
		x"43",	--2634
		x"02",	--2635
		x"41",	--2636
		x"53",	--2637
		x"02",	--2638
		x"41",	--2639
		x"43",	--2640
		x"41",	--2641
		x"12",	--2642
		x"12",	--2643
		x"4e",	--2644
		x"4f",	--2645
		x"43",	--2646
		x"40",	--2647
		x"4f",	--2648
		x"12",	--2649
		x"db",	--2650
		x"93",	--2651
		x"34",	--2652
		x"4a",	--2653
		x"4b",	--2654
		x"12",	--2655
		x"dd",	--2656
		x"41",	--2657
		x"41",	--2658
		x"41",	--2659
		x"43",	--2660
		x"40",	--2661
		x"4f",	--2662
		x"4a",	--2663
		x"4b",	--2664
		x"12",	--2665
		x"d7",	--2666
		x"12",	--2667
		x"dd",	--2668
		x"53",	--2669
		x"60",	--2670
		x"80",	--2671
		x"41",	--2672
		x"41",	--2673
		x"41",	--2674
		x"12",	--2675
		x"12",	--2676
		x"12",	--2677
		x"12",	--2678
		x"12",	--2679
		x"12",	--2680
		x"12",	--2681
		x"12",	--2682
		x"50",	--2683
		x"ff",	--2684
		x"4d",	--2685
		x"4f",	--2686
		x"93",	--2687
		x"28",	--2688
		x"4e",	--2689
		x"93",	--2690
		x"28",	--2691
		x"92",	--2692
		x"20",	--2693
		x"40",	--2694
		x"d7",	--2695
		x"92",	--2696
		x"24",	--2697
		x"93",	--2698
		x"24",	--2699
		x"93",	--2700
		x"24",	--2701
		x"4f",	--2702
		x"00",	--2703
		x"00",	--2704
		x"4e",	--2705
		x"00",	--2706
		x"4f",	--2707
		x"00",	--2708
		x"4f",	--2709
		x"00",	--2710
		x"4e",	--2711
		x"00",	--2712
		x"4e",	--2713
		x"00",	--2714
		x"41",	--2715
		x"8b",	--2716
		x"4c",	--2717
		x"93",	--2718
		x"38",	--2719
		x"90",	--2720
		x"00",	--2721
		x"34",	--2722
		x"93",	--2723
		x"38",	--2724
		x"46",	--2725
		x"00",	--2726
		x"47",	--2727
		x"00",	--2728
		x"49",	--2729
		x"f0",	--2730
		x"00",	--2731
		x"24",	--2732
		x"46",	--2733
		x"47",	--2734
		x"c3",	--2735
		x"10",	--2736
		x"10",	--2737
		x"53",	--2738
		x"23",	--2739
		x"4a",	--2740
		x"00",	--2741
		x"4b",	--2742
		x"00",	--2743
		x"43",	--2744
		x"43",	--2745
		x"f0",	--2746
		x"00",	--2747
		x"24",	--2748
		x"5c",	--2749
		x"6d",	--2750
		x"53",	--2751
		x"23",	--2752
		x"53",	--2753
		x"63",	--2754
		x"f6",	--2755
		x"f7",	--2756
		x"43",	--2757
		x"43",	--2758
		x"93",	--2759
		x"20",	--2760
		x"93",	--2761
		x"24",	--2762
		x"41",	--2763
		x"00",	--2764
		x"41",	--2765
		x"00",	--2766
		x"da",	--2767
		x"db",	--2768
		x"4f",	--2769
		x"00",	--2770
		x"9e",	--2771
		x"00",	--2772
		x"20",	--2773
		x"4f",	--2774
		x"00",	--2775
		x"41",	--2776
		x"00",	--2777
		x"46",	--2778
		x"47",	--2779
		x"54",	--2780
		x"65",	--2781
		x"4e",	--2782
		x"00",	--2783
		x"4f",	--2784
		x"00",	--2785
		x"40",	--2786
		x"00",	--2787
		x"00",	--2788
		x"93",	--2789
		x"38",	--2790
		x"48",	--2791
		x"50",	--2792
		x"00",	--2793
		x"41",	--2794
		x"41",	--2795
		x"41",	--2796
		x"41",	--2797
		x"41",	--2798
		x"41",	--2799
		x"41",	--2800
		x"41",	--2801
		x"41",	--2802
		x"91",	--2803
		x"38",	--2804
		x"4b",	--2805
		x"00",	--2806
		x"43",	--2807
		x"43",	--2808
		x"4f",	--2809
		x"00",	--2810
		x"9e",	--2811
		x"00",	--2812
		x"27",	--2813
		x"93",	--2814
		x"24",	--2815
		x"46",	--2816
		x"47",	--2817
		x"84",	--2818
		x"75",	--2819
		x"93",	--2820
		x"38",	--2821
		x"43",	--2822
		x"00",	--2823
		x"41",	--2824
		x"00",	--2825
		x"4e",	--2826
		x"00",	--2827
		x"4f",	--2828
		x"00",	--2829
		x"4e",	--2830
		x"4f",	--2831
		x"53",	--2832
		x"63",	--2833
		x"90",	--2834
		x"3f",	--2835
		x"28",	--2836
		x"90",	--2837
		x"40",	--2838
		x"2c",	--2839
		x"93",	--2840
		x"2c",	--2841
		x"48",	--2842
		x"00",	--2843
		x"53",	--2844
		x"5e",	--2845
		x"6f",	--2846
		x"4b",	--2847
		x"53",	--2848
		x"4e",	--2849
		x"4f",	--2850
		x"53",	--2851
		x"63",	--2852
		x"90",	--2853
		x"3f",	--2854
		x"2b",	--2855
		x"24",	--2856
		x"4e",	--2857
		x"00",	--2858
		x"4f",	--2859
		x"00",	--2860
		x"4a",	--2861
		x"00",	--2862
		x"40",	--2863
		x"00",	--2864
		x"00",	--2865
		x"93",	--2866
		x"37",	--2867
		x"4e",	--2868
		x"4f",	--2869
		x"f3",	--2870
		x"f3",	--2871
		x"c3",	--2872
		x"10",	--2873
		x"10",	--2874
		x"4c",	--2875
		x"4d",	--2876
		x"de",	--2877
		x"df",	--2878
		x"4a",	--2879
		x"00",	--2880
		x"4b",	--2881
		x"00",	--2882
		x"53",	--2883
		x"00",	--2884
		x"48",	--2885
		x"3f",	--2886
		x"93",	--2887
		x"23",	--2888
		x"4f",	--2889
		x"00",	--2890
		x"4f",	--2891
		x"00",	--2892
		x"00",	--2893
		x"4f",	--2894
		x"00",	--2895
		x"00",	--2896
		x"4f",	--2897
		x"00",	--2898
		x"00",	--2899
		x"4e",	--2900
		x"00",	--2901
		x"ff",	--2902
		x"00",	--2903
		x"4e",	--2904
		x"00",	--2905
		x"4d",	--2906
		x"3f",	--2907
		x"43",	--2908
		x"43",	--2909
		x"3f",	--2910
		x"e3",	--2911
		x"53",	--2912
		x"90",	--2913
		x"00",	--2914
		x"37",	--2915
		x"3f",	--2916
		x"93",	--2917
		x"2b",	--2918
		x"3f",	--2919
		x"44",	--2920
		x"45",	--2921
		x"86",	--2922
		x"77",	--2923
		x"3f",	--2924
		x"4e",	--2925
		x"3f",	--2926
		x"43",	--2927
		x"00",	--2928
		x"41",	--2929
		x"00",	--2930
		x"e3",	--2931
		x"e3",	--2932
		x"53",	--2933
		x"63",	--2934
		x"4e",	--2935
		x"00",	--2936
		x"4f",	--2937
		x"00",	--2938
		x"3f",	--2939
		x"93",	--2940
		x"27",	--2941
		x"59",	--2942
		x"00",	--2943
		x"44",	--2944
		x"00",	--2945
		x"45",	--2946
		x"00",	--2947
		x"49",	--2948
		x"f0",	--2949
		x"00",	--2950
		x"24",	--2951
		x"4d",	--2952
		x"44",	--2953
		x"45",	--2954
		x"c3",	--2955
		x"10",	--2956
		x"10",	--2957
		x"53",	--2958
		x"23",	--2959
		x"4c",	--2960
		x"00",	--2961
		x"4d",	--2962
		x"00",	--2963
		x"43",	--2964
		x"43",	--2965
		x"f0",	--2966
		x"00",	--2967
		x"24",	--2968
		x"5c",	--2969
		x"6d",	--2970
		x"53",	--2971
		x"23",	--2972
		x"53",	--2973
		x"63",	--2974
		x"f4",	--2975
		x"f5",	--2976
		x"43",	--2977
		x"43",	--2978
		x"93",	--2979
		x"20",	--2980
		x"93",	--2981
		x"20",	--2982
		x"43",	--2983
		x"43",	--2984
		x"41",	--2985
		x"00",	--2986
		x"41",	--2987
		x"00",	--2988
		x"da",	--2989
		x"db",	--2990
		x"3f",	--2991
		x"43",	--2992
		x"43",	--2993
		x"3f",	--2994
		x"92",	--2995
		x"23",	--2996
		x"9e",	--2997
		x"00",	--2998
		x"00",	--2999
		x"27",	--3000
		x"40",	--3001
		x"f0",	--3002
		x"3f",	--3003
		x"50",	--3004
		x"ff",	--3005
		x"4e",	--3006
		x"00",	--3007
		x"4f",	--3008
		x"00",	--3009
		x"4c",	--3010
		x"00",	--3011
		x"4d",	--3012
		x"00",	--3013
		x"41",	--3014
		x"50",	--3015
		x"00",	--3016
		x"41",	--3017
		x"52",	--3018
		x"12",	--3019
		x"e0",	--3020
		x"41",	--3021
		x"50",	--3022
		x"00",	--3023
		x"41",	--3024
		x"12",	--3025
		x"e0",	--3026
		x"41",	--3027
		x"52",	--3028
		x"41",	--3029
		x"50",	--3030
		x"00",	--3031
		x"41",	--3032
		x"50",	--3033
		x"00",	--3034
		x"12",	--3035
		x"d4",	--3036
		x"12",	--3037
		x"df",	--3038
		x"50",	--3039
		x"00",	--3040
		x"41",	--3041
		x"50",	--3042
		x"ff",	--3043
		x"4e",	--3044
		x"00",	--3045
		x"4f",	--3046
		x"00",	--3047
		x"4c",	--3048
		x"00",	--3049
		x"4d",	--3050
		x"00",	--3051
		x"41",	--3052
		x"50",	--3053
		x"00",	--3054
		x"41",	--3055
		x"52",	--3056
		x"12",	--3057
		x"e0",	--3058
		x"41",	--3059
		x"50",	--3060
		x"00",	--3061
		x"41",	--3062
		x"12",	--3063
		x"e0",	--3064
		x"e3",	--3065
		x"00",	--3066
		x"41",	--3067
		x"52",	--3068
		x"41",	--3069
		x"50",	--3070
		x"00",	--3071
		x"41",	--3072
		x"50",	--3073
		x"00",	--3074
		x"12",	--3075
		x"d4",	--3076
		x"12",	--3077
		x"df",	--3078
		x"50",	--3079
		x"00",	--3080
		x"41",	--3081
		x"12",	--3082
		x"12",	--3083
		x"12",	--3084
		x"12",	--3085
		x"12",	--3086
		x"12",	--3087
		x"12",	--3088
		x"12",	--3089
		x"50",	--3090
		x"ff",	--3091
		x"4e",	--3092
		x"00",	--3093
		x"4f",	--3094
		x"00",	--3095
		x"4c",	--3096
		x"00",	--3097
		x"4d",	--3098
		x"00",	--3099
		x"41",	--3100
		x"50",	--3101
		x"00",	--3102
		x"41",	--3103
		x"52",	--3104
		x"12",	--3105
		x"e0",	--3106
		x"41",	--3107
		x"50",	--3108
		x"00",	--3109
		x"41",	--3110
		x"12",	--3111
		x"e0",	--3112
		x"41",	--3113
		x"00",	--3114
		x"93",	--3115
		x"28",	--3116
		x"41",	--3117
		x"00",	--3118
		x"93",	--3119
		x"28",	--3120
		x"92",	--3121
		x"24",	--3122
		x"92",	--3123
		x"24",	--3124
		x"93",	--3125
		x"24",	--3126
		x"93",	--3127
		x"24",	--3128
		x"41",	--3129
		x"00",	--3130
		x"41",	--3131
		x"00",	--3132
		x"41",	--3133
		x"00",	--3134
		x"41",	--3135
		x"00",	--3136
		x"40",	--3137
		x"00",	--3138
		x"43",	--3139
		x"43",	--3140
		x"43",	--3141
		x"43",	--3142
		x"43",	--3143
		x"00",	--3144
		x"43",	--3145
		x"00",	--3146
		x"43",	--3147
		x"43",	--3148
		x"4c",	--3149
		x"00",	--3150
		x"3c",	--3151
		x"58",	--3152
		x"69",	--3153
		x"c3",	--3154
		x"10",	--3155
		x"10",	--3156
		x"53",	--3157
		x"00",	--3158
		x"24",	--3159
		x"b3",	--3160
		x"24",	--3161
		x"58",	--3162
		x"69",	--3163
		x"56",	--3164
		x"67",	--3165
		x"43",	--3166
		x"43",	--3167
		x"99",	--3168
		x"28",	--3169
		x"24",	--3170
		x"43",	--3171
		x"43",	--3172
		x"5c",	--3173
		x"6d",	--3174
		x"56",	--3175
		x"67",	--3176
		x"93",	--3177
		x"37",	--3178
		x"d3",	--3179
		x"d3",	--3180
		x"3f",	--3181
		x"98",	--3182
		x"2b",	--3183
		x"3f",	--3184
		x"4a",	--3185
		x"00",	--3186
		x"4b",	--3187
		x"00",	--3188
		x"4f",	--3189
		x"41",	--3190
		x"00",	--3191
		x"51",	--3192
		x"00",	--3193
		x"4a",	--3194
		x"53",	--3195
		x"46",	--3196
		x"00",	--3197
		x"43",	--3198
		x"91",	--3199
		x"00",	--3200
		x"00",	--3201
		x"24",	--3202
		x"4d",	--3203
		x"00",	--3204
		x"93",	--3205
		x"38",	--3206
		x"90",	--3207
		x"40",	--3208
		x"2c",	--3209
		x"41",	--3210
		x"00",	--3211
		x"53",	--3212
		x"41",	--3213
		x"00",	--3214
		x"41",	--3215
		x"00",	--3216
		x"4d",	--3217
		x"5e",	--3218
		x"6f",	--3219
		x"93",	--3220
		x"38",	--3221
		x"5a",	--3222
		x"6b",	--3223
		x"53",	--3224
		x"90",	--3225
		x"40",	--3226
		x"2b",	--3227
		x"4a",	--3228
		x"00",	--3229
		x"4b",	--3230
		x"00",	--3231
		x"4c",	--3232
		x"00",	--3233
		x"4e",	--3234
		x"4f",	--3235
		x"f0",	--3236
		x"00",	--3237
		x"f3",	--3238
		x"90",	--3239
		x"00",	--3240
		x"24",	--3241
		x"4e",	--3242
		x"00",	--3243
		x"4f",	--3244
		x"00",	--3245
		x"40",	--3246
		x"00",	--3247
		x"00",	--3248
		x"41",	--3249
		x"52",	--3250
		x"12",	--3251
		x"df",	--3252
		x"50",	--3253
		x"00",	--3254
		x"41",	--3255
		x"41",	--3256
		x"41",	--3257
		x"41",	--3258
		x"41",	--3259
		x"41",	--3260
		x"41",	--3261
		x"41",	--3262
		x"41",	--3263
		x"d3",	--3264
		x"d3",	--3265
		x"3f",	--3266
		x"50",	--3267
		x"00",	--3268
		x"4a",	--3269
		x"b3",	--3270
		x"24",	--3271
		x"41",	--3272
		x"00",	--3273
		x"41",	--3274
		x"00",	--3275
		x"c3",	--3276
		x"10",	--3277
		x"10",	--3278
		x"4c",	--3279
		x"4d",	--3280
		x"d3",	--3281
		x"d0",	--3282
		x"80",	--3283
		x"46",	--3284
		x"00",	--3285
		x"47",	--3286
		x"00",	--3287
		x"c3",	--3288
		x"10",	--3289
		x"10",	--3290
		x"53",	--3291
		x"93",	--3292
		x"3b",	--3293
		x"48",	--3294
		x"00",	--3295
		x"3f",	--3296
		x"93",	--3297
		x"24",	--3298
		x"43",	--3299
		x"91",	--3300
		x"00",	--3301
		x"00",	--3302
		x"24",	--3303
		x"4f",	--3304
		x"00",	--3305
		x"41",	--3306
		x"50",	--3307
		x"00",	--3308
		x"3f",	--3309
		x"93",	--3310
		x"23",	--3311
		x"4e",	--3312
		x"4f",	--3313
		x"f0",	--3314
		x"00",	--3315
		x"f3",	--3316
		x"93",	--3317
		x"23",	--3318
		x"93",	--3319
		x"23",	--3320
		x"93",	--3321
		x"00",	--3322
		x"20",	--3323
		x"93",	--3324
		x"00",	--3325
		x"27",	--3326
		x"50",	--3327
		x"00",	--3328
		x"63",	--3329
		x"f0",	--3330
		x"ff",	--3331
		x"f3",	--3332
		x"3f",	--3333
		x"43",	--3334
		x"3f",	--3335
		x"43",	--3336
		x"3f",	--3337
		x"43",	--3338
		x"91",	--3339
		x"00",	--3340
		x"00",	--3341
		x"24",	--3342
		x"4f",	--3343
		x"00",	--3344
		x"41",	--3345
		x"50",	--3346
		x"00",	--3347
		x"3f",	--3348
		x"43",	--3349
		x"3f",	--3350
		x"93",	--3351
		x"23",	--3352
		x"40",	--3353
		x"f0",	--3354
		x"3f",	--3355
		x"12",	--3356
		x"12",	--3357
		x"12",	--3358
		x"12",	--3359
		x"12",	--3360
		x"50",	--3361
		x"ff",	--3362
		x"4e",	--3363
		x"00",	--3364
		x"4f",	--3365
		x"00",	--3366
		x"4c",	--3367
		x"00",	--3368
		x"4d",	--3369
		x"00",	--3370
		x"41",	--3371
		x"50",	--3372
		x"00",	--3373
		x"41",	--3374
		x"52",	--3375
		x"12",	--3376
		x"e0",	--3377
		x"41",	--3378
		x"52",	--3379
		x"41",	--3380
		x"12",	--3381
		x"e0",	--3382
		x"41",	--3383
		x"00",	--3384
		x"93",	--3385
		x"28",	--3386
		x"41",	--3387
		x"00",	--3388
		x"93",	--3389
		x"28",	--3390
		x"e1",	--3391
		x"00",	--3392
		x"00",	--3393
		x"92",	--3394
		x"24",	--3395
		x"93",	--3396
		x"24",	--3397
		x"92",	--3398
		x"24",	--3399
		x"93",	--3400
		x"24",	--3401
		x"41",	--3402
		x"00",	--3403
		x"81",	--3404
		x"00",	--3405
		x"4d",	--3406
		x"00",	--3407
		x"41",	--3408
		x"00",	--3409
		x"41",	--3410
		x"00",	--3411
		x"41",	--3412
		x"00",	--3413
		x"41",	--3414
		x"00",	--3415
		x"99",	--3416
		x"2c",	--3417
		x"5e",	--3418
		x"6f",	--3419
		x"53",	--3420
		x"4d",	--3421
		x"00",	--3422
		x"40",	--3423
		x"00",	--3424
		x"43",	--3425
		x"40",	--3426
		x"40",	--3427
		x"43",	--3428
		x"43",	--3429
		x"3c",	--3430
		x"dc",	--3431
		x"dd",	--3432
		x"88",	--3433
		x"79",	--3434
		x"c3",	--3435
		x"10",	--3436
		x"10",	--3437
		x"5e",	--3438
		x"6f",	--3439
		x"53",	--3440
		x"24",	--3441
		x"99",	--3442
		x"2b",	--3443
		x"23",	--3444
		x"98",	--3445
		x"2b",	--3446
		x"3f",	--3447
		x"9f",	--3448
		x"2b",	--3449
		x"98",	--3450
		x"2f",	--3451
		x"3f",	--3452
		x"4a",	--3453
		x"4b",	--3454
		x"f0",	--3455
		x"00",	--3456
		x"f3",	--3457
		x"90",	--3458
		x"00",	--3459
		x"24",	--3460
		x"4a",	--3461
		x"00",	--3462
		x"4b",	--3463
		x"00",	--3464
		x"41",	--3465
		x"50",	--3466
		x"00",	--3467
		x"12",	--3468
		x"df",	--3469
		x"50",	--3470
		x"00",	--3471
		x"41",	--3472
		x"41",	--3473
		x"41",	--3474
		x"41",	--3475
		x"41",	--3476
		x"41",	--3477
		x"42",	--3478
		x"00",	--3479
		x"41",	--3480
		x"50",	--3481
		x"00",	--3482
		x"3f",	--3483
		x"9e",	--3484
		x"23",	--3485
		x"40",	--3486
		x"f0",	--3487
		x"3f",	--3488
		x"93",	--3489
		x"23",	--3490
		x"4a",	--3491
		x"4b",	--3492
		x"f0",	--3493
		x"00",	--3494
		x"f3",	--3495
		x"93",	--3496
		x"23",	--3497
		x"93",	--3498
		x"23",	--3499
		x"93",	--3500
		x"20",	--3501
		x"93",	--3502
		x"27",	--3503
		x"50",	--3504
		x"00",	--3505
		x"63",	--3506
		x"f0",	--3507
		x"ff",	--3508
		x"f3",	--3509
		x"3f",	--3510
		x"43",	--3511
		x"00",	--3512
		x"43",	--3513
		x"00",	--3514
		x"43",	--3515
		x"00",	--3516
		x"41",	--3517
		x"50",	--3518
		x"00",	--3519
		x"3f",	--3520
		x"41",	--3521
		x"52",	--3522
		x"3f",	--3523
		x"50",	--3524
		x"ff",	--3525
		x"4e",	--3526
		x"00",	--3527
		x"4f",	--3528
		x"00",	--3529
		x"4c",	--3530
		x"00",	--3531
		x"4d",	--3532
		x"00",	--3533
		x"41",	--3534
		x"50",	--3535
		x"00",	--3536
		x"41",	--3537
		x"52",	--3538
		x"12",	--3539
		x"e0",	--3540
		x"41",	--3541
		x"52",	--3542
		x"41",	--3543
		x"12",	--3544
		x"e0",	--3545
		x"93",	--3546
		x"00",	--3547
		x"28",	--3548
		x"93",	--3549
		x"00",	--3550
		x"28",	--3551
		x"41",	--3552
		x"52",	--3553
		x"41",	--3554
		x"50",	--3555
		x"00",	--3556
		x"12",	--3557
		x"e2",	--3558
		x"50",	--3559
		x"00",	--3560
		x"41",	--3561
		x"43",	--3562
		x"3f",	--3563
		x"50",	--3564
		x"ff",	--3565
		x"4e",	--3566
		x"00",	--3567
		x"4f",	--3568
		x"00",	--3569
		x"4c",	--3570
		x"00",	--3571
		x"4d",	--3572
		x"00",	--3573
		x"41",	--3574
		x"50",	--3575
		x"00",	--3576
		x"41",	--3577
		x"52",	--3578
		x"12",	--3579
		x"e0",	--3580
		x"41",	--3581
		x"52",	--3582
		x"41",	--3583
		x"12",	--3584
		x"e0",	--3585
		x"93",	--3586
		x"00",	--3587
		x"28",	--3588
		x"93",	--3589
		x"00",	--3590
		x"28",	--3591
		x"41",	--3592
		x"52",	--3593
		x"41",	--3594
		x"50",	--3595
		x"00",	--3596
		x"12",	--3597
		x"e2",	--3598
		x"50",	--3599
		x"00",	--3600
		x"41",	--3601
		x"43",	--3602
		x"3f",	--3603
		x"50",	--3604
		x"ff",	--3605
		x"4e",	--3606
		x"00",	--3607
		x"4f",	--3608
		x"00",	--3609
		x"4c",	--3610
		x"00",	--3611
		x"4d",	--3612
		x"00",	--3613
		x"41",	--3614
		x"50",	--3615
		x"00",	--3616
		x"41",	--3617
		x"52",	--3618
		x"12",	--3619
		x"e0",	--3620
		x"41",	--3621
		x"52",	--3622
		x"41",	--3623
		x"12",	--3624
		x"e0",	--3625
		x"93",	--3626
		x"00",	--3627
		x"28",	--3628
		x"93",	--3629
		x"00",	--3630
		x"28",	--3631
		x"41",	--3632
		x"52",	--3633
		x"41",	--3634
		x"50",	--3635
		x"00",	--3636
		x"12",	--3637
		x"e2",	--3638
		x"50",	--3639
		x"00",	--3640
		x"41",	--3641
		x"43",	--3642
		x"3f",	--3643
		x"12",	--3644
		x"12",	--3645
		x"82",	--3646
		x"40",	--3647
		x"00",	--3648
		x"00",	--3649
		x"4f",	--3650
		x"5d",	--3651
		x"43",	--3652
		x"6d",	--3653
		x"4d",	--3654
		x"4d",	--3655
		x"00",	--3656
		x"93",	--3657
		x"20",	--3658
		x"93",	--3659
		x"20",	--3660
		x"43",	--3661
		x"00",	--3662
		x"41",	--3663
		x"12",	--3664
		x"df",	--3665
		x"52",	--3666
		x"41",	--3667
		x"41",	--3668
		x"41",	--3669
		x"40",	--3670
		x"00",	--3671
		x"00",	--3672
		x"93",	--3673
		x"20",	--3674
		x"4e",	--3675
		x"4f",	--3676
		x"4a",	--3677
		x"00",	--3678
		x"4b",	--3679
		x"00",	--3680
		x"4a",	--3681
		x"4b",	--3682
		x"12",	--3683
		x"de",	--3684
		x"53",	--3685
		x"93",	--3686
		x"3b",	--3687
		x"4a",	--3688
		x"00",	--3689
		x"4b",	--3690
		x"00",	--3691
		x"4f",	--3692
		x"f0",	--3693
		x"00",	--3694
		x"20",	--3695
		x"40",	--3696
		x"00",	--3697
		x"8f",	--3698
		x"4e",	--3699
		x"00",	--3700
		x"3f",	--3701
		x"93",	--3702
		x"24",	--3703
		x"4e",	--3704
		x"4f",	--3705
		x"e3",	--3706
		x"e3",	--3707
		x"53",	--3708
		x"63",	--3709
		x"3f",	--3710
		x"51",	--3711
		x"00",	--3712
		x"00",	--3713
		x"61",	--3714
		x"00",	--3715
		x"00",	--3716
		x"53",	--3717
		x"23",	--3718
		x"3f",	--3719
		x"90",	--3720
		x"80",	--3721
		x"23",	--3722
		x"43",	--3723
		x"40",	--3724
		x"cf",	--3725
		x"3f",	--3726
		x"50",	--3727
		x"ff",	--3728
		x"4e",	--3729
		x"00",	--3730
		x"4f",	--3731
		x"00",	--3732
		x"41",	--3733
		x"52",	--3734
		x"41",	--3735
		x"12",	--3736
		x"e0",	--3737
		x"41",	--3738
		x"00",	--3739
		x"93",	--3740
		x"24",	--3741
		x"28",	--3742
		x"92",	--3743
		x"24",	--3744
		x"41",	--3745
		x"00",	--3746
		x"93",	--3747
		x"38",	--3748
		x"90",	--3749
		x"00",	--3750
		x"38",	--3751
		x"93",	--3752
		x"00",	--3753
		x"20",	--3754
		x"43",	--3755
		x"40",	--3756
		x"7f",	--3757
		x"50",	--3758
		x"00",	--3759
		x"41",	--3760
		x"41",	--3761
		x"00",	--3762
		x"41",	--3763
		x"00",	--3764
		x"40",	--3765
		x"00",	--3766
		x"8d",	--3767
		x"4c",	--3768
		x"f0",	--3769
		x"00",	--3770
		x"20",	--3771
		x"93",	--3772
		x"00",	--3773
		x"27",	--3774
		x"e3",	--3775
		x"e3",	--3776
		x"53",	--3777
		x"63",	--3778
		x"50",	--3779
		x"00",	--3780
		x"41",	--3781
		x"43",	--3782
		x"43",	--3783
		x"50",	--3784
		x"00",	--3785
		x"41",	--3786
		x"c3",	--3787
		x"10",	--3788
		x"10",	--3789
		x"53",	--3790
		x"23",	--3791
		x"3f",	--3792
		x"43",	--3793
		x"40",	--3794
		x"80",	--3795
		x"50",	--3796
		x"00",	--3797
		x"41",	--3798
		x"12",	--3799
		x"12",	--3800
		x"12",	--3801
		x"12",	--3802
		x"82",	--3803
		x"4e",	--3804
		x"4f",	--3805
		x"43",	--3806
		x"00",	--3807
		x"93",	--3808
		x"20",	--3809
		x"93",	--3810
		x"20",	--3811
		x"43",	--3812
		x"00",	--3813
		x"41",	--3814
		x"12",	--3815
		x"df",	--3816
		x"52",	--3817
		x"41",	--3818
		x"41",	--3819
		x"41",	--3820
		x"41",	--3821
		x"41",	--3822
		x"40",	--3823
		x"00",	--3824
		x"00",	--3825
		x"40",	--3826
		x"00",	--3827
		x"00",	--3828
		x"4a",	--3829
		x"00",	--3830
		x"4b",	--3831
		x"00",	--3832
		x"4a",	--3833
		x"4b",	--3834
		x"12",	--3835
		x"de",	--3836
		x"53",	--3837
		x"93",	--3838
		x"38",	--3839
		x"27",	--3840
		x"4a",	--3841
		x"00",	--3842
		x"4b",	--3843
		x"00",	--3844
		x"4f",	--3845
		x"f0",	--3846
		x"00",	--3847
		x"20",	--3848
		x"40",	--3849
		x"00",	--3850
		x"8f",	--3851
		x"4e",	--3852
		x"00",	--3853
		x"3f",	--3854
		x"51",	--3855
		x"00",	--3856
		x"00",	--3857
		x"61",	--3858
		x"00",	--3859
		x"00",	--3860
		x"53",	--3861
		x"23",	--3862
		x"3f",	--3863
		x"4f",	--3864
		x"e3",	--3865
		x"53",	--3866
		x"43",	--3867
		x"43",	--3868
		x"4e",	--3869
		x"f0",	--3870
		x"00",	--3871
		x"24",	--3872
		x"5c",	--3873
		x"6d",	--3874
		x"53",	--3875
		x"23",	--3876
		x"53",	--3877
		x"63",	--3878
		x"fa",	--3879
		x"fb",	--3880
		x"43",	--3881
		x"43",	--3882
		x"93",	--3883
		x"20",	--3884
		x"93",	--3885
		x"20",	--3886
		x"43",	--3887
		x"43",	--3888
		x"f0",	--3889
		x"00",	--3890
		x"20",	--3891
		x"48",	--3892
		x"49",	--3893
		x"da",	--3894
		x"db",	--3895
		x"4d",	--3896
		x"00",	--3897
		x"4e",	--3898
		x"00",	--3899
		x"40",	--3900
		x"00",	--3901
		x"8f",	--3902
		x"4e",	--3903
		x"00",	--3904
		x"3f",	--3905
		x"c3",	--3906
		x"10",	--3907
		x"10",	--3908
		x"53",	--3909
		x"23",	--3910
		x"3f",	--3911
		x"12",	--3912
		x"12",	--3913
		x"12",	--3914
		x"93",	--3915
		x"2c",	--3916
		x"90",	--3917
		x"01",	--3918
		x"28",	--3919
		x"40",	--3920
		x"00",	--3921
		x"43",	--3922
		x"42",	--3923
		x"4e",	--3924
		x"4f",	--3925
		x"49",	--3926
		x"93",	--3927
		x"20",	--3928
		x"50",	--3929
		x"f0",	--3930
		x"4c",	--3931
		x"43",	--3932
		x"8e",	--3933
		x"7f",	--3934
		x"4a",	--3935
		x"41",	--3936
		x"41",	--3937
		x"41",	--3938
		x"41",	--3939
		x"90",	--3940
		x"01",	--3941
		x"28",	--3942
		x"42",	--3943
		x"43",	--3944
		x"40",	--3945
		x"00",	--3946
		x"4e",	--3947
		x"4f",	--3948
		x"49",	--3949
		x"93",	--3950
		x"27",	--3951
		x"c3",	--3952
		x"10",	--3953
		x"10",	--3954
		x"53",	--3955
		x"23",	--3956
		x"3f",	--3957
		x"40",	--3958
		x"00",	--3959
		x"43",	--3960
		x"40",	--3961
		x"00",	--3962
		x"3f",	--3963
		x"40",	--3964
		x"00",	--3965
		x"43",	--3966
		x"43",	--3967
		x"3f",	--3968
		x"12",	--3969
		x"12",	--3970
		x"12",	--3971
		x"12",	--3972
		x"12",	--3973
		x"4f",	--3974
		x"4f",	--3975
		x"00",	--3976
		x"4f",	--3977
		x"00",	--3978
		x"4d",	--3979
		x"00",	--3980
		x"4d",	--3981
		x"93",	--3982
		x"28",	--3983
		x"92",	--3984
		x"24",	--3985
		x"93",	--3986
		x"24",	--3987
		x"93",	--3988
		x"24",	--3989
		x"4d",	--3990
		x"00",	--3991
		x"90",	--3992
		x"ff",	--3993
		x"38",	--3994
		x"90",	--3995
		x"00",	--3996
		x"34",	--3997
		x"4e",	--3998
		x"4f",	--3999
		x"f0",	--4000
		x"00",	--4001
		x"f3",	--4002
		x"90",	--4003
		x"00",	--4004
		x"24",	--4005
		x"50",	--4006
		x"00",	--4007
		x"63",	--4008
		x"93",	--4009
		x"38",	--4010
		x"4b",	--4011
		x"50",	--4012
		x"00",	--4013
		x"c3",	--4014
		x"10",	--4015
		x"10",	--4016
		x"c3",	--4017
		x"10",	--4018
		x"10",	--4019
		x"c3",	--4020
		x"10",	--4021
		x"10",	--4022
		x"c3",	--4023
		x"10",	--4024
		x"10",	--4025
		x"c3",	--4026
		x"10",	--4027
		x"10",	--4028
		x"c3",	--4029
		x"10",	--4030
		x"10",	--4031
		x"c3",	--4032
		x"10",	--4033
		x"10",	--4034
		x"f3",	--4035
		x"f0",	--4036
		x"00",	--4037
		x"4d",	--4038
		x"3c",	--4039
		x"93",	--4040
		x"23",	--4041
		x"43",	--4042
		x"43",	--4043
		x"43",	--4044
		x"4d",	--4045
		x"5d",	--4046
		x"5d",	--4047
		x"5d",	--4048
		x"5d",	--4049
		x"5d",	--4050
		x"5d",	--4051
		x"5d",	--4052
		x"4f",	--4053
		x"f0",	--4054
		x"00",	--4055
		x"dd",	--4056
		x"4a",	--4057
		x"11",	--4058
		x"43",	--4059
		x"10",	--4060
		x"4c",	--4061
		x"df",	--4062
		x"4d",	--4063
		x"41",	--4064
		x"41",	--4065
		x"41",	--4066
		x"41",	--4067
		x"41",	--4068
		x"41",	--4069
		x"93",	--4070
		x"23",	--4071
		x"4e",	--4072
		x"4f",	--4073
		x"f0",	--4074
		x"00",	--4075
		x"f3",	--4076
		x"93",	--4077
		x"20",	--4078
		x"93",	--4079
		x"27",	--4080
		x"50",	--4081
		x"00",	--4082
		x"63",	--4083
		x"3f",	--4084
		x"c3",	--4085
		x"10",	--4086
		x"10",	--4087
		x"4b",	--4088
		x"50",	--4089
		x"00",	--4090
		x"3f",	--4091
		x"43",	--4092
		x"43",	--4093
		x"43",	--4094
		x"3f",	--4095
		x"d3",	--4096
		x"d0",	--4097
		x"00",	--4098
		x"f3",	--4099
		x"f0",	--4100
		x"00",	--4101
		x"43",	--4102
		x"3f",	--4103
		x"40",	--4104
		x"ff",	--4105
		x"8b",	--4106
		x"90",	--4107
		x"00",	--4108
		x"34",	--4109
		x"4e",	--4110
		x"4f",	--4111
		x"47",	--4112
		x"f0",	--4113
		x"00",	--4114
		x"24",	--4115
		x"c3",	--4116
		x"10",	--4117
		x"10",	--4118
		x"53",	--4119
		x"23",	--4120
		x"43",	--4121
		x"43",	--4122
		x"f0",	--4123
		x"00",	--4124
		x"24",	--4125
		x"58",	--4126
		x"69",	--4127
		x"53",	--4128
		x"23",	--4129
		x"53",	--4130
		x"63",	--4131
		x"fe",	--4132
		x"ff",	--4133
		x"43",	--4134
		x"43",	--4135
		x"93",	--4136
		x"20",	--4137
		x"93",	--4138
		x"20",	--4139
		x"43",	--4140
		x"43",	--4141
		x"4e",	--4142
		x"4f",	--4143
		x"dc",	--4144
		x"dd",	--4145
		x"48",	--4146
		x"49",	--4147
		x"f0",	--4148
		x"00",	--4149
		x"f3",	--4150
		x"90",	--4151
		x"00",	--4152
		x"24",	--4153
		x"50",	--4154
		x"00",	--4155
		x"63",	--4156
		x"48",	--4157
		x"49",	--4158
		x"c3",	--4159
		x"10",	--4160
		x"10",	--4161
		x"c3",	--4162
		x"10",	--4163
		x"10",	--4164
		x"c3",	--4165
		x"10",	--4166
		x"10",	--4167
		x"c3",	--4168
		x"10",	--4169
		x"10",	--4170
		x"c3",	--4171
		x"10",	--4172
		x"10",	--4173
		x"c3",	--4174
		x"10",	--4175
		x"10",	--4176
		x"c3",	--4177
		x"10",	--4178
		x"10",	--4179
		x"f3",	--4180
		x"f0",	--4181
		x"00",	--4182
		x"43",	--4183
		x"90",	--4184
		x"40",	--4185
		x"2f",	--4186
		x"43",	--4187
		x"3f",	--4188
		x"43",	--4189
		x"43",	--4190
		x"3f",	--4191
		x"93",	--4192
		x"23",	--4193
		x"48",	--4194
		x"49",	--4195
		x"f0",	--4196
		x"00",	--4197
		x"f3",	--4198
		x"93",	--4199
		x"24",	--4200
		x"50",	--4201
		x"00",	--4202
		x"63",	--4203
		x"3f",	--4204
		x"93",	--4205
		x"27",	--4206
		x"3f",	--4207
		x"12",	--4208
		x"12",	--4209
		x"4f",	--4210
		x"4f",	--4211
		x"00",	--4212
		x"f0",	--4213
		x"00",	--4214
		x"4f",	--4215
		x"00",	--4216
		x"c3",	--4217
		x"10",	--4218
		x"c3",	--4219
		x"10",	--4220
		x"c3",	--4221
		x"10",	--4222
		x"c3",	--4223
		x"10",	--4224
		x"c3",	--4225
		x"10",	--4226
		x"c3",	--4227
		x"10",	--4228
		x"c3",	--4229
		x"10",	--4230
		x"4d",	--4231
		x"4f",	--4232
		x"00",	--4233
		x"b0",	--4234
		x"00",	--4235
		x"43",	--4236
		x"6f",	--4237
		x"4f",	--4238
		x"00",	--4239
		x"93",	--4240
		x"20",	--4241
		x"93",	--4242
		x"24",	--4243
		x"40",	--4244
		x"ff",	--4245
		x"00",	--4246
		x"4a",	--4247
		x"4b",	--4248
		x"5c",	--4249
		x"6d",	--4250
		x"5c",	--4251
		x"6d",	--4252
		x"5c",	--4253
		x"6d",	--4254
		x"5c",	--4255
		x"6d",	--4256
		x"5c",	--4257
		x"6d",	--4258
		x"5c",	--4259
		x"6d",	--4260
		x"5c",	--4261
		x"6d",	--4262
		x"40",	--4263
		x"00",	--4264
		x"00",	--4265
		x"90",	--4266
		x"40",	--4267
		x"2c",	--4268
		x"40",	--4269
		x"ff",	--4270
		x"5c",	--4271
		x"6d",	--4272
		x"4f",	--4273
		x"53",	--4274
		x"90",	--4275
		x"40",	--4276
		x"2b",	--4277
		x"4a",	--4278
		x"00",	--4279
		x"4c",	--4280
		x"00",	--4281
		x"4d",	--4282
		x"00",	--4283
		x"41",	--4284
		x"41",	--4285
		x"41",	--4286
		x"90",	--4287
		x"00",	--4288
		x"24",	--4289
		x"50",	--4290
		x"ff",	--4291
		x"4d",	--4292
		x"00",	--4293
		x"40",	--4294
		x"00",	--4295
		x"00",	--4296
		x"4a",	--4297
		x"4b",	--4298
		x"5c",	--4299
		x"6d",	--4300
		x"5c",	--4301
		x"6d",	--4302
		x"5c",	--4303
		x"6d",	--4304
		x"5c",	--4305
		x"6d",	--4306
		x"5c",	--4307
		x"6d",	--4308
		x"5c",	--4309
		x"6d",	--4310
		x"5c",	--4311
		x"6d",	--4312
		x"4c",	--4313
		x"4d",	--4314
		x"d3",	--4315
		x"d0",	--4316
		x"40",	--4317
		x"4a",	--4318
		x"00",	--4319
		x"4b",	--4320
		x"00",	--4321
		x"41",	--4322
		x"41",	--4323
		x"41",	--4324
		x"93",	--4325
		x"23",	--4326
		x"43",	--4327
		x"00",	--4328
		x"41",	--4329
		x"41",	--4330
		x"41",	--4331
		x"93",	--4332
		x"24",	--4333
		x"4a",	--4334
		x"4b",	--4335
		x"f3",	--4336
		x"f0",	--4337
		x"00",	--4338
		x"93",	--4339
		x"20",	--4340
		x"93",	--4341
		x"24",	--4342
		x"43",	--4343
		x"00",	--4344
		x"3f",	--4345
		x"93",	--4346
		x"23",	--4347
		x"42",	--4348
		x"00",	--4349
		x"3f",	--4350
		x"43",	--4351
		x"00",	--4352
		x"3f",	--4353
		x"12",	--4354
		x"4f",	--4355
		x"93",	--4356
		x"28",	--4357
		x"4e",	--4358
		x"93",	--4359
		x"28",	--4360
		x"92",	--4361
		x"24",	--4362
		x"92",	--4363
		x"24",	--4364
		x"93",	--4365
		x"24",	--4366
		x"93",	--4367
		x"24",	--4368
		x"4f",	--4369
		x"00",	--4370
		x"9e",	--4371
		x"00",	--4372
		x"24",	--4373
		x"93",	--4374
		x"20",	--4375
		x"43",	--4376
		x"4e",	--4377
		x"41",	--4378
		x"41",	--4379
		x"93",	--4380
		x"24",	--4381
		x"93",	--4382
		x"00",	--4383
		x"23",	--4384
		x"43",	--4385
		x"4e",	--4386
		x"41",	--4387
		x"41",	--4388
		x"93",	--4389
		x"00",	--4390
		x"27",	--4391
		x"43",	--4392
		x"3f",	--4393
		x"4f",	--4394
		x"00",	--4395
		x"4e",	--4396
		x"00",	--4397
		x"9b",	--4398
		x"3b",	--4399
		x"9c",	--4400
		x"38",	--4401
		x"4f",	--4402
		x"00",	--4403
		x"4f",	--4404
		x"00",	--4405
		x"4e",	--4406
		x"00",	--4407
		x"4e",	--4408
		x"00",	--4409
		x"9f",	--4410
		x"2b",	--4411
		x"9e",	--4412
		x"28",	--4413
		x"9b",	--4414
		x"2b",	--4415
		x"9e",	--4416
		x"28",	--4417
		x"9f",	--4418
		x"28",	--4419
		x"9c",	--4420
		x"28",	--4421
		x"43",	--4422
		x"3f",	--4423
		x"93",	--4424
		x"23",	--4425
		x"43",	--4426
		x"3f",	--4427
		x"92",	--4428
		x"23",	--4429
		x"4e",	--4430
		x"00",	--4431
		x"4f",	--4432
		x"00",	--4433
		x"8f",	--4434
		x"3f",	--4435
		x"42",	--4436
		x"02",	--4437
		x"93",	--4438
		x"38",	--4439
		x"42",	--4440
		x"02",	--4441
		x"4f",	--4442
		x"00",	--4443
		x"53",	--4444
		x"4d",	--4445
		x"02",	--4446
		x"53",	--4447
		x"4e",	--4448
		x"02",	--4449
		x"41",	--4450
		x"43",	--4451
		x"41",	--4452
		x"12",	--4453
		x"12",	--4454
		x"83",	--4455
		x"4e",	--4456
		x"00",	--4457
		x"42",	--4458
		x"02",	--4459
		x"42",	--4460
		x"02",	--4461
		x"4e",	--4462
		x"4f",	--4463
		x"40",	--4464
		x"e2",	--4465
		x"12",	--4466
		x"e4",	--4467
		x"9b",	--4468
		x"38",	--4469
		x"4a",	--4470
		x"5b",	--4471
		x"43",	--4472
		x"ff",	--4473
		x"3c",	--4474
		x"42",	--4475
		x"02",	--4476
		x"43",	--4477
		x"00",	--4478
		x"53",	--4479
		x"41",	--4480
		x"41",	--4481
		x"41",	--4482
		x"41",	--4483
		x"00",	--4484
		x"02",	--4485
		x"40",	--4486
		x"7f",	--4487
		x"02",	--4488
		x"41",	--4489
		x"50",	--4490
		x"00",	--4491
		x"41",	--4492
		x"00",	--4493
		x"12",	--4494
		x"e2",	--4495
		x"41",	--4496
		x"41",	--4497
		x"00",	--4498
		x"02",	--4499
		x"41",	--4500
		x"00",	--4501
		x"02",	--4502
		x"41",	--4503
		x"52",	--4504
		x"41",	--4505
		x"00",	--4506
		x"12",	--4507
		x"e2",	--4508
		x"41",	--4509
		x"4e",	--4510
		x"4f",	--4511
		x"02",	--4512
		x"40",	--4513
		x"7f",	--4514
		x"02",	--4515
		x"4d",	--4516
		x"4c",	--4517
		x"12",	--4518
		x"e2",	--4519
		x"41",	--4520
		x"4f",	--4521
		x"02",	--4522
		x"4e",	--4523
		x"02",	--4524
		x"4c",	--4525
		x"4d",	--4526
		x"12",	--4527
		x"e2",	--4528
		x"41",	--4529
		x"12",	--4530
		x"12",	--4531
		x"12",	--4532
		x"12",	--4533
		x"12",	--4534
		x"12",	--4535
		x"12",	--4536
		x"12",	--4537
		x"82",	--4538
		x"4f",	--4539
		x"4e",	--4540
		x"00",	--4541
		x"4d",	--4542
		x"41",	--4543
		x"00",	--4544
		x"41",	--4545
		x"00",	--4546
		x"4d",	--4547
		x"4d",	--4548
		x"10",	--4549
		x"44",	--4550
		x"4f",	--4551
		x"b0",	--4552
		x"00",	--4553
		x"24",	--4554
		x"40",	--4555
		x"00",	--4556
		x"00",	--4557
		x"4f",	--4558
		x"10",	--4559
		x"f3",	--4560
		x"24",	--4561
		x"40",	--4562
		x"00",	--4563
		x"3c",	--4564
		x"40",	--4565
		x"00",	--4566
		x"4e",	--4567
		x"00",	--4568
		x"41",	--4569
		x"53",	--4570
		x"3c",	--4571
		x"f0",	--4572
		x"00",	--4573
		x"24",	--4574
		x"40",	--4575
		x"00",	--4576
		x"00",	--4577
		x"3c",	--4578
		x"93",	--4579
		x"24",	--4580
		x"4d",	--4581
		x"00",	--4582
		x"41",	--4583
		x"53",	--4584
		x"3c",	--4585
		x"41",	--4586
		x"4c",	--4587
		x"10",	--4588
		x"11",	--4589
		x"10",	--4590
		x"11",	--4591
		x"4c",	--4592
		x"41",	--4593
		x"41",	--4594
		x"10",	--4595
		x"11",	--4596
		x"10",	--4597
		x"11",	--4598
		x"4c",	--4599
		x"86",	--4600
		x"77",	--4601
		x"4f",	--4602
		x"10",	--4603
		x"4e",	--4604
		x"00",	--4605
		x"f2",	--4606
		x"24",	--4607
		x"45",	--4608
		x"3c",	--4609
		x"43",	--4610
		x"4f",	--4611
		x"b0",	--4612
		x"00",	--4613
		x"20",	--4614
		x"41",	--4615
		x"00",	--4616
		x"53",	--4617
		x"53",	--4618
		x"93",	--4619
		x"00",	--4620
		x"23",	--4621
		x"81",	--4622
		x"00",	--4623
		x"9a",	--4624
		x"28",	--4625
		x"8a",	--4626
		x"3c",	--4627
		x"43",	--4628
		x"b3",	--4629
		x"00",	--4630
		x"24",	--4631
		x"95",	--4632
		x"28",	--4633
		x"85",	--4634
		x"3c",	--4635
		x"43",	--4636
		x"4d",	--4637
		x"9d",	--4638
		x"2c",	--4639
		x"47",	--4640
		x"93",	--4641
		x"38",	--4642
		x"40",	--4643
		x"00",	--4644
		x"00",	--4645
		x"43",	--4646
		x"43",	--4647
		x"3c",	--4648
		x"41",	--4649
		x"56",	--4650
		x"4f",	--4651
		x"11",	--4652
		x"53",	--4653
		x"12",	--4654
		x"3c",	--4655
		x"43",	--4656
		x"9a",	--4657
		x"3b",	--4658
		x"4a",	--4659
		x"40",	--4660
		x"00",	--4661
		x"00",	--4662
		x"8b",	--4663
		x"3c",	--4664
		x"41",	--4665
		x"00",	--4666
		x"11",	--4667
		x"12",	--4668
		x"53",	--4669
		x"45",	--4670
		x"5b",	--4671
		x"99",	--4672
		x"2b",	--4673
		x"3c",	--4674
		x"43",	--4675
		x"43",	--4676
		x"3c",	--4677
		x"53",	--4678
		x"41",	--4679
		x"56",	--4680
		x"4f",	--4681
		x"11",	--4682
		x"53",	--4683
		x"12",	--4684
		x"9a",	--4685
		x"3b",	--4686
		x"b3",	--4687
		x"00",	--4688
		x"24",	--4689
		x"44",	--4690
		x"3c",	--4691
		x"41",	--4692
		x"00",	--4693
		x"8b",	--4694
		x"3c",	--4695
		x"40",	--4696
		x"00",	--4697
		x"12",	--4698
		x"53",	--4699
		x"93",	--4700
		x"23",	--4701
		x"44",	--4702
		x"54",	--4703
		x"3f",	--4704
		x"53",	--4705
		x"11",	--4706
		x"12",	--4707
		x"53",	--4708
		x"4a",	--4709
		x"5b",	--4710
		x"4f",	--4711
		x"93",	--4712
		x"24",	--4713
		x"93",	--4714
		x"23",	--4715
		x"3c",	--4716
		x"40",	--4717
		x"00",	--4718
		x"12",	--4719
		x"53",	--4720
		x"99",	--4721
		x"2b",	--4722
		x"4b",	--4723
		x"52",	--4724
		x"41",	--4725
		x"41",	--4726
		x"41",	--4727
		x"41",	--4728
		x"41",	--4729
		x"41",	--4730
		x"41",	--4731
		x"41",	--4732
		x"41",	--4733
		x"12",	--4734
		x"12",	--4735
		x"12",	--4736
		x"12",	--4737
		x"12",	--4738
		x"12",	--4739
		x"12",	--4740
		x"12",	--4741
		x"50",	--4742
		x"ff",	--4743
		x"4f",	--4744
		x"00",	--4745
		x"4e",	--4746
		x"4d",	--4747
		x"4e",	--4748
		x"00",	--4749
		x"43",	--4750
		x"00",	--4751
		x"43",	--4752
		x"00",	--4753
		x"43",	--4754
		x"00",	--4755
		x"43",	--4756
		x"00",	--4757
		x"43",	--4758
		x"00",	--4759
		x"43",	--4760
		x"00",	--4761
		x"43",	--4762
		x"43",	--4763
		x"00",	--4764
		x"41",	--4765
		x"50",	--4766
		x"00",	--4767
		x"4e",	--4768
		x"00",	--4769
		x"40",	--4770
		x"eb",	--4771
		x"46",	--4772
		x"53",	--4773
		x"4f",	--4774
		x"00",	--4775
		x"93",	--4776
		x"20",	--4777
		x"90",	--4778
		x"00",	--4779
		x"20",	--4780
		x"43",	--4781
		x"00",	--4782
		x"43",	--4783
		x"00",	--4784
		x"46",	--4785
		x"00",	--4786
		x"43",	--4787
		x"00",	--4788
		x"43",	--4789
		x"00",	--4790
		x"43",	--4791
		x"00",	--4792
		x"43",	--4793
		x"00",	--4794
		x"43",	--4795
		x"00",	--4796
		x"40",	--4797
		x"eb",	--4798
		x"47",	--4799
		x"11",	--4800
		x"4e",	--4801
		x"12",	--4802
		x"00",	--4803
		x"53",	--4804
		x"00",	--4805
		x"40",	--4806
		x"eb",	--4807
		x"90",	--4808
		x"00",	--4809
		x"24",	--4810
		x"90",	--4811
		x"00",	--4812
		x"34",	--4813
		x"90",	--4814
		x"00",	--4815
		x"24",	--4816
		x"90",	--4817
		x"00",	--4818
		x"34",	--4819
		x"90",	--4820
		x"00",	--4821
		x"24",	--4822
		x"90",	--4823
		x"00",	--4824
		x"34",	--4825
		x"90",	--4826
		x"00",	--4827
		x"24",	--4828
		x"90",	--4829
		x"00",	--4830
		x"27",	--4831
		x"90",	--4832
		x"00",	--4833
		x"20",	--4834
		x"3c",	--4835
		x"90",	--4836
		x"00",	--4837
		x"24",	--4838
		x"90",	--4839
		x"00",	--4840
		x"24",	--4841
		x"90",	--4842
		x"00",	--4843
		x"20",	--4844
		x"3c",	--4845
		x"90",	--4846
		x"00",	--4847
		x"38",	--4848
		x"90",	--4849
		x"00",	--4850
		x"20",	--4851
		x"3c",	--4852
		x"90",	--4853
		x"00",	--4854
		x"24",	--4855
		x"90",	--4856
		x"00",	--4857
		x"34",	--4858
		x"90",	--4859
		x"00",	--4860
		x"24",	--4861
		x"90",	--4862
		x"00",	--4863
		x"24",	--4864
		x"90",	--4865
		x"00",	--4866
		x"20",	--4867
		x"3c",	--4868
		x"90",	--4869
		x"00",	--4870
		x"24",	--4871
		x"90",	--4872
		x"00",	--4873
		x"34",	--4874
		x"90",	--4875
		x"00",	--4876
		x"20",	--4877
		x"3c",	--4878
		x"90",	--4879
		x"00",	--4880
		x"24",	--4881
		x"90",	--4882
		x"00",	--4883
		x"24",	--4884
		x"41",	--4885
		x"00",	--4886
		x"41",	--4887
		x"00",	--4888
		x"89",	--4889
		x"40",	--4890
		x"eb",	--4891
		x"42",	--4892
		x"00",	--4893
		x"3c",	--4894
		x"d2",	--4895
		x"00",	--4896
		x"40",	--4897
		x"eb",	--4898
		x"41",	--4899
		x"f3",	--4900
		x"41",	--4901
		x"24",	--4902
		x"f0",	--4903
		x"ff",	--4904
		x"d3",	--4905
		x"3c",	--4906
		x"d3",	--4907
		x"4e",	--4908
		x"00",	--4909
		x"40",	--4910
		x"eb",	--4911
		x"d0",	--4912
		x"00",	--4913
		x"00",	--4914
		x"40",	--4915
		x"eb",	--4916
		x"40",	--4917
		x"00",	--4918
		x"00",	--4919
		x"40",	--4920
		x"eb",	--4921
		x"90",	--4922
		x"00",	--4923
		x"00",	--4924
		x"20",	--4925
		x"40",	--4926
		x"eb",	--4927
		x"40",	--4928
		x"00",	--4929
		x"00",	--4930
		x"40",	--4931
		x"eb",	--4932
		x"93",	--4933
		x"00",	--4934
		x"24",	--4935
		x"40",	--4936
		x"eb",	--4937
		x"43",	--4938
		x"00",	--4939
		x"40",	--4940
		x"eb",	--4941
		x"45",	--4942
		x"53",	--4943
		x"45",	--4944
		x"93",	--4945
		x"38",	--4946
		x"4a",	--4947
		x"00",	--4948
		x"3c",	--4949
		x"93",	--4950
		x"00",	--4951
		x"24",	--4952
		x"40",	--4953
		x"eb",	--4954
		x"d0",	--4955
		x"00",	--4956
		x"00",	--4957
		x"e3",	--4958
		x"4a",	--4959
		x"00",	--4960
		x"53",	--4961
		x"00",	--4962
		x"4e",	--4963
		x"3c",	--4964
		x"93",	--4965
		x"00",	--4966
		x"20",	--4967
		x"93",	--4968
		x"00",	--4969
		x"20",	--4970
		x"41",	--4971
		x"f0",	--4972
		x"00",	--4973
		x"43",	--4974
		x"24",	--4975
		x"43",	--4976
		x"4e",	--4977
		x"11",	--4978
		x"43",	--4979
		x"10",	--4980
		x"41",	--4981
		x"f0",	--4982
		x"00",	--4983
		x"de",	--4984
		x"4a",	--4985
		x"00",	--4986
		x"40",	--4987
		x"eb",	--4988
		x"41",	--4989
		x"00",	--4990
		x"5a",	--4991
		x"4a",	--4992
		x"5c",	--4993
		x"5c",	--4994
		x"5c",	--4995
		x"4a",	--4996
		x"00",	--4997
		x"50",	--4998
		x"ff",	--4999
		x"00",	--5000
		x"11",	--5001
		x"5e",	--5002
		x"00",	--5003
		x"43",	--5004
		x"00",	--5005
		x"40",	--5006
		x"eb",	--5007
		x"45",	--5008
		x"53",	--5009
		x"45",	--5010
		x"93",	--5011
		x"00",	--5012
		x"20",	--5013
		x"93",	--5014
		x"00",	--5015
		x"27",	--5016
		x"4e",	--5017
		x"00",	--5018
		x"43",	--5019
		x"00",	--5020
		x"41",	--5021
		x"52",	--5022
		x"3c",	--5023
		x"45",	--5024
		x"53",	--5025
		x"45",	--5026
		x"93",	--5027
		x"00",	--5028
		x"24",	--5029
		x"d2",	--5030
		x"00",	--5031
		x"41",	--5032
		x"00",	--5033
		x"4f",	--5034
		x"00",	--5035
		x"3c",	--5036
		x"93",	--5037
		x"00",	--5038
		x"24",	--5039
		x"41",	--5040
		x"00",	--5041
		x"00",	--5042
		x"93",	--5043
		x"20",	--5044
		x"40",	--5045
		x"f1",	--5046
		x"12",	--5047
		x"00",	--5048
		x"12",	--5049
		x"00",	--5050
		x"41",	--5051
		x"00",	--5052
		x"41",	--5053
		x"00",	--5054
		x"12",	--5055
		x"e3",	--5056
		x"52",	--5057
		x"5f",	--5058
		x"00",	--5059
		x"47",	--5060
		x"40",	--5061
		x"eb",	--5062
		x"45",	--5063
		x"53",	--5064
		x"45",	--5065
		x"49",	--5066
		x"00",	--5067
		x"43",	--5068
		x"93",	--5069
		x"20",	--5070
		x"43",	--5071
		x"5e",	--5072
		x"5e",	--5073
		x"5e",	--5074
		x"41",	--5075
		x"f0",	--5076
		x"ff",	--5077
		x"de",	--5078
		x"4a",	--5079
		x"00",	--5080
		x"47",	--5081
		x"40",	--5082
		x"00",	--5083
		x"00",	--5084
		x"3c",	--5085
		x"d3",	--5086
		x"00",	--5087
		x"3c",	--5088
		x"d2",	--5089
		x"00",	--5090
		x"40",	--5091
		x"00",	--5092
		x"00",	--5093
		x"3c",	--5094
		x"40",	--5095
		x"00",	--5096
		x"00",	--5097
		x"41",	--5098
		x"b3",	--5099
		x"24",	--5100
		x"45",	--5101
		x"52",	--5102
		x"45",	--5103
		x"45",	--5104
		x"00",	--5105
		x"45",	--5106
		x"00",	--5107
		x"45",	--5108
		x"00",	--5109
		x"48",	--5110
		x"00",	--5111
		x"47",	--5112
		x"00",	--5113
		x"46",	--5114
		x"00",	--5115
		x"4b",	--5116
		x"00",	--5117
		x"43",	--5118
		x"00",	--5119
		x"93",	--5120
		x"20",	--5121
		x"93",	--5122
		x"20",	--5123
		x"93",	--5124
		x"20",	--5125
		x"93",	--5126
		x"24",	--5127
		x"43",	--5128
		x"00",	--5129
		x"5b",	--5130
		x"43",	--5131
		x"6b",	--5132
		x"4b",	--5133
		x"00",	--5134
		x"4c",	--5135
		x"3c",	--5136
		x"f3",	--5137
		x"45",	--5138
		x"24",	--5139
		x"52",	--5140
		x"45",	--5141
		x"45",	--5142
		x"00",	--5143
		x"48",	--5144
		x"00",	--5145
		x"4b",	--5146
		x"00",	--5147
		x"43",	--5148
		x"00",	--5149
		x"93",	--5150
		x"20",	--5151
		x"3c",	--5152
		x"53",	--5153
		x"45",	--5154
		x"4b",	--5155
		x"00",	--5156
		x"43",	--5157
		x"00",	--5158
		x"93",	--5159
		x"24",	--5160
		x"43",	--5161
		x"00",	--5162
		x"5b",	--5163
		x"43",	--5164
		x"6b",	--5165
		x"4b",	--5166
		x"00",	--5167
		x"47",	--5168
		x"b2",	--5169
		x"00",	--5170
		x"24",	--5171
		x"93",	--5172
		x"00",	--5173
		x"20",	--5174
		x"41",	--5175
		x"90",	--5176
		x"00",	--5177
		x"00",	--5178
		x"20",	--5179
		x"d0",	--5180
		x"00",	--5181
		x"3c",	--5182
		x"92",	--5183
		x"00",	--5184
		x"20",	--5185
		x"d0",	--5186
		x"00",	--5187
		x"48",	--5188
		x"00",	--5189
		x"41",	--5190
		x"b2",	--5191
		x"24",	--5192
		x"93",	--5193
		x"00",	--5194
		x"24",	--5195
		x"40",	--5196
		x"00",	--5197
		x"00",	--5198
		x"b3",	--5199
		x"24",	--5200
		x"e3",	--5201
		x"00",	--5202
		x"e3",	--5203
		x"00",	--5204
		x"e3",	--5205
		x"00",	--5206
		x"e3",	--5207
		x"00",	--5208
		x"53",	--5209
		x"00",	--5210
		x"63",	--5211
		x"00",	--5212
		x"63",	--5213
		x"00",	--5214
		x"63",	--5215
		x"00",	--5216
		x"3c",	--5217
		x"b3",	--5218
		x"24",	--5219
		x"41",	--5220
		x"00",	--5221
		x"41",	--5222
		x"00",	--5223
		x"e3",	--5224
		x"e3",	--5225
		x"4a",	--5226
		x"4b",	--5227
		x"53",	--5228
		x"63",	--5229
		x"4e",	--5230
		x"00",	--5231
		x"4f",	--5232
		x"00",	--5233
		x"3c",	--5234
		x"41",	--5235
		x"00",	--5236
		x"e3",	--5237
		x"53",	--5238
		x"4a",	--5239
		x"00",	--5240
		x"43",	--5241
		x"00",	--5242
		x"b3",	--5243
		x"24",	--5244
		x"41",	--5245
		x"00",	--5246
		x"41",	--5247
		x"00",	--5248
		x"00",	--5249
		x"41",	--5250
		x"00",	--5251
		x"41",	--5252
		x"00",	--5253
		x"41",	--5254
		x"50",	--5255
		x"00",	--5256
		x"46",	--5257
		x"41",	--5258
		x"00",	--5259
		x"00",	--5260
		x"41",	--5261
		x"00",	--5262
		x"10",	--5263
		x"11",	--5264
		x"10",	--5265
		x"11",	--5266
		x"4b",	--5267
		x"00",	--5268
		x"4b",	--5269
		x"00",	--5270
		x"4b",	--5271
		x"00",	--5272
		x"12",	--5273
		x"00",	--5274
		x"12",	--5275
		x"00",	--5276
		x"12",	--5277
		x"00",	--5278
		x"12",	--5279
		x"00",	--5280
		x"49",	--5281
		x"41",	--5282
		x"00",	--5283
		x"48",	--5284
		x"44",	--5285
		x"12",	--5286
		x"ed",	--5287
		x"52",	--5288
		x"4c",	--5289
		x"90",	--5290
		x"00",	--5291
		x"34",	--5292
		x"50",	--5293
		x"00",	--5294
		x"4b",	--5295
		x"00",	--5296
		x"3c",	--5297
		x"4c",	--5298
		x"b3",	--5299
		x"00",	--5300
		x"24",	--5301
		x"40",	--5302
		x"00",	--5303
		x"3c",	--5304
		x"40",	--5305
		x"00",	--5306
		x"5b",	--5307
		x"4a",	--5308
		x"00",	--5309
		x"47",	--5310
		x"53",	--5311
		x"12",	--5312
		x"00",	--5313
		x"12",	--5314
		x"00",	--5315
		x"12",	--5316
		x"00",	--5317
		x"12",	--5318
		x"00",	--5319
		x"49",	--5320
		x"41",	--5321
		x"00",	--5322
		x"48",	--5323
		x"44",	--5324
		x"12",	--5325
		x"ec",	--5326
		x"52",	--5327
		x"4c",	--5328
		x"4d",	--5329
		x"00",	--5330
		x"4e",	--5331
		x"4f",	--5332
		x"53",	--5333
		x"93",	--5334
		x"23",	--5335
		x"93",	--5336
		x"23",	--5337
		x"93",	--5338
		x"23",	--5339
		x"93",	--5340
		x"23",	--5341
		x"43",	--5342
		x"00",	--5343
		x"43",	--5344
		x"00",	--5345
		x"43",	--5346
		x"00",	--5347
		x"43",	--5348
		x"00",	--5349
		x"3c",	--5350
		x"b3",	--5351
		x"24",	--5352
		x"41",	--5353
		x"00",	--5354
		x"41",	--5355
		x"00",	--5356
		x"41",	--5357
		x"50",	--5358
		x"00",	--5359
		x"41",	--5360
		x"00",	--5361
		x"10",	--5362
		x"11",	--5363
		x"10",	--5364
		x"11",	--5365
		x"41",	--5366
		x"00",	--5367
		x"49",	--5368
		x"44",	--5369
		x"47",	--5370
		x"12",	--5371
		x"ec",	--5372
		x"4e",	--5373
		x"90",	--5374
		x"00",	--5375
		x"34",	--5376
		x"50",	--5377
		x"00",	--5378
		x"4b",	--5379
		x"00",	--5380
		x"3c",	--5381
		x"4e",	--5382
		x"b3",	--5383
		x"00",	--5384
		x"24",	--5385
		x"40",	--5386
		x"00",	--5387
		x"3c",	--5388
		x"40",	--5389
		x"00",	--5390
		x"5b",	--5391
		x"4a",	--5392
		x"00",	--5393
		x"48",	--5394
		x"53",	--5395
		x"41",	--5396
		x"00",	--5397
		x"49",	--5398
		x"44",	--5399
		x"47",	--5400
		x"12",	--5401
		x"eb",	--5402
		x"4e",	--5403
		x"4f",	--5404
		x"53",	--5405
		x"93",	--5406
		x"23",	--5407
		x"93",	--5408
		x"23",	--5409
		x"43",	--5410
		x"00",	--5411
		x"43",	--5412
		x"00",	--5413
		x"3c",	--5414
		x"41",	--5415
		x"00",	--5416
		x"41",	--5417
		x"50",	--5418
		x"00",	--5419
		x"41",	--5420
		x"00",	--5421
		x"47",	--5422
		x"12",	--5423
		x"ec",	--5424
		x"4f",	--5425
		x"90",	--5426
		x"00",	--5427
		x"34",	--5428
		x"50",	--5429
		x"00",	--5430
		x"4d",	--5431
		x"00",	--5432
		x"3c",	--5433
		x"4f",	--5434
		x"b3",	--5435
		x"00",	--5436
		x"24",	--5437
		x"40",	--5438
		x"00",	--5439
		x"3c",	--5440
		x"40",	--5441
		x"00",	--5442
		x"5d",	--5443
		x"4c",	--5444
		x"00",	--5445
		x"48",	--5446
		x"53",	--5447
		x"41",	--5448
		x"00",	--5449
		x"47",	--5450
		x"12",	--5451
		x"ec",	--5452
		x"4f",	--5453
		x"53",	--5454
		x"93",	--5455
		x"23",	--5456
		x"43",	--5457
		x"00",	--5458
		x"90",	--5459
		x"00",	--5460
		x"00",	--5461
		x"24",	--5462
		x"43",	--5463
		x"00",	--5464
		x"93",	--5465
		x"00",	--5466
		x"24",	--5467
		x"41",	--5468
		x"50",	--5469
		x"00",	--5470
		x"4f",	--5471
		x"00",	--5472
		x"41",	--5473
		x"00",	--5474
		x"10",	--5475
		x"11",	--5476
		x"10",	--5477
		x"11",	--5478
		x"4a",	--5479
		x"00",	--5480
		x"46",	--5481
		x"00",	--5482
		x"46",	--5483
		x"10",	--5484
		x"11",	--5485
		x"10",	--5486
		x"11",	--5487
		x"4a",	--5488
		x"00",	--5489
		x"41",	--5490
		x"00",	--5491
		x"41",	--5492
		x"00",	--5493
		x"81",	--5494
		x"00",	--5495
		x"71",	--5496
		x"00",	--5497
		x"83",	--5498
		x"91",	--5499
		x"00",	--5500
		x"2c",	--5501
		x"d3",	--5502
		x"00",	--5503
		x"41",	--5504
		x"00",	--5505
		x"8c",	--5506
		x"4e",	--5507
		x"00",	--5508
		x"3c",	--5509
		x"93",	--5510
		x"00",	--5511
		x"24",	--5512
		x"41",	--5513
		x"00",	--5514
		x"00",	--5515
		x"12",	--5516
		x"00",	--5517
		x"12",	--5518
		x"00",	--5519
		x"41",	--5520
		x"00",	--5521
		x"46",	--5522
		x"53",	--5523
		x"41",	--5524
		x"00",	--5525
		x"12",	--5526
		x"e3",	--5527
		x"52",	--5528
		x"5f",	--5529
		x"00",	--5530
		x"3c",	--5531
		x"49",	--5532
		x"11",	--5533
		x"12",	--5534
		x"00",	--5535
		x"49",	--5536
		x"58",	--5537
		x"91",	--5538
		x"00",	--5539
		x"2b",	--5540
		x"49",	--5541
		x"00",	--5542
		x"4e",	--5543
		x"00",	--5544
		x"43",	--5545
		x"3c",	--5546
		x"41",	--5547
		x"00",	--5548
		x"00",	--5549
		x"43",	--5550
		x"00",	--5551
		x"43",	--5552
		x"00",	--5553
		x"3c",	--5554
		x"4e",	--5555
		x"43",	--5556
		x"00",	--5557
		x"43",	--5558
		x"00",	--5559
		x"43",	--5560
		x"41",	--5561
		x"00",	--5562
		x"46",	--5563
		x"93",	--5564
		x"24",	--5565
		x"40",	--5566
		x"e5",	--5567
		x"41",	--5568
		x"00",	--5569
		x"50",	--5570
		x"00",	--5571
		x"41",	--5572
		x"41",	--5573
		x"41",	--5574
		x"41",	--5575
		x"41",	--5576
		x"41",	--5577
		x"41",	--5578
		x"41",	--5579
		x"41",	--5580
		x"43",	--5581
		x"93",	--5582
		x"34",	--5583
		x"40",	--5584
		x"00",	--5585
		x"e3",	--5586
		x"53",	--5587
		x"93",	--5588
		x"34",	--5589
		x"e3",	--5590
		x"e3",	--5591
		x"53",	--5592
		x"12",	--5593
		x"12",	--5594
		x"ec",	--5595
		x"41",	--5596
		x"b3",	--5597
		x"24",	--5598
		x"e3",	--5599
		x"53",	--5600
		x"b3",	--5601
		x"24",	--5602
		x"e3",	--5603
		x"53",	--5604
		x"41",	--5605
		x"12",	--5606
		x"eb",	--5607
		x"4e",	--5608
		x"41",	--5609
		x"12",	--5610
		x"12",	--5611
		x"12",	--5612
		x"40",	--5613
		x"00",	--5614
		x"4c",	--5615
		x"4d",	--5616
		x"43",	--5617
		x"43",	--5618
		x"5e",	--5619
		x"6f",	--5620
		x"6c",	--5621
		x"6d",	--5622
		x"9b",	--5623
		x"28",	--5624
		x"20",	--5625
		x"9a",	--5626
		x"28",	--5627
		x"8a",	--5628
		x"7b",	--5629
		x"d3",	--5630
		x"83",	--5631
		x"23",	--5632
		x"41",	--5633
		x"41",	--5634
		x"41",	--5635
		x"41",	--5636
		x"12",	--5637
		x"eb",	--5638
		x"4c",	--5639
		x"4d",	--5640
		x"41",	--5641
		x"12",	--5642
		x"43",	--5643
		x"93",	--5644
		x"34",	--5645
		x"40",	--5646
		x"00",	--5647
		x"e3",	--5648
		x"e3",	--5649
		x"53",	--5650
		x"63",	--5651
		x"93",	--5652
		x"34",	--5653
		x"e3",	--5654
		x"e3",	--5655
		x"e3",	--5656
		x"53",	--5657
		x"63",	--5658
		x"12",	--5659
		x"eb",	--5660
		x"b3",	--5661
		x"24",	--5662
		x"e3",	--5663
		x"e3",	--5664
		x"53",	--5665
		x"63",	--5666
		x"b3",	--5667
		x"24",	--5668
		x"e3",	--5669
		x"e3",	--5670
		x"53",	--5671
		x"63",	--5672
		x"41",	--5673
		x"41",	--5674
		x"12",	--5675
		x"ec",	--5676
		x"4c",	--5677
		x"4d",	--5678
		x"41",	--5679
		x"40",	--5680
		x"00",	--5681
		x"4e",	--5682
		x"43",	--5683
		x"5f",	--5684
		x"6e",	--5685
		x"9d",	--5686
		x"28",	--5687
		x"8d",	--5688
		x"d3",	--5689
		x"83",	--5690
		x"23",	--5691
		x"41",	--5692
		x"12",	--5693
		x"ec",	--5694
		x"4e",	--5695
		x"41",	--5696
		x"12",	--5697
		x"12",	--5698
		x"12",	--5699
		x"12",	--5700
		x"12",	--5701
		x"00",	--5702
		x"48",	--5703
		x"49",	--5704
		x"4a",	--5705
		x"4b",	--5706
		x"43",	--5707
		x"43",	--5708
		x"43",	--5709
		x"43",	--5710
		x"5c",	--5711
		x"6d",	--5712
		x"6e",	--5713
		x"6f",	--5714
		x"68",	--5715
		x"69",	--5716
		x"6a",	--5717
		x"6b",	--5718
		x"97",	--5719
		x"28",	--5720
		x"20",	--5721
		x"96",	--5722
		x"28",	--5723
		x"20",	--5724
		x"95",	--5725
		x"28",	--5726
		x"20",	--5727
		x"94",	--5728
		x"28",	--5729
		x"84",	--5730
		x"75",	--5731
		x"76",	--5732
		x"77",	--5733
		x"d3",	--5734
		x"83",	--5735
		x"00",	--5736
		x"23",	--5737
		x"53",	--5738
		x"41",	--5739
		x"41",	--5740
		x"41",	--5741
		x"41",	--5742
		x"41",	--5743
		x"12",	--5744
		x"12",	--5745
		x"12",	--5746
		x"12",	--5747
		x"41",	--5748
		x"00",	--5749
		x"41",	--5750
		x"00",	--5751
		x"41",	--5752
		x"00",	--5753
		x"41",	--5754
		x"00",	--5755
		x"12",	--5756
		x"ec",	--5757
		x"41",	--5758
		x"41",	--5759
		x"41",	--5760
		x"41",	--5761
		x"41",	--5762
		x"12",	--5763
		x"12",	--5764
		x"12",	--5765
		x"12",	--5766
		x"41",	--5767
		x"00",	--5768
		x"41",	--5769
		x"00",	--5770
		x"41",	--5771
		x"00",	--5772
		x"41",	--5773
		x"00",	--5774
		x"12",	--5775
		x"ec",	--5776
		x"48",	--5777
		x"49",	--5778
		x"4a",	--5779
		x"4b",	--5780
		x"41",	--5781
		x"41",	--5782
		x"41",	--5783
		x"41",	--5784
		x"41",	--5785
		x"12",	--5786
		x"12",	--5787
		x"12",	--5788
		x"12",	--5789
		x"12",	--5790
		x"41",	--5791
		x"00",	--5792
		x"41",	--5793
		x"00",	--5794
		x"41",	--5795
		x"00",	--5796
		x"41",	--5797
		x"00",	--5798
		x"12",	--5799
		x"ec",	--5800
		x"41",	--5801
		x"00",	--5802
		x"48",	--5803
		x"00",	--5804
		x"49",	--5805
		x"00",	--5806
		x"4a",	--5807
		x"00",	--5808
		x"4b",	--5809
		x"00",	--5810
		x"41",	--5811
		x"41",	--5812
		x"41",	--5813
		x"41",	--5814
		x"41",	--5815
		x"41",	--5816
		x"13",	--5817
		x"d0",	--5818
		x"00",	--5819
		x"3f",	--5820
		x"74",	--5821
		x"70",	--5822
		x"0a",	--5823
		x"63",	--5824
		x"72",	--5825
		x"65",	--5826
		x"74",	--5827
		x"75",	--5828
		x"61",	--5829
		x"65",	--5830
		x"0d",	--5831
		x"00",	--5832
		x"25",	--5833
		x"20",	--5834
		x"45",	--5835
		x"54",	--5836
		x"52",	--5837
		x"47",	--5838
		x"54",	--5839
		x"3c",	--5840
		x"49",	--5841
		x"45",	--5842
		x"55",	--5843
		x"3e",	--5844
		x"0a",	--5845
		x"25",	--5846
		x"20",	--5847
		x"64",	--5848
		x"0a",	--5849
		x"4e",	--5850
		x"74",	--5851
		x"69",	--5852
		x"70",	--5853
		x"65",	--5854
		x"65",	--5855
		x"74",	--5856
		x"64",	--5857
		x"59",	--5858
		x"74",	--5859
		x"0a",	--5860
		x"57",	--5861
		x"69",	--5862
		x"69",	--5863
		x"67",	--5864
		x"66",	--5865
		x"72",	--5866
		x"61",	--5867
		x"6e",	--5868
		x"77",	--5869
		x"2e",	--5870
		x"69",	--5871
		x"20",	--5872
		x"69",	--5873
		x"65",	--5874
		x"0a",	--5875
		x"57",	--5876
		x"20",	--5877
		x"68",	--5878
		x"75",	--5879
		x"64",	--5880
		x"6e",	--5881
		x"74",	--5882
		x"73",	--5883
		x"65",	--5884
		x"74",	--5885
		x"61",	--5886
		x"0d",	--5887
		x"00",	--5888
		x"74",	--5889
		x"70",	--5890
		x"0a",	--5891
		x"65",	--5892
		x"72",	--5893
		x"72",	--5894
		x"20",	--5895
		x"69",	--5896
		x"73",	--5897
		x"6e",	--5898
		x"20",	--5899
		x"72",	--5900
		x"75",	--5901
		x"65",	--5902
		x"74",	--5903
		x"0a",	--5904
		x"63",	--5905
		x"72",	--5906
		x"65",	--5907
		x"74",	--5908
		x"75",	--5909
		x"61",	--5910
		x"65",	--5911
		x"0d",	--5912
		x"00",	--5913
		x"25",	--5914
		x"20",	--5915
		x"45",	--5916
		x"54",	--5917
		x"52",	--5918
		x"47",	--5919
		x"54",	--5920
		x"3c",	--5921
		x"49",	--5922
		x"45",	--5923
		x"55",	--5924
		x"3e",	--5925
		x"0a",	--5926
		x"25",	--5927
		x"20",	--5928
		x"64",	--5929
		x"0a",	--5930
		x"25",	--5931
		x"64",	--5932
		x"25",	--5933
		x"64",	--5934
		x"25",	--5935
		x"0d",	--5936
		x"00",	--5937
		x"64",	--5938
		x"25",	--5939
		x"0d",	--5940
		x"00",	--5941
		x"c9",	--5942
		x"c9",	--5943
		x"c9",	--5944
		x"c9",	--5945
		x"c9",	--5946
		x"c9",	--5947
		x"c9",	--5948
		x"c9",	--5949
		x"0a",	--5950
		x"3d",	--5951
		x"3d",	--5952
		x"3d",	--5953
		x"4d",	--5954
		x"72",	--5955
		x"65",	--5956
		x"20",	--5957
		x"43",	--5958
		x"20",	--5959
		x"3d",	--5960
		x"3d",	--5961
		x"3d",	--5962
		x"0a",	--5963
		x"69",	--5964
		x"74",	--5965
		x"72",	--5966
		x"63",	--5967
		x"69",	--5968
		x"65",	--5969
		x"6d",	--5970
		x"64",	--5971
		x"00",	--5972
		x"72",	--5973
		x"74",	--5974
		x"00",	--5975
		x"65",	--5976
		x"64",	--5977
		x"62",	--5978
		x"7a",	--5979
		x"65",	--5980
		x"00",	--5981
		x"77",	--5982
		x"00",	--5983
		x"6e",	--5984
		x"6f",	--5985
		x"65",	--5986
		x"00",	--5987
		x"70",	--5988
		x"65",	--5989
		x"20",	--5990
		x"6f",	--5991
		x"74",	--5992
		x"6f",	--5993
		x"6c",	--5994
		x"72",	--5995
		x"73",	--5996
		x"65",	--5997
		x"64",	--5998
		x"63",	--5999
		x"6e",	--6000
		x"69",	--6001
		x"75",	--6002
		x"61",	--6003
		x"69",	--6004
		x"6e",	--6005
		x"62",	--6006
		x"6f",	--6007
		x"6c",	--6008
		x"61",	--6009
		x"65",	--6010
		x"00",	--6011
		x"0a",	--6012
		x"08",	--6013
		x"08",	--6014
		x"25",	--6015
		x"00",	--6016
		x"50",	--6017
		x"0a",	--6018
		x"44",	--6019
		x"57",	--6020
		x"0d",	--6021
		x"00",	--6022
		x"49",	--6023
		x"48",	--6024
		x"0d",	--6025
		x"00",	--6026
		x"45",	--6027
		x"54",	--6028
		x"0a",	--6029
		x"00",	--6030
		x"72",	--6031
		x"74",	--6032
		x"0a",	--6033
		x"00",	--6034
		x"72",	--6035
		x"6f",	--6036
		x"3a",	--6037
		x"6d",	--6038
		x"73",	--6039
		x"69",	--6040
		x"67",	--6041
		x"61",	--6042
		x"67",	--6043
		x"6d",	--6044
		x"6e",	--6045
		x"0d",	--6046
		x"00",	--6047
		x"6f",	--6048
		x"72",	--6049
		x"63",	--6050
		x"20",	--6051
		x"73",	--6052
		x"67",	--6053
		x"3a",	--6054
		x"0a",	--6055
		x"09",	--6056
		x"73",	--6057
		x"52",	--6058
		x"47",	--6059
		x"53",	--6060
		x"45",	--6061
		x"20",	--6062
		x"41",	--6063
		x"55",	--6064
		x"0d",	--6065
		x"00",	--6066
		x"3d",	--6067
		x"64",	--6068
		x"76",	--6069
		x"25",	--6070
		x"0d",	--6071
		x"00",	--6072
		x"25",	--6073
		x"20",	--6074
		x"45",	--6075
		x"49",	--6076
		x"54",	--6077
		x"52",	--6078
		x"0a",	--6079
		x"72",	--6080
		x"61",	--6081
		x"0a",	--6082
		x"00",	--6083
		x"63",	--6084
		x"69",	--6085
		x"20",	--6086
		x"6f",	--6087
		x"20",	--6088
		x"20",	--6089
		x"75",	--6090
		x"62",	--6091
		x"72",	--6092
		x"0a",	--6093
		x"25",	--6094
		x"20",	--6095
		x"73",	--6096
		x"0a",	--6097
		x"25",	--6098
		x"3a",	--6099
		x"6e",	--6100
		x"20",	--6101
		x"75",	--6102
		x"68",	--6103
		x"63",	--6104
		x"6d",	--6105
		x"61",	--6106
		x"64",	--6107
		x"0a",	--6108
		x"00",	--6109
		x"d3",	--6110
		x"d3",	--6111
		x"d3",	--6112
		x"d3",	--6113
		x"d3",	--6114
		x"d3",	--6115
		x"d3",	--6116
		x"d3",	--6117
		x"d3",	--6118
		x"d3",	--6119
		x"d3",	--6120
		x"d3",	--6121
		x"d3",	--6122
		x"d3",	--6123
		x"d3",	--6124
		x"d3",	--6125
		x"d3",	--6126
		x"d3",	--6127
		x"d3",	--6128
		x"d3",	--6129
		x"d3",	--6130
		x"d3",	--6131
		x"d3",	--6132
		x"d3",	--6133
		x"d3",	--6134
		x"d3",	--6135
		x"d3",	--6136
		x"d3",	--6137
		x"d3",	--6138
		x"d3",	--6139
		x"d3",	--6140
		x"d3",	--6141
		x"d3",	--6142
		x"d3",	--6143
		x"d3",	--6144
		x"d3",	--6145
		x"d3",	--6146
		x"d3",	--6147
		x"d3",	--6148
		x"d3",	--6149
		x"d3",	--6150
		x"d3",	--6151
		x"d3",	--6152
		x"d3",	--6153
		x"d3",	--6154
		x"d3",	--6155
		x"d3",	--6156
		x"d3",	--6157
		x"d3",	--6158
		x"d3",	--6159
		x"d3",	--6160
		x"d3",	--6161
		x"d3",	--6162
		x"d3",	--6163
		x"d3",	--6164
		x"d3",	--6165
		x"d3",	--6166
		x"d3",	--6167
		x"d3",	--6168
		x"d3",	--6169
		x"d3",	--6170
		x"d3",	--6171
		x"d3",	--6172
		x"d3",	--6173
		x"d3",	--6174
		x"d3",	--6175
		x"d3",	--6176
		x"d3",	--6177
		x"d3",	--6178
		x"d3",	--6179
		x"d3",	--6180
		x"d3",	--6181
		x"d3",	--6182
		x"d3",	--6183
		x"d3",	--6184
		x"d3",	--6185
		x"d3",	--6186
		x"d3",	--6187
		x"d3",	--6188
		x"d3",	--6189
		x"d3",	--6190
		x"d3",	--6191
		x"d3",	--6192
		x"d3",	--6193
		x"31",	--6194
		x"33",	--6195
		x"35",	--6196
		x"37",	--6197
		x"39",	--6198
		x"62",	--6199
		x"64",	--6200
		x"66",	--6201
		x"00",	--6202
		x"00",	--6203
		x"00",	--6204
		x"00",	--6205
		x"00",	--6206
		x"01",	--6207
		x"02",	--6208
		x"03",	--6209
		x"03",	--6210
		x"04",	--6211
		x"04",	--6212
		x"04",	--6213
		x"04",	--6214
		x"05",	--6215
		x"05",	--6216
		x"05",	--6217
		x"05",	--6218
		x"05",	--6219
		x"05",	--6220
		x"05",	--6221
		x"05",	--6222
		x"06",	--6223
		x"06",	--6224
		x"06",	--6225
		x"06",	--6226
		x"06",	--6227
		x"06",	--6228
		x"06",	--6229
		x"06",	--6230
		x"06",	--6231
		x"06",	--6232
		x"06",	--6233
		x"06",	--6234
		x"06",	--6235
		x"06",	--6236
		x"06",	--6237
		x"06",	--6238
		x"07",	--6239
		x"07",	--6240
		x"07",	--6241
		x"07",	--6242
		x"07",	--6243
		x"07",	--6244
		x"07",	--6245
		x"07",	--6246
		x"07",	--6247
		x"07",	--6248
		x"07",	--6249
		x"07",	--6250
		x"07",	--6251
		x"07",	--6252
		x"07",	--6253
		x"07",	--6254
		x"07",	--6255
		x"07",	--6256
		x"07",	--6257
		x"07",	--6258
		x"07",	--6259
		x"07",	--6260
		x"07",	--6261
		x"07",	--6262
		x"07",	--6263
		x"07",	--6264
		x"07",	--6265
		x"07",	--6266
		x"07",	--6267
		x"07",	--6268
		x"07",	--6269
		x"07",	--6270
		x"08",	--6271
		x"08",	--6272
		x"08",	--6273
		x"08",	--6274
		x"08",	--6275
		x"08",	--6276
		x"08",	--6277
		x"08",	--6278
		x"08",	--6279
		x"08",	--6280
		x"08",	--6281
		x"08",	--6282
		x"08",	--6283
		x"08",	--6284
		x"08",	--6285
		x"08",	--6286
		x"08",	--6287
		x"08",	--6288
		x"08",	--6289
		x"08",	--6290
		x"08",	--6291
		x"08",	--6292
		x"08",	--6293
		x"08",	--6294
		x"08",	--6295
		x"08",	--6296
		x"08",	--6297
		x"08",	--6298
		x"08",	--6299
		x"08",	--6300
		x"08",	--6301
		x"08",	--6302
		x"08",	--6303
		x"08",	--6304
		x"08",	--6305
		x"08",	--6306
		x"08",	--6307
		x"08",	--6308
		x"08",	--6309
		x"08",	--6310
		x"08",	--6311
		x"08",	--6312
		x"08",	--6313
		x"08",	--6314
		x"08",	--6315
		x"08",	--6316
		x"08",	--6317
		x"08",	--6318
		x"08",	--6319
		x"08",	--6320
		x"08",	--6321
		x"08",	--6322
		x"08",	--6323
		x"08",	--6324
		x"08",	--6325
		x"08",	--6326
		x"08",	--6327
		x"08",	--6328
		x"08",	--6329
		x"08",	--6330
		x"08",	--6331
		x"08",	--6332
		x"08",	--6333
		x"08",	--6334
		x"6e",	--6335
		x"6c",	--6336
		x"29",	--6337
		x"00",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"65",	--6342
		x"70",	--6343
		x"00",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"c3",	--8176
		x"c3",	--8177
		x"c3",	--8178
		x"c3",	--8179
		x"c3",	--8180
		x"c3",	--8181
		x"c3",	--8182
		x"d3",	--8183
		x"d0",	--8184
		x"c3",	--8185
		x"c3",	--8186
		x"c3",	--8187
		x"c3",	--8188
		x"c3",	--8189
		x"c3",	--8190
		x"c0");	--8191

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
