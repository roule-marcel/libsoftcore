library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"4c",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"10",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"4c",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"4e",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"3c",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"4c",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"10",	--29
		x"f9",	--30
		x"31",	--31
		x"3e",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"76",	--44
		x"b0",	--45
		x"b2",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"8a",	--50
		x"b0",	--51
		x"3a",	--52
		x"21",	--53
		x"3d",	--54
		x"a7",	--55
		x"3e",	--56
		x"8a",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"e2",	--61
		x"3d",	--62
		x"b8",	--63
		x"3e",	--64
		x"f4",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"e2",	--69
		x"3d",	--70
		x"be",	--71
		x"3e",	--72
		x"68",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"e2",	--77
		x"3d",	--78
		x"c3",	--79
		x"3e",	--80
		x"36",	--81
		x"7f",	--82
		x"61",	--83
		x"b0",	--84
		x"e2",	--85
		x"3d",	--86
		x"ca",	--87
		x"3e",	--88
		x"98",	--89
		x"7f",	--90
		x"70",	--91
		x"b0",	--92
		x"e2",	--93
		x"3d",	--94
		x"ce",	--95
		x"3e",	--96
		x"d8",	--97
		x"7f",	--98
		x"65",	--99
		x"b0",	--100
		x"e2",	--101
		x"3d",	--102
		x"d6",	--103
		x"3e",	--104
		x"68",	--105
		x"7f",	--106
		x"73",	--107
		x"b0",	--108
		x"e2",	--109
		x"3d",	--110
		x"e7",	--111
		x"3e",	--112
		x"06",	--113
		x"7f",	--114
		x"7a",	--115
		x"b0",	--116
		x"e2",	--117
		x"3d",	--118
		x"f0",	--119
		x"3e",	--120
		x"90",	--121
		x"7f",	--122
		x"63",	--123
		x"b0",	--124
		x"e2",	--125
		x"3d",	--126
		x"04",	--127
		x"3e",	--128
		x"c2",	--129
		x"7f",	--130
		x"6f",	--131
		x"b0",	--132
		x"e2",	--133
		x"3d",	--134
		x"17",	--135
		x"3e",	--136
		x"9a",	--137
		x"7f",	--138
		x"74",	--139
		x"b0",	--140
		x"e2",	--141
		x"3d",	--142
		x"1c",	--143
		x"3e",	--144
		x"9e",	--145
		x"7f",	--146
		x"62",	--147
		x"b0",	--148
		x"e2",	--149
		x"0e",	--150
		x"0f",	--151
		x"b0",	--152
		x"78",	--153
		x"2c",	--154
		x"3d",	--155
		x"20",	--156
		x"3e",	--157
		x"80",	--158
		x"0f",	--159
		x"3f",	--160
		x"12",	--161
		x"b0",	--162
		x"80",	--163
		x"0f",	--164
		x"3f",	--165
		x"12",	--166
		x"b0",	--167
		x"c8",	--168
		x"2c",	--169
		x"3d",	--170
		x"20",	--171
		x"3e",	--172
		x"88",	--173
		x"0f",	--174
		x"3f",	--175
		x"b0",	--176
		x"80",	--177
		x"0f",	--178
		x"3f",	--179
		x"b0",	--180
		x"c8",	--181
		x"0e",	--182
		x"3e",	--183
		x"0f",	--184
		x"3f",	--185
		x"12",	--186
		x"b0",	--187
		x"8e",	--188
		x"3e",	--189
		x"98",	--190
		x"0f",	--191
		x"3f",	--192
		x"06",	--193
		x"b0",	--194
		x"1c",	--195
		x"3e",	--196
		x"9c",	--197
		x"0f",	--198
		x"2f",	--199
		x"b0",	--200
		x"1c",	--201
		x"0e",	--202
		x"2e",	--203
		x"0f",	--204
		x"3f",	--205
		x"06",	--206
		x"b0",	--207
		x"c4",	--208
		x"0e",	--209
		x"3e",	--210
		x"0f",	--211
		x"3f",	--212
		x"12",	--213
		x"b0",	--214
		x"ce",	--215
		x"b0",	--216
		x"f4",	--217
		x"3e",	--218
		x"a0",	--219
		x"0f",	--220
		x"2f",	--221
		x"b0",	--222
		x"34",	--223
		x"0f",	--224
		x"2f",	--225
		x"b0",	--226
		x"30",	--227
		x"3d",	--228
		x"64",	--229
		x"3e",	--230
		x"2a",	--231
		x"0f",	--232
		x"2f",	--233
		x"b0",	--234
		x"48",	--235
		x"3e",	--236
		x"b0",	--237
		x"0f",	--238
		x"b0",	--239
		x"ae",	--240
		x"0f",	--241
		x"b0",	--242
		x"bc",	--243
		x"30",	--244
		x"a0",	--245
		x"03",	--246
		x"03",	--247
		x"03",	--248
		x"30",	--249
		x"d1",	--250
		x"30",	--251
		x"17",	--252
		x"30",	--253
		x"1d",	--254
		x"30",	--255
		x"52",	--256
		x"3c",	--257
		x"32",	--258
		x"0d",	--259
		x"3d",	--260
		x"16",	--261
		x"0e",	--262
		x"3e",	--263
		x"22",	--264
		x"0f",	--265
		x"3f",	--266
		x"a4",	--267
		x"b0",	--268
		x"a6",	--269
		x"31",	--270
		x"10",	--271
		x"30",	--272
		x"a0",	--273
		x"03",	--274
		x"03",	--275
		x"03",	--276
		x"30",	--277
		x"d1",	--278
		x"30",	--279
		x"17",	--280
		x"30",	--281
		x"1d",	--282
		x"30",	--283
		x"52",	--284
		x"3c",	--285
		x"32",	--286
		x"0d",	--287
		x"3d",	--288
		x"14",	--289
		x"0e",	--290
		x"3e",	--291
		x"18",	--292
		x"0f",	--293
		x"3f",	--294
		x"78",	--295
		x"b0",	--296
		x"a6",	--297
		x"31",	--298
		x"10",	--299
		x"0e",	--300
		x"3e",	--301
		x"68",	--302
		x"0f",	--303
		x"3f",	--304
		x"94",	--305
		x"b0",	--306
		x"58",	--307
		x"0f",	--308
		x"b0",	--309
		x"62",	--310
		x"b0",	--311
		x"30",	--312
		x"30",	--313
		x"b0",	--314
		x"30",	--315
		x"19",	--316
		x"30",	--317
		x"9a",	--318
		x"3d",	--319
		x"8f",	--320
		x"3e",	--321
		x"75",	--322
		x"0f",	--323
		x"3f",	--324
		x"22",	--325
		x"b0",	--326
		x"4e",	--327
		x"31",	--328
		x"06",	--329
		x"0d",	--330
		x"3d",	--331
		x"06",	--332
		x"0e",	--333
		x"2e",	--334
		x"0f",	--335
		x"3f",	--336
		x"1c",	--337
		x"b0",	--338
		x"a6",	--339
		x"3e",	--340
		x"64",	--341
		x"0f",	--342
		x"3f",	--343
		x"1c",	--344
		x"b0",	--345
		x"6a",	--346
		x"0f",	--347
		x"3f",	--348
		x"1c",	--349
		x"b0",	--350
		x"00",	--351
		x"0e",	--352
		x"3e",	--353
		x"68",	--354
		x"0f",	--355
		x"3f",	--356
		x"94",	--357
		x"b0",	--358
		x"6c",	--359
		x"0f",	--360
		x"b0",	--361
		x"76",	--362
		x"3f",	--363
		x"64",	--364
		x"b0",	--365
		x"7c",	--366
		x"f2",	--367
		x"80",	--368
		x"19",	--369
		x"32",	--370
		x"0b",	--371
		x"0a",	--372
		x"05",	--373
		x"1b",	--374
		x"03",	--375
		x"2b",	--376
		x"01",	--377
		x"0b",	--378
		x"b0",	--379
		x"94",	--380
		x"0f",	--381
		x"fc",	--382
		x"b0",	--383
		x"bc",	--384
		x"0b",	--385
		x"3e",	--386
		x"7f",	--387
		x"0d",	--388
		x"06",	--389
		x"7f",	--390
		x"1b",	--391
		x"ed",	--392
		x"7f",	--393
		x"1c",	--394
		x"12",	--395
		x"30",	--396
		x"27",	--397
		x"b0",	--398
		x"3a",	--399
		x"21",	--400
		x"3f",	--401
		x"40",	--402
		x"0f",	--403
		x"0a",	--404
		x"ca",	--405
		x"00",	--406
		x"0e",	--407
		x"5f",	--408
		x"40",	--409
		x"b0",	--410
		x"16",	--411
		x"0a",	--412
		x"dd",	--413
		x"0a",	--414
		x"db",	--415
		x"3a",	--416
		x"30",	--417
		x"2a",	--418
		x"b0",	--419
		x"3a",	--420
		x"21",	--421
		x"d4",	--422
		x"3a",	--423
		x"28",	--424
		x"d1",	--425
		x"82",	--426
		x"18",	--427
		x"0c",	--428
		x"4e",	--429
		x"8e",	--430
		x"0e",	--431
		x"30",	--432
		x"2e",	--433
		x"81",	--434
		x"c4",	--435
		x"b0",	--436
		x"3a",	--437
		x"21",	--438
		x"1f",	--439
		x"c0",	--440
		x"3e",	--441
		x"40",	--442
		x"0e",	--443
		x"0e",	--444
		x"ce",	--445
		x"00",	--446
		x"1a",	--447
		x"ba",	--448
		x"1b",	--449
		x"04",	--450
		x"7f",	--451
		x"5b",	--452
		x"b5",	--453
		x"b1",	--454
		x"2b",	--455
		x"b2",	--456
		x"7f",	--457
		x"42",	--458
		x"17",	--459
		x"7f",	--460
		x"43",	--461
		x"04",	--462
		x"7f",	--463
		x"41",	--464
		x"a8",	--465
		x"07",	--466
		x"7f",	--467
		x"43",	--468
		x"16",	--469
		x"7f",	--470
		x"44",	--471
		x"a1",	--472
		x"1b",	--473
		x"30",	--474
		x"31",	--475
		x"b0",	--476
		x"3a",	--477
		x"21",	--478
		x"b0",	--479
		x"f0",	--480
		x"0b",	--481
		x"98",	--482
		x"30",	--483
		x"36",	--484
		x"b0",	--485
		x"3a",	--486
		x"21",	--487
		x"b0",	--488
		x"18",	--489
		x"0b",	--490
		x"8f",	--491
		x"30",	--492
		x"3d",	--493
		x"b0",	--494
		x"3a",	--495
		x"21",	--496
		x"b0",	--497
		x"40",	--498
		x"0b",	--499
		x"86",	--500
		x"30",	--501
		x"45",	--502
		x"b0",	--503
		x"3a",	--504
		x"21",	--505
		x"b0",	--506
		x"68",	--507
		x"0b",	--508
		x"7d",	--509
		x"30",	--510
		x"56",	--511
		x"82",	--512
		x"10",	--513
		x"30",	--514
		x"0b",	--515
		x"30",	--516
		x"5e",	--517
		x"b0",	--518
		x"3a",	--519
		x"21",	--520
		x"1b",	--521
		x"10",	--522
		x"0c",	--523
		x"3d",	--524
		x"7a",	--525
		x"1e",	--526
		x"12",	--527
		x"1f",	--528
		x"14",	--529
		x"b0",	--530
		x"58",	--531
		x"b0",	--532
		x"02",	--533
		x"0e",	--534
		x"0c",	--535
		x"3d",	--536
		x"7a",	--537
		x"1e",	--538
		x"0e",	--539
		x"1f",	--540
		x"10",	--541
		x"b0",	--542
		x"58",	--543
		x"b0",	--544
		x"02",	--545
		x"0e",	--546
		x"0c",	--547
		x"3d",	--548
		x"7a",	--549
		x"1e",	--550
		x"0a",	--551
		x"1f",	--552
		x"0c",	--553
		x"b0",	--554
		x"58",	--555
		x"b0",	--556
		x"02",	--557
		x"0e",	--558
		x"30",	--559
		x"61",	--560
		x"30",	--561
		x"4c",	--562
		x"b0",	--563
		x"ea",	--564
		x"31",	--565
		x"0a",	--566
		x"30",	--567
		x"4c",	--568
		x"30",	--569
		x"6a",	--570
		x"b0",	--571
		x"3a",	--572
		x"21",	--573
		x"0f",	--574
		x"3b",	--575
		x"30",	--576
		x"0b",	--577
		x"30",	--578
		x"6f",	--579
		x"b0",	--580
		x"3a",	--581
		x"21",	--582
		x"0b",	--583
		x"0e",	--584
		x"1f",	--585
		x"12",	--586
		x"b0",	--587
		x"be",	--588
		x"0f",	--589
		x"30",	--590
		x"72",	--591
		x"b0",	--592
		x"3a",	--593
		x"21",	--594
		x"1b",	--595
		x"3b",	--596
		x"05",	--597
		x"f1",	--598
		x"30",	--599
		x"76",	--600
		x"b0",	--601
		x"3a",	--602
		x"21",	--603
		x"3b",	--604
		x"30",	--605
		x"82",	--606
		x"12",	--607
		x"30",	--608
		x"0b",	--609
		x"21",	--610
		x"0b",	--611
		x"81",	--612
		x"00",	--613
		x"1f",	--614
		x"14",	--615
		x"b2",	--616
		x"00",	--617
		x"25",	--618
		x"92",	--619
		x"14",	--620
		x"0e",	--621
		x"1f",	--622
		x"02",	--623
		x"b0",	--624
		x"cc",	--625
		x"0d",	--626
		x"0e",	--627
		x"1f",	--628
		x"00",	--629
		x"b0",	--630
		x"48",	--631
		x"0f",	--632
		x"21",	--633
		x"3b",	--634
		x"30",	--635
		x"82",	--636
		x"14",	--637
		x"0a",	--638
		x"82",	--639
		x"14",	--640
		x"1f",	--641
		x"00",	--642
		x"b0",	--643
		x"70",	--644
		x"0f",	--645
		x"21",	--646
		x"3b",	--647
		x"30",	--648
		x"0f",	--649
		x"b0",	--650
		x"82",	--651
		x"0f",	--652
		x"21",	--653
		x"3b",	--654
		x"30",	--655
		x"0e",	--656
		x"3f",	--657
		x"82",	--658
		x"b0",	--659
		x"04",	--660
		x"82",	--661
		x"00",	--662
		x"d3",	--663
		x"82",	--664
		x"16",	--665
		x"30",	--666
		x"0b",	--667
		x"0a",	--668
		x"21",	--669
		x"0a",	--670
		x"0b",	--671
		x"2f",	--672
		x"1b",	--673
		x"0e",	--674
		x"1f",	--675
		x"02",	--676
		x"b0",	--677
		x"cc",	--678
		x"0d",	--679
		x"2a",	--680
		x"18",	--681
		x"0e",	--682
		x"1f",	--683
		x"04",	--684
		x"81",	--685
		x"02",	--686
		x"b0",	--687
		x"cc",	--688
		x"0e",	--689
		x"1d",	--690
		x"02",	--691
		x"1f",	--692
		x"16",	--693
		x"b0",	--694
		x"48",	--695
		x"0f",	--696
		x"21",	--697
		x"3a",	--698
		x"3b",	--699
		x"30",	--700
		x"3d",	--701
		x"64",	--702
		x"3e",	--703
		x"2a",	--704
		x"f2",	--705
		x"3e",	--706
		x"2a",	--707
		x"ef",	--708
		x"1f",	--709
		x"82",	--710
		x"18",	--711
		x"01",	--712
		x"0f",	--713
		x"82",	--714
		x"18",	--715
		x"0f",	--716
		x"30",	--717
		x"5e",	--718
		x"19",	--719
		x"4e",	--720
		x"0f",	--721
		x"03",	--722
		x"c2",	--723
		x"19",	--724
		x"30",	--725
		x"c2",	--726
		x"19",	--727
		x"30",	--728
		x"1e",	--729
		x"1a",	--730
		x"3e",	--731
		x"06",	--732
		x"0f",	--733
		x"0f",	--734
		x"10",	--735
		x"7a",	--736
		x"c2",	--737
		x"19",	--738
		x"3e",	--739
		x"07",	--740
		x"03",	--741
		x"82",	--742
		x"1a",	--743
		x"30",	--744
		x"1e",	--745
		x"82",	--746
		x"1a",	--747
		x"30",	--748
		x"f2",	--749
		x"0e",	--750
		x"19",	--751
		x"f2",	--752
		x"f2",	--753
		x"0a",	--754
		x"19",	--755
		x"ee",	--756
		x"e2",	--757
		x"19",	--758
		x"eb",	--759
		x"f2",	--760
		x"0d",	--761
		x"19",	--762
		x"e7",	--763
		x"f2",	--764
		x"09",	--765
		x"19",	--766
		x"e3",	--767
		x"f2",	--768
		x"03",	--769
		x"19",	--770
		x"df",	--771
		x"f2",	--772
		x"07",	--773
		x"19",	--774
		x"db",	--775
		x"0e",	--776
		x"1f",	--777
		x"1c",	--778
		x"b0",	--779
		x"3a",	--780
		x"0e",	--781
		x"1f",	--782
		x"1e",	--783
		x"b0",	--784
		x"3a",	--785
		x"30",	--786
		x"4c",	--787
		x"b0",	--788
		x"3a",	--789
		x"21",	--790
		x"30",	--791
		x"b2",	--792
		x"02",	--793
		x"09",	--794
		x"1f",	--795
		x"1c",	--796
		x"b0",	--797
		x"f6",	--798
		x"1f",	--799
		x"1e",	--800
		x"b0",	--801
		x"f6",	--802
		x"30",	--803
		x"0e",	--804
		x"3f",	--805
		x"10",	--806
		x"b0",	--807
		x"04",	--808
		x"82",	--809
		x"02",	--810
		x"ef",	--811
		x"82",	--812
		x"1c",	--813
		x"82",	--814
		x"1e",	--815
		x"30",	--816
		x"82",	--817
		x"20",	--818
		x"30",	--819
		x"0b",	--820
		x"0a",	--821
		x"21",	--822
		x"0b",	--823
		x"3f",	--824
		x"03",	--825
		x"30",	--826
		x"23",	--827
		x"0e",	--828
		x"1f",	--829
		x"02",	--830
		x"b0",	--831
		x"9a",	--832
		x"0a",	--833
		x"0e",	--834
		x"1f",	--835
		x"04",	--836
		x"b0",	--837
		x"9a",	--838
		x"0b",	--839
		x"0f",	--840
		x"0a",	--841
		x"30",	--842
		x"83",	--843
		x"b0",	--844
		x"3a",	--845
		x"31",	--846
		x"06",	--847
		x"0e",	--848
		x"1f",	--849
		x"1c",	--850
		x"b0",	--851
		x"3a",	--852
		x"0e",	--853
		x"1f",	--854
		x"1e",	--855
		x"b0",	--856
		x"3a",	--857
		x"0f",	--858
		x"21",	--859
		x"3a",	--860
		x"3b",	--861
		x"30",	--862
		x"0e",	--863
		x"1f",	--864
		x"06",	--865
		x"b0",	--866
		x"cc",	--867
		x"1d",	--868
		x"0e",	--869
		x"1f",	--870
		x"02",	--871
		x"b0",	--872
		x"48",	--873
		x"d1",	--874
		x"30",	--875
		x"53",	--876
		x"b0",	--877
		x"3a",	--878
		x"a1",	--879
		x"00",	--880
		x"30",	--881
		x"64",	--882
		x"b0",	--883
		x"3a",	--884
		x"21",	--885
		x"3f",	--886
		x"e3",	--887
		x"3e",	--888
		x"64",	--889
		x"1f",	--890
		x"1c",	--891
		x"b0",	--892
		x"3a",	--893
		x"3e",	--894
		x"9c",	--895
		x"1f",	--896
		x"1e",	--897
		x"b0",	--898
		x"3a",	--899
		x"1d",	--900
		x"3e",	--901
		x"c8",	--902
		x"1f",	--903
		x"02",	--904
		x"b0",	--905
		x"48",	--906
		x"30",	--907
		x"3e",	--908
		x"9c",	--909
		x"1f",	--910
		x"1c",	--911
		x"b0",	--912
		x"3a",	--913
		x"3e",	--914
		x"64",	--915
		x"1f",	--916
		x"1e",	--917
		x"b0",	--918
		x"3a",	--919
		x"1d",	--920
		x"3e",	--921
		x"c8",	--922
		x"1f",	--923
		x"02",	--924
		x"b0",	--925
		x"48",	--926
		x"30",	--927
		x"3e",	--928
		x"c4",	--929
		x"1f",	--930
		x"1c",	--931
		x"b0",	--932
		x"3a",	--933
		x"3e",	--934
		x"c4",	--935
		x"1f",	--936
		x"1e",	--937
		x"b0",	--938
		x"3a",	--939
		x"1d",	--940
		x"3e",	--941
		x"c8",	--942
		x"1f",	--943
		x"02",	--944
		x"b0",	--945
		x"48",	--946
		x"30",	--947
		x"3e",	--948
		x"3c",	--949
		x"1f",	--950
		x"1c",	--951
		x"b0",	--952
		x"3a",	--953
		x"3e",	--954
		x"3c",	--955
		x"1f",	--956
		x"1e",	--957
		x"b0",	--958
		x"3a",	--959
		x"1d",	--960
		x"3e",	--961
		x"c8",	--962
		x"1f",	--963
		x"02",	--964
		x"b0",	--965
		x"48",	--966
		x"30",	--967
		x"30",	--968
		x"8b",	--969
		x"b0",	--970
		x"3a",	--971
		x"21",	--972
		x"0f",	--973
		x"30",	--974
		x"b2",	--975
		x"00",	--976
		x"92",	--977
		x"b2",	--978
		x"30",	--979
		x"94",	--980
		x"b2",	--981
		x"41",	--982
		x"96",	--983
		x"30",	--984
		x"a1",	--985
		x"b0",	--986
		x"3a",	--987
		x"92",	--988
		x"90",	--989
		x"b1",	--990
		x"bf",	--991
		x"00",	--992
		x"b0",	--993
		x"3a",	--994
		x"21",	--995
		x"0f",	--996
		x"30",	--997
		x"0b",	--998
		x"0a",	--999
		x"8e",	--1000
		x"00",	--1001
		x"6d",	--1002
		x"4d",	--1003
		x"5e",	--1004
		x"1f",	--1005
		x"0a",	--1006
		x"0c",	--1007
		x"0f",	--1008
		x"7b",	--1009
		x"0a",	--1010
		x"2b",	--1011
		x"0c",	--1012
		x"0c",	--1013
		x"0c",	--1014
		x"0c",	--1015
		x"8d",	--1016
		x"0c",	--1017
		x"3c",	--1018
		x"d0",	--1019
		x"1a",	--1020
		x"7d",	--1021
		x"4d",	--1022
		x"17",	--1023
		x"7d",	--1024
		x"78",	--1025
		x"1a",	--1026
		x"4b",	--1027
		x"7b",	--1028
		x"d0",	--1029
		x"0a",	--1030
		x"e9",	--1031
		x"7b",	--1032
		x"0a",	--1033
		x"34",	--1034
		x"0c",	--1035
		x"0b",	--1036
		x"0b",	--1037
		x"0b",	--1038
		x"0c",	--1039
		x"8d",	--1040
		x"0c",	--1041
		x"3c",	--1042
		x"d0",	--1043
		x"7d",	--1044
		x"4d",	--1045
		x"e9",	--1046
		x"9e",	--1047
		x"00",	--1048
		x"0f",	--1049
		x"3a",	--1050
		x"3b",	--1051
		x"30",	--1052
		x"1a",	--1053
		x"de",	--1054
		x"4b",	--1055
		x"7b",	--1056
		x"9f",	--1057
		x"7b",	--1058
		x"06",	--1059
		x"0a",	--1060
		x"0c",	--1061
		x"0c",	--1062
		x"0c",	--1063
		x"0c",	--1064
		x"8d",	--1065
		x"0c",	--1066
		x"3c",	--1067
		x"a9",	--1068
		x"1a",	--1069
		x"ce",	--1070
		x"4b",	--1071
		x"7b",	--1072
		x"bf",	--1073
		x"7b",	--1074
		x"06",	--1075
		x"0a",	--1076
		x"0c",	--1077
		x"0c",	--1078
		x"0c",	--1079
		x"0c",	--1080
		x"8d",	--1081
		x"0c",	--1082
		x"3c",	--1083
		x"c9",	--1084
		x"1a",	--1085
		x"be",	--1086
		x"8d",	--1087
		x"0d",	--1088
		x"30",	--1089
		x"d8",	--1090
		x"b0",	--1091
		x"3a",	--1092
		x"21",	--1093
		x"0c",	--1094
		x"0f",	--1095
		x"3a",	--1096
		x"3b",	--1097
		x"30",	--1098
		x"0c",	--1099
		x"ca",	--1100
		x"0b",	--1101
		x"0a",	--1102
		x"8e",	--1103
		x"00",	--1104
		x"6b",	--1105
		x"4b",	--1106
		x"37",	--1107
		x"1f",	--1108
		x"1a",	--1109
		x"0c",	--1110
		x"12",	--1111
		x"4d",	--1112
		x"7d",	--1113
		x"d0",	--1114
		x"7d",	--1115
		x"0a",	--1116
		x"22",	--1117
		x"0c",	--1118
		x"0d",	--1119
		x"0d",	--1120
		x"0d",	--1121
		x"0c",	--1122
		x"8b",	--1123
		x"0c",	--1124
		x"3c",	--1125
		x"d0",	--1126
		x"7b",	--1127
		x"4b",	--1128
		x"07",	--1129
		x"7b",	--1130
		x"2d",	--1131
		x"eb",	--1132
		x"3a",	--1133
		x"7b",	--1134
		x"4b",	--1135
		x"f9",	--1136
		x"02",	--1137
		x"32",	--1138
		x"03",	--1139
		x"82",	--1140
		x"32",	--1141
		x"82",	--1142
		x"38",	--1143
		x"1f",	--1144
		x"3a",	--1145
		x"32",	--1146
		x"9e",	--1147
		x"00",	--1148
		x"3a",	--1149
		x"3b",	--1150
		x"30",	--1151
		x"8b",	--1152
		x"0b",	--1153
		x"30",	--1154
		x"d8",	--1155
		x"b0",	--1156
		x"3a",	--1157
		x"21",	--1158
		x"0f",	--1159
		x"3a",	--1160
		x"3b",	--1161
		x"30",	--1162
		x"0f",	--1163
		x"ee",	--1164
		x"0b",	--1165
		x"0a",	--1166
		x"09",	--1167
		x"09",	--1168
		x"1f",	--1169
		x"22",	--1170
		x"b0",	--1171
		x"24",	--1172
		x"0a",	--1173
		x"0b",	--1174
		x"1e",	--1175
		x"24",	--1176
		x"1f",	--1177
		x"26",	--1178
		x"b0",	--1179
		x"5c",	--1180
		x"89",	--1181
		x"24",	--1182
		x"89",	--1183
		x"26",	--1184
		x"0d",	--1185
		x"0e",	--1186
		x"0f",	--1187
		x"b0",	--1188
		x"d6",	--1189
		x"0c",	--1190
		x"3d",	--1191
		x"00",	--1192
		x"b0",	--1193
		x"bc",	--1194
		x"0a",	--1195
		x"0b",	--1196
		x"3c",	--1197
		x"66",	--1198
		x"3d",	--1199
		x"66",	--1200
		x"b0",	--1201
		x"1c",	--1202
		x"0f",	--1203
		x"01",	--1204
		x"18",	--1205
		x"3c",	--1206
		x"cd",	--1207
		x"3d",	--1208
		x"cc",	--1209
		x"0e",	--1210
		x"0f",	--1211
		x"b0",	--1212
		x"bc",	--1213
		x"0f",	--1214
		x"04",	--1215
		x"3a",	--1216
		x"cd",	--1217
		x"3b",	--1218
		x"cc",	--1219
		x"0d",	--1220
		x"0e",	--1221
		x"1f",	--1222
		x"20",	--1223
		x"b0",	--1224
		x"1c",	--1225
		x"39",	--1226
		x"3a",	--1227
		x"3b",	--1228
		x"30",	--1229
		x"3a",	--1230
		x"66",	--1231
		x"3b",	--1232
		x"66",	--1233
		x"f1",	--1234
		x"0b",	--1235
		x"0a",	--1236
		x"0b",	--1237
		x"0a",	--1238
		x"8f",	--1239
		x"20",	--1240
		x"8f",	--1241
		x"22",	--1242
		x"11",	--1243
		x"16",	--1244
		x"11",	--1245
		x"16",	--1246
		x"11",	--1247
		x"16",	--1248
		x"11",	--1249
		x"16",	--1250
		x"11",	--1251
		x"16",	--1252
		x"11",	--1253
		x"16",	--1254
		x"1d",	--1255
		x"12",	--1256
		x"1e",	--1257
		x"14",	--1258
		x"b0",	--1259
		x"3c",	--1260
		x"31",	--1261
		x"0c",	--1262
		x"8b",	--1263
		x"28",	--1264
		x"0e",	--1265
		x"3f",	--1266
		x"1a",	--1267
		x"b0",	--1268
		x"04",	--1269
		x"8b",	--1270
		x"2a",	--1271
		x"3a",	--1272
		x"3b",	--1273
		x"30",	--1274
		x"0b",	--1275
		x"0b",	--1276
		x"1f",	--1277
		x"22",	--1278
		x"b0",	--1279
		x"24",	--1280
		x"8b",	--1281
		x"24",	--1282
		x"8b",	--1283
		x"26",	--1284
		x"0d",	--1285
		x"1e",	--1286
		x"28",	--1287
		x"1f",	--1288
		x"2a",	--1289
		x"b0",	--1290
		x"48",	--1291
		x"3b",	--1292
		x"30",	--1293
		x"0b",	--1294
		x"0b",	--1295
		x"0d",	--1296
		x"3e",	--1297
		x"00",	--1298
		x"1f",	--1299
		x"20",	--1300
		x"b0",	--1301
		x"1c",	--1302
		x"1f",	--1303
		x"2a",	--1304
		x"b0",	--1305
		x"70",	--1306
		x"3b",	--1307
		x"30",	--1308
		x"0b",	--1309
		x"0b",	--1310
		x"0d",	--1311
		x"8d",	--1312
		x"8d",	--1313
		x"8d",	--1314
		x"8d",	--1315
		x"0f",	--1316
		x"b0",	--1317
		x"5c",	--1318
		x"0d",	--1319
		x"0e",	--1320
		x"0f",	--1321
		x"b0",	--1322
		x"c2",	--1323
		x"3b",	--1324
		x"30",	--1325
		x"0b",	--1326
		x"0a",	--1327
		x"0a",	--1328
		x"3b",	--1329
		x"00",	--1330
		x"0d",	--1331
		x"0e",	--1332
		x"1f",	--1333
		x"22",	--1334
		x"b0",	--1335
		x"1c",	--1336
		x"0d",	--1337
		x"0e",	--1338
		x"1f",	--1339
		x"24",	--1340
		x"b0",	--1341
		x"1c",	--1342
		x"30",	--1343
		x"ed",	--1344
		x"b0",	--1345
		x"3a",	--1346
		x"21",	--1347
		x"3a",	--1348
		x"3b",	--1349
		x"30",	--1350
		x"82",	--1351
		x"22",	--1352
		x"82",	--1353
		x"24",	--1354
		x"30",	--1355
		x"0b",	--1356
		x"0a",	--1357
		x"21",	--1358
		x"0a",	--1359
		x"0b",	--1360
		x"b2",	--1361
		x"04",	--1362
		x"4e",	--1363
		x"3a",	--1364
		x"03",	--1365
		x"53",	--1366
		x"3e",	--1367
		x"0e",	--1368
		x"1f",	--1369
		x"02",	--1370
		x"b0",	--1371
		x"cc",	--1372
		x"0a",	--1373
		x"0e",	--1374
		x"1f",	--1375
		x"04",	--1376
		x"b0",	--1377
		x"cc",	--1378
		x"0b",	--1379
		x"0f",	--1380
		x"0a",	--1381
		x"30",	--1382
		x"3a",	--1383
		x"b0",	--1384
		x"3a",	--1385
		x"31",	--1386
		x"06",	--1387
		x"0e",	--1388
		x"0f",	--1389
		x"b0",	--1390
		x"92",	--1391
		x"0c",	--1392
		x"3d",	--1393
		x"c8",	--1394
		x"b0",	--1395
		x"7c",	--1396
		x"0c",	--1397
		x"0d",	--1398
		x"0e",	--1399
		x"3f",	--1400
		x"80",	--1401
		x"b0",	--1402
		x"08",	--1403
		x"0d",	--1404
		x"0e",	--1405
		x"1f",	--1406
		x"22",	--1407
		x"b0",	--1408
		x"1c",	--1409
		x"0e",	--1410
		x"0f",	--1411
		x"b0",	--1412
		x"92",	--1413
		x"0c",	--1414
		x"3d",	--1415
		x"c8",	--1416
		x"b0",	--1417
		x"7c",	--1418
		x"0d",	--1419
		x"0e",	--1420
		x"1f",	--1421
		x"24",	--1422
		x"b0",	--1423
		x"1c",	--1424
		x"0f",	--1425
		x"21",	--1426
		x"3a",	--1427
		x"3b",	--1428
		x"30",	--1429
		x"0e",	--1430
		x"1f",	--1431
		x"06",	--1432
		x"b0",	--1433
		x"cc",	--1434
		x"1d",	--1435
		x"0e",	--1436
		x"1f",	--1437
		x"04",	--1438
		x"b0",	--1439
		x"48",	--1440
		x"b6",	--1441
		x"0e",	--1442
		x"3f",	--1443
		x"5c",	--1444
		x"b0",	--1445
		x"04",	--1446
		x"82",	--1447
		x"04",	--1448
		x"aa",	--1449
		x"30",	--1450
		x"f4",	--1451
		x"b0",	--1452
		x"3a",	--1453
		x"b1",	--1454
		x"0e",	--1455
		x"00",	--1456
		x"b0",	--1457
		x"3a",	--1458
		x"a1",	--1459
		x"00",	--1460
		x"30",	--1461
		x"1f",	--1462
		x"b0",	--1463
		x"3a",	--1464
		x"21",	--1465
		x"3f",	--1466
		x"d6",	--1467
		x"0b",	--1468
		x"0a",	--1469
		x"1f",	--1470
		x"28",	--1471
		x"b0",	--1472
		x"24",	--1473
		x"0a",	--1474
		x"0b",	--1475
		x"1f",	--1476
		x"26",	--1477
		x"b0",	--1478
		x"24",	--1479
		x"0b",	--1480
		x"0a",	--1481
		x"3e",	--1482
		x"3f",	--1483
		x"1e",	--1484
		x"0f",	--1485
		x"0f",	--1486
		x"0e",	--1487
		x"30",	--1488
		x"42",	--1489
		x"30",	--1490
		x"4c",	--1491
		x"b0",	--1492
		x"ea",	--1493
		x"31",	--1494
		x"0c",	--1495
		x"30",	--1496
		x"4c",	--1497
		x"30",	--1498
		x"4a",	--1499
		x"b0",	--1500
		x"3a",	--1501
		x"21",	--1502
		x"3a",	--1503
		x"3b",	--1504
		x"30",	--1505
		x"82",	--1506
		x"26",	--1507
		x"82",	--1508
		x"28",	--1509
		x"30",	--1510
		x"82",	--1511
		x"2a",	--1512
		x"82",	--1513
		x"2c",	--1514
		x"30",	--1515
		x"0b",	--1516
		x"0a",	--1517
		x"09",	--1518
		x"08",	--1519
		x"21",	--1520
		x"0a",	--1521
		x"0b",	--1522
		x"81",	--1523
		x"00",	--1524
		x"1f",	--1525
		x"1c",	--1526
		x"b2",	--1527
		x"06",	--1528
		x"6f",	--1529
		x"92",	--1530
		x"2e",	--1531
		x"0e",	--1532
		x"1f",	--1533
		x"02",	--1534
		x"b0",	--1535
		x"cc",	--1536
		x"08",	--1537
		x"3a",	--1538
		x"03",	--1539
		x"1e",	--1540
		x"09",	--1541
		x"0d",	--1542
		x"0e",	--1543
		x"1f",	--1544
		x"06",	--1545
		x"b0",	--1546
		x"48",	--1547
		x"0f",	--1548
		x"21",	--1549
		x"38",	--1550
		x"39",	--1551
		x"3a",	--1552
		x"3b",	--1553
		x"30",	--1554
		x"82",	--1555
		x"2e",	--1556
		x"49",	--1557
		x"82",	--1558
		x"2e",	--1559
		x"1f",	--1560
		x"06",	--1561
		x"b0",	--1562
		x"70",	--1563
		x"0f",	--1564
		x"21",	--1565
		x"38",	--1566
		x"39",	--1567
		x"3a",	--1568
		x"3b",	--1569
		x"30",	--1570
		x"0e",	--1571
		x"1f",	--1572
		x"04",	--1573
		x"b0",	--1574
		x"cc",	--1575
		x"09",	--1576
		x"3a",	--1577
		x"05",	--1578
		x"da",	--1579
		x"0e",	--1580
		x"1f",	--1581
		x"06",	--1582
		x"b0",	--1583
		x"cc",	--1584
		x"0a",	--1585
		x"0e",	--1586
		x"1f",	--1587
		x"08",	--1588
		x"b0",	--1589
		x"cc",	--1590
		x"0b",	--1591
		x"0f",	--1592
		x"0a",	--1593
		x"30",	--1594
		x"4f",	--1595
		x"b0",	--1596
		x"3a",	--1597
		x"31",	--1598
		x"06",	--1599
		x"0e",	--1600
		x"0f",	--1601
		x"b0",	--1602
		x"92",	--1603
		x"0c",	--1604
		x"3d",	--1605
		x"c8",	--1606
		x"b0",	--1607
		x"7c",	--1608
		x"0d",	--1609
		x"0e",	--1610
		x"1f",	--1611
		x"2a",	--1612
		x"b0",	--1613
		x"1c",	--1614
		x"0e",	--1615
		x"0f",	--1616
		x"b0",	--1617
		x"92",	--1618
		x"0c",	--1619
		x"3d",	--1620
		x"c8",	--1621
		x"b0",	--1622
		x"7c",	--1623
		x"0d",	--1624
		x"0e",	--1625
		x"1f",	--1626
		x"2c",	--1627
		x"b0",	--1628
		x"1c",	--1629
		x"a7",	--1630
		x"0f",	--1631
		x"b0",	--1632
		x"78",	--1633
		x"0f",	--1634
		x"21",	--1635
		x"38",	--1636
		x"39",	--1637
		x"3a",	--1638
		x"3b",	--1639
		x"30",	--1640
		x"0e",	--1641
		x"3f",	--1642
		x"78",	--1643
		x"b0",	--1644
		x"04",	--1645
		x"82",	--1646
		x"06",	--1647
		x"89",	--1648
		x"0b",	--1649
		x"0a",	--1650
		x"09",	--1651
		x"08",	--1652
		x"08",	--1653
		x"3a",	--1654
		x"08",	--1655
		x"09",	--1656
		x"0b",	--1657
		x"0e",	--1658
		x"0f",	--1659
		x"b0",	--1660
		x"be",	--1661
		x"2f",	--1662
		x"09",	--1663
		x"1e",	--1664
		x"4d",	--1665
		x"7d",	--1666
		x"0f",	--1667
		x"03",	--1668
		x"0e",	--1669
		x"7d",	--1670
		x"fd",	--1671
		x"09",	--1672
		x"1b",	--1673
		x"2a",	--1674
		x"3b",	--1675
		x"05",	--1676
		x"ec",	--1677
		x"0f",	--1678
		x"38",	--1679
		x"39",	--1680
		x"3a",	--1681
		x"3b",	--1682
		x"30",	--1683
		x"0b",	--1684
		x"0a",	--1685
		x"82",	--1686
		x"30",	--1687
		x"03",	--1688
		x"3a",	--1689
		x"3b",	--1690
		x"30",	--1691
		x"1f",	--1692
		x"32",	--1693
		x"b0",	--1694
		x"e2",	--1695
		x"0a",	--1696
		x"0b",	--1697
		x"0e",	--1698
		x"1f",	--1699
		x"32",	--1700
		x"b0",	--1701
		x"be",	--1702
		x"0f",	--1703
		x"30",	--1704
		x"58",	--1705
		x"b0",	--1706
		x"3a",	--1707
		x"21",	--1708
		x"1b",	--1709
		x"3b",	--1710
		x"05",	--1711
		x"f1",	--1712
		x"30",	--1713
		x"5c",	--1714
		x"b0",	--1715
		x"3a",	--1716
		x"21",	--1717
		x"1f",	--1718
		x"34",	--1719
		x"0f",	--1720
		x"22",	--1721
		x"0a",	--1722
		x"74",	--1723
		x"3a",	--1724
		x"7f",	--1725
		x"2a",	--1726
		x"83",	--1727
		x"1a",	--1728
		x"99",	--1729
		x"2a",	--1730
		x"47",	--1731
		x"a2",	--1732
		x"34",	--1733
		x"0e",	--1734
		x"1f",	--1735
		x"36",	--1736
		x"b0",	--1737
		x"3a",	--1738
		x"0e",	--1739
		x"1f",	--1740
		x"38",	--1741
		x"b0",	--1742
		x"3a",	--1743
		x"b2",	--1744
		x"14",	--1745
		x"3a",	--1746
		x"b2",	--1747
		x"0a",	--1748
		x"3c",	--1749
		x"30",	--1750
		x"8e",	--1751
		x"b0",	--1752
		x"3a",	--1753
		x"21",	--1754
		x"bd",	--1755
		x"82",	--1756
		x"3a",	--1757
		x"12",	--1758
		x"1e",	--1759
		x"3c",	--1760
		x"0e",	--1761
		x"0b",	--1762
		x"1f",	--1763
		x"8f",	--1764
		x"2f",	--1765
		x"ae",	--1766
		x"3f",	--1767
		x"03",	--1768
		x"32",	--1769
		x"3e",	--1770
		x"82",	--1771
		x"3c",	--1772
		x"ab",	--1773
		x"82",	--1774
		x"34",	--1775
		x"a8",	--1776
		x"0e",	--1777
		x"1f",	--1778
		x"36",	--1779
		x"b0",	--1780
		x"3a",	--1781
		x"0e",	--1782
		x"1f",	--1783
		x"38",	--1784
		x"b0",	--1785
		x"3a",	--1786
		x"30",	--1787
		x"a4",	--1788
		x"b0",	--1789
		x"3a",	--1790
		x"21",	--1791
		x"b2",	--1792
		x"3a",	--1793
		x"0a",	--1794
		x"95",	--1795
		x"82",	--1796
		x"3a",	--1797
		x"82",	--1798
		x"3c",	--1799
		x"82",	--1800
		x"34",	--1801
		x"8e",	--1802
		x"0e",	--1803
		x"1f",	--1804
		x"36",	--1805
		x"b0",	--1806
		x"3a",	--1807
		x"0e",	--1808
		x"1f",	--1809
		x"38",	--1810
		x"b0",	--1811
		x"3a",	--1812
		x"0a",	--1813
		x"30",	--1814
		x"9f",	--1815
		x"b0",	--1816
		x"3a",	--1817
		x"21",	--1818
		x"7d",	--1819
		x"3e",	--1820
		x"1e",	--1821
		x"1f",	--1822
		x"36",	--1823
		x"b0",	--1824
		x"3a",	--1825
		x"3e",	--1826
		x"1e",	--1827
		x"1f",	--1828
		x"38",	--1829
		x"b0",	--1830
		x"3a",	--1831
		x"30",	--1832
		x"cc",	--1833
		x"b0",	--1834
		x"3a",	--1835
		x"21",	--1836
		x"1e",	--1837
		x"3c",	--1838
		x"ba",	--1839
		x"3e",	--1840
		x"3c",	--1841
		x"1f",	--1842
		x"36",	--1843
		x"b0",	--1844
		x"3a",	--1845
		x"3e",	--1846
		x"c4",	--1847
		x"1f",	--1848
		x"38",	--1849
		x"b0",	--1850
		x"3a",	--1851
		x"5c",	--1852
		x"30",	--1853
		x"5f",	--1854
		x"b0",	--1855
		x"3a",	--1856
		x"21",	--1857
		x"56",	--1858
		x"92",	--1859
		x"34",	--1860
		x"0e",	--1861
		x"1f",	--1862
		x"36",	--1863
		x"b0",	--1864
		x"3a",	--1865
		x"0e",	--1866
		x"1f",	--1867
		x"38",	--1868
		x"b0",	--1869
		x"3a",	--1870
		x"b2",	--1871
		x"14",	--1872
		x"3a",	--1873
		x"b2",	--1874
		x"14",	--1875
		x"3c",	--1876
		x"30",	--1877
		x"6e",	--1878
		x"b0",	--1879
		x"3a",	--1880
		x"21",	--1881
		x"3e",	--1882
		x"b2",	--1883
		x"03",	--1884
		x"34",	--1885
		x"0e",	--1886
		x"1f",	--1887
		x"36",	--1888
		x"b0",	--1889
		x"3a",	--1890
		x"0e",	--1891
		x"1f",	--1892
		x"38",	--1893
		x"b0",	--1894
		x"3a",	--1895
		x"b2",	--1896
		x"14",	--1897
		x"3a",	--1898
		x"b2",	--1899
		x"0a",	--1900
		x"3c",	--1901
		x"30",	--1902
		x"7c",	--1903
		x"b0",	--1904
		x"3a",	--1905
		x"21",	--1906
		x"25",	--1907
		x"0e",	--1908
		x"1f",	--1909
		x"32",	--1910
		x"b0",	--1911
		x"be",	--1912
		x"0b",	--1913
		x"2e",	--1914
		x"1f",	--1915
		x"32",	--1916
		x"b0",	--1917
		x"be",	--1918
		x"0b",	--1919
		x"28",	--1920
		x"3e",	--1921
		x"1e",	--1922
		x"1f",	--1923
		x"36",	--1924
		x"b0",	--1925
		x"3a",	--1926
		x"3e",	--1927
		x"1e",	--1928
		x"1f",	--1929
		x"38",	--1930
		x"b0",	--1931
		x"3a",	--1932
		x"30",	--1933
		x"ab",	--1934
		x"b0",	--1935
		x"3a",	--1936
		x"21",	--1937
		x"1e",	--1938
		x"3c",	--1939
		x"55",	--1940
		x"3e",	--1941
		x"e2",	--1942
		x"1f",	--1943
		x"36",	--1944
		x"b0",	--1945
		x"3a",	--1946
		x"3e",	--1947
		x"e2",	--1948
		x"1f",	--1949
		x"38",	--1950
		x"b0",	--1951
		x"3a",	--1952
		x"30",	--1953
		x"bc",	--1954
		x"b0",	--1955
		x"3a",	--1956
		x"21",	--1957
		x"1e",	--1958
		x"3c",	--1959
		x"41",	--1960
		x"3e",	--1961
		x"e2",	--1962
		x"1f",	--1963
		x"36",	--1964
		x"b0",	--1965
		x"3a",	--1966
		x"3e",	--1967
		x"e2",	--1968
		x"1f",	--1969
		x"38",	--1970
		x"b0",	--1971
		x"3a",	--1972
		x"d7",	--1973
		x"82",	--1974
		x"36",	--1975
		x"82",	--1976
		x"38",	--1977
		x"30",	--1978
		x"82",	--1979
		x"32",	--1980
		x"30",	--1981
		x"0b",	--1982
		x"0b",	--1983
		x"0e",	--1984
		x"3f",	--1985
		x"28",	--1986
		x"b0",	--1987
		x"04",	--1988
		x"82",	--1989
		x"3e",	--1990
		x"0d",	--1991
		x"0e",	--1992
		x"b0",	--1993
		x"48",	--1994
		x"3b",	--1995
		x"30",	--1996
		x"0b",	--1997
		x"0b",	--1998
		x"1f",	--1999
		x"0e",	--2000
		x"2f",	--2001
		x"09",	--2002
		x"1f",	--2003
		x"02",	--2004
		x"6f",	--2005
		x"7f",	--2006
		x"30",	--2007
		x"30",	--2008
		x"7f",	--2009
		x"31",	--2010
		x"2a",	--2011
		x"0f",	--2012
		x"3b",	--2013
		x"30",	--2014
		x"82",	--2015
		x"30",	--2016
		x"1e",	--2017
		x"82",	--2018
		x"30",	--2019
		x"0f",	--2020
		x"08",	--2021
		x"30",	--2022
		x"dd",	--2023
		x"b0",	--2024
		x"3a",	--2025
		x"21",	--2026
		x"0f",	--2027
		x"3b",	--2028
		x"30",	--2029
		x"0e",	--2030
		x"1f",	--2031
		x"36",	--2032
		x"b0",	--2033
		x"3a",	--2034
		x"0e",	--2035
		x"1f",	--2036
		x"38",	--2037
		x"b0",	--2038
		x"3a",	--2039
		x"30",	--2040
		x"f1",	--2041
		x"b0",	--2042
		x"3a",	--2043
		x"21",	--2044
		x"0f",	--2045
		x"3b",	--2046
		x"30",	--2047
		x"0f",	--2048
		x"82",	--2049
		x"30",	--2050
		x"0f",	--2051
		x"e9",	--2052
		x"e0",	--2053
		x"92",	--2054
		x"30",	--2055
		x"dd",	--2056
		x"82",	--2057
		x"30",	--2058
		x"30",	--2059
		x"f1",	--2060
		x"b0",	--2061
		x"3a",	--2062
		x"21",	--2063
		x"0e",	--2064
		x"1f",	--2065
		x"36",	--2066
		x"b0",	--2067
		x"3a",	--2068
		x"0e",	--2069
		x"1f",	--2070
		x"38",	--2071
		x"b0",	--2072
		x"3a",	--2073
		x"1f",	--2074
		x"02",	--2075
		x"6f",	--2076
		x"bb",	--2077
		x"8f",	--2078
		x"00",	--2079
		x"8f",	--2080
		x"02",	--2081
		x"9f",	--2082
		x"02",	--2083
		x"04",	--2084
		x"9f",	--2085
		x"04",	--2086
		x"06",	--2087
		x"9f",	--2088
		x"06",	--2089
		x"08",	--2090
		x"9f",	--2091
		x"08",	--2092
		x"0a",	--2093
		x"9f",	--2094
		x"0a",	--2095
		x"10",	--2096
		x"9f",	--2097
		x"0c",	--2098
		x"12",	--2099
		x"8f",	--2100
		x"14",	--2101
		x"8f",	--2102
		x"16",	--2103
		x"8f",	--2104
		x"0c",	--2105
		x"8f",	--2106
		x"0e",	--2107
		x"8f",	--2108
		x"18",	--2109
		x"8f",	--2110
		x"1a",	--2111
		x"8f",	--2112
		x"1c",	--2113
		x"8f",	--2114
		x"1e",	--2115
		x"30",	--2116
		x"8f",	--2117
		x"0c",	--2118
		x"8f",	--2119
		x"0e",	--2120
		x"8f",	--2121
		x"18",	--2122
		x"8f",	--2123
		x"1a",	--2124
		x"8f",	--2125
		x"1c",	--2126
		x"8f",	--2127
		x"1e",	--2128
		x"30",	--2129
		x"8f",	--2130
		x"00",	--2131
		x"8f",	--2132
		x"02",	--2133
		x"30",	--2134
		x"8f",	--2135
		x"04",	--2136
		x"8f",	--2137
		x"06",	--2138
		x"30",	--2139
		x"8f",	--2140
		x"08",	--2141
		x"8f",	--2142
		x"0a",	--2143
		x"30",	--2144
		x"8f",	--2145
		x"0c",	--2146
		x"8f",	--2147
		x"0e",	--2148
		x"30",	--2149
		x"8f",	--2150
		x"10",	--2151
		x"8f",	--2152
		x"12",	--2153
		x"30",	--2154
		x"0b",	--2155
		x"0a",	--2156
		x"09",	--2157
		x"07",	--2158
		x"06",	--2159
		x"05",	--2160
		x"04",	--2161
		x"09",	--2162
		x"04",	--2163
		x"05",	--2164
		x"16",	--2165
		x"14",	--2166
		x"17",	--2167
		x"16",	--2168
		x"1a",	--2169
		x"0c",	--2170
		x"1b",	--2171
		x"0e",	--2172
		x"0c",	--2173
		x"0d",	--2174
		x"0e",	--2175
		x"0f",	--2176
		x"b0",	--2177
		x"bc",	--2178
		x"1c",	--2179
		x"10",	--2180
		x"1d",	--2181
		x"12",	--2182
		x"0f",	--2183
		x"5b",	--2184
		x"0e",	--2185
		x"0f",	--2186
		x"b0",	--2187
		x"bc",	--2188
		x"06",	--2189
		x"07",	--2190
		x"89",	--2191
		x"14",	--2192
		x"89",	--2193
		x"16",	--2194
		x"0c",	--2195
		x"0d",	--2196
		x"0e",	--2197
		x"0f",	--2198
		x"b0",	--2199
		x"bc",	--2200
		x"0f",	--2201
		x"5c",	--2202
		x"89",	--2203
		x"14",	--2204
		x"89",	--2205
		x"16",	--2206
		x"0c",	--2207
		x"0d",	--2208
		x"0e",	--2209
		x"0f",	--2210
		x"b0",	--2211
		x"08",	--2212
		x"0a",	--2213
		x"0b",	--2214
		x"1c",	--2215
		x"18",	--2216
		x"1d",	--2217
		x"1a",	--2218
		x"b0",	--2219
		x"bc",	--2220
		x"06",	--2221
		x"07",	--2222
		x"89",	--2223
		x"18",	--2224
		x"89",	--2225
		x"1a",	--2226
		x"2c",	--2227
		x"1d",	--2228
		x"02",	--2229
		x"0e",	--2230
		x"0f",	--2231
		x"b0",	--2232
		x"58",	--2233
		x"04",	--2234
		x"05",	--2235
		x"1c",	--2236
		x"04",	--2237
		x"1d",	--2238
		x"06",	--2239
		x"0e",	--2240
		x"0f",	--2241
		x"b0",	--2242
		x"58",	--2243
		x"0c",	--2244
		x"0d",	--2245
		x"b0",	--2246
		x"bc",	--2247
		x"06",	--2248
		x"07",	--2249
		x"1c",	--2250
		x"1c",	--2251
		x"1d",	--2252
		x"1e",	--2253
		x"0e",	--2254
		x"0f",	--2255
		x"b0",	--2256
		x"08",	--2257
		x"1c",	--2258
		x"08",	--2259
		x"1d",	--2260
		x"0a",	--2261
		x"b0",	--2262
		x"58",	--2263
		x"0c",	--2264
		x"0d",	--2265
		x"b0",	--2266
		x"bc",	--2267
		x"34",	--2268
		x"35",	--2269
		x"36",	--2270
		x"37",	--2271
		x"39",	--2272
		x"3a",	--2273
		x"3b",	--2274
		x"30",	--2275
		x"0e",	--2276
		x"0f",	--2277
		x"b0",	--2278
		x"08",	--2279
		x"06",	--2280
		x"07",	--2281
		x"89",	--2282
		x"14",	--2283
		x"89",	--2284
		x"16",	--2285
		x"0c",	--2286
		x"0d",	--2287
		x"0e",	--2288
		x"0f",	--2289
		x"b0",	--2290
		x"1c",	--2291
		x"0f",	--2292
		x"01",	--2293
		x"a4",	--2294
		x"0a",	--2295
		x"0b",	--2296
		x"a5",	--2297
		x"0b",	--2298
		x"0a",	--2299
		x"21",	--2300
		x"0a",	--2301
		x"0b",	--2302
		x"30",	--2303
		x"12",	--2304
		x"b0",	--2305
		x"3a",	--2306
		x"21",	--2307
		x"3a",	--2308
		x"03",	--2309
		x"1b",	--2310
		x"0e",	--2311
		x"1f",	--2312
		x"02",	--2313
		x"b0",	--2314
		x"cc",	--2315
		x"0a",	--2316
		x"0e",	--2317
		x"1f",	--2318
		x"04",	--2319
		x"b0",	--2320
		x"cc",	--2321
		x"0b",	--2322
		x"0f",	--2323
		x"0a",	--2324
		x"30",	--2325
		x"5a",	--2326
		x"b0",	--2327
		x"3a",	--2328
		x"31",	--2329
		x"06",	--2330
		x"8a",	--2331
		x"00",	--2332
		x"0f",	--2333
		x"21",	--2334
		x"3a",	--2335
		x"3b",	--2336
		x"30",	--2337
		x"30",	--2338
		x"1a",	--2339
		x"b0",	--2340
		x"3a",	--2341
		x"b1",	--2342
		x"34",	--2343
		x"00",	--2344
		x"b0",	--2345
		x"3a",	--2346
		x"a1",	--2347
		x"00",	--2348
		x"30",	--2349
		x"45",	--2350
		x"b0",	--2351
		x"3a",	--2352
		x"21",	--2353
		x"3f",	--2354
		x"ea",	--2355
		x"0b",	--2356
		x"21",	--2357
		x"0b",	--2358
		x"1f",	--2359
		x"17",	--2360
		x"16",	--2361
		x"30",	--2362
		x"75",	--2363
		x"b0",	--2364
		x"3a",	--2365
		x"21",	--2366
		x"0e",	--2367
		x"1f",	--2368
		x"02",	--2369
		x"b0",	--2370
		x"cc",	--2371
		x"2f",	--2372
		x"0f",	--2373
		x"30",	--2374
		x"5a",	--2375
		x"b0",	--2376
		x"3a",	--2377
		x"31",	--2378
		x"06",	--2379
		x"0f",	--2380
		x"21",	--2381
		x"3b",	--2382
		x"30",	--2383
		x"30",	--2384
		x"1a",	--2385
		x"b0",	--2386
		x"3a",	--2387
		x"b1",	--2388
		x"34",	--2389
		x"00",	--2390
		x"b0",	--2391
		x"3a",	--2392
		x"a1",	--2393
		x"00",	--2394
		x"30",	--2395
		x"66",	--2396
		x"b0",	--2397
		x"3a",	--2398
		x"21",	--2399
		x"3f",	--2400
		x"eb",	--2401
		x"0b",	--2402
		x"0a",	--2403
		x"09",	--2404
		x"08",	--2405
		x"07",	--2406
		x"06",	--2407
		x"06",	--2408
		x"07",	--2409
		x"08",	--2410
		x"09",	--2411
		x"b0",	--2412
		x"bc",	--2413
		x"0a",	--2414
		x"0b",	--2415
		x"3c",	--2416
		x"db",	--2417
		x"3d",	--2418
		x"49",	--2419
		x"b0",	--2420
		x"0c",	--2421
		x"0f",	--2422
		x"20",	--2423
		x"1f",	--2424
		x"3c",	--2425
		x"db",	--2426
		x"3d",	--2427
		x"49",	--2428
		x"0e",	--2429
		x"0f",	--2430
		x"b0",	--2431
		x"1c",	--2432
		x"0f",	--2433
		x"01",	--2434
		x"09",	--2435
		x"0e",	--2436
		x"0f",	--2437
		x"36",	--2438
		x"37",	--2439
		x"38",	--2440
		x"39",	--2441
		x"3a",	--2442
		x"3b",	--2443
		x"30",	--2444
		x"3c",	--2445
		x"db",	--2446
		x"3d",	--2447
		x"c9",	--2448
		x"0e",	--2449
		x"0f",	--2450
		x"b0",	--2451
		x"08",	--2452
		x"0a",	--2453
		x"0b",	--2454
		x"ec",	--2455
		x"3c",	--2456
		x"db",	--2457
		x"3d",	--2458
		x"c9",	--2459
		x"0e",	--2460
		x"0f",	--2461
		x"b0",	--2462
		x"bc",	--2463
		x"0c",	--2464
		x"0d",	--2465
		x"b0",	--2466
		x"bc",	--2467
		x"0a",	--2468
		x"0b",	--2469
		x"dd",	--2470
		x"0b",	--2471
		x"0b",	--2472
		x"8f",	--2473
		x"0a",	--2474
		x"8f",	--2475
		x"0c",	--2476
		x"8f",	--2477
		x"0e",	--2478
		x"8f",	--2479
		x"10",	--2480
		x"8f",	--2481
		x"12",	--2482
		x"8f",	--2483
		x"14",	--2484
		x"8f",	--2485
		x"00",	--2486
		x"8f",	--2487
		x"02",	--2488
		x"9f",	--2489
		x"04",	--2490
		x"04",	--2491
		x"9f",	--2492
		x"06",	--2493
		x"06",	--2494
		x"9f",	--2495
		x"08",	--2496
		x"08",	--2497
		x"8f",	--2498
		x"16",	--2499
		x"8f",	--2500
		x"18",	--2501
		x"8f",	--2502
		x"1a",	--2503
		x"8f",	--2504
		x"1c",	--2505
		x"0e",	--2506
		x"3f",	--2507
		x"2a",	--2508
		x"b0",	--2509
		x"04",	--2510
		x"8b",	--2511
		x"22",	--2512
		x"3b",	--2513
		x"30",	--2514
		x"8f",	--2515
		x"20",	--2516
		x"8f",	--2517
		x"1e",	--2518
		x"30",	--2519
		x"0b",	--2520
		x"0a",	--2521
		x"09",	--2522
		x"08",	--2523
		x"07",	--2524
		x"05",	--2525
		x"04",	--2526
		x"31",	--2527
		x"f4",	--2528
		x"07",	--2529
		x"81",	--2530
		x"04",	--2531
		x"81",	--2532
		x"06",	--2533
		x"3c",	--2534
		x"db",	--2535
		x"3d",	--2536
		x"c9",	--2537
		x"2e",	--2538
		x"1f",	--2539
		x"02",	--2540
		x"b0",	--2541
		x"58",	--2542
		x"0a",	--2543
		x"0b",	--2544
		x"1e",	--2545
		x"08",	--2546
		x"0f",	--2547
		x"8f",	--2548
		x"8f",	--2549
		x"8f",	--2550
		x"8f",	--2551
		x"b0",	--2552
		x"5c",	--2553
		x"0c",	--2554
		x"0d",	--2555
		x"0e",	--2556
		x"0f",	--2557
		x"b0",	--2558
		x"7c",	--2559
		x"0a",	--2560
		x"0b",	--2561
		x"18",	--2562
		x"04",	--2563
		x"19",	--2564
		x"06",	--2565
		x"18",	--2566
		x"16",	--2567
		x"19",	--2568
		x"18",	--2569
		x"14",	--2570
		x"1c",	--2571
		x"15",	--2572
		x"1e",	--2573
		x"14",	--2574
		x"1a",	--2575
		x"15",	--2576
		x"1c",	--2577
		x"0e",	--2578
		x"0f",	--2579
		x"b0",	--2580
		x"5c",	--2581
		x"0c",	--2582
		x"0d",	--2583
		x"b0",	--2584
		x"58",	--2585
		x"81",	--2586
		x"00",	--2587
		x"81",	--2588
		x"02",	--2589
		x"0e",	--2590
		x"0f",	--2591
		x"b0",	--2592
		x"5c",	--2593
		x"0c",	--2594
		x"0d",	--2595
		x"b0",	--2596
		x"58",	--2597
		x"0a",	--2598
		x"0b",	--2599
		x"0c",	--2600
		x"0d",	--2601
		x"2e",	--2602
		x"1f",	--2603
		x"02",	--2604
		x"b0",	--2605
		x"bc",	--2606
		x"81",	--2607
		x"08",	--2608
		x"81",	--2609
		x"0a",	--2610
		x"08",	--2611
		x"a0",	--2612
		x"09",	--2613
		x"9e",	--2614
		x"04",	--2615
		x"02",	--2616
		x"30",	--2617
		x"22",	--2618
		x"18",	--2619
		x"04",	--2620
		x"19",	--2621
		x"06",	--2622
		x"2c",	--2623
		x"1d",	--2624
		x"02",	--2625
		x"0e",	--2626
		x"0f",	--2627
		x"b0",	--2628
		x"08",	--2629
		x"0a",	--2630
		x"0b",	--2631
		x"0c",	--2632
		x"0d",	--2633
		x"1e",	--2634
		x"08",	--2635
		x"1f",	--2636
		x"0a",	--2637
		x"b0",	--2638
		x"58",	--2639
		x"0c",	--2640
		x"0d",	--2641
		x"b0",	--2642
		x"7c",	--2643
		x"04",	--2644
		x"05",	--2645
		x"0c",	--2646
		x"0d",	--2647
		x"0e",	--2648
		x"0f",	--2649
		x"b0",	--2650
		x"bc",	--2651
		x"0c",	--2652
		x"0d",	--2653
		x"0e",	--2654
		x"0f",	--2655
		x"b0",	--2656
		x"7c",	--2657
		x"b0",	--2658
		x"3e",	--2659
		x"81",	--2660
		x"00",	--2661
		x"81",	--2662
		x"02",	--2663
		x"1a",	--2664
		x"12",	--2665
		x"1b",	--2666
		x"14",	--2667
		x"0e",	--2668
		x"0f",	--2669
		x"b0",	--2670
		x"e4",	--2671
		x"0c",	--2672
		x"0d",	--2673
		x"b0",	--2674
		x"58",	--2675
		x"0c",	--2676
		x"0d",	--2677
		x"1e",	--2678
		x"0a",	--2679
		x"1f",	--2680
		x"0c",	--2681
		x"b0",	--2682
		x"08",	--2683
		x"81",	--2684
		x"08",	--2685
		x"81",	--2686
		x"0a",	--2687
		x"0e",	--2688
		x"0f",	--2689
		x"b0",	--2690
		x"be",	--2691
		x"0c",	--2692
		x"0d",	--2693
		x"b0",	--2694
		x"58",	--2695
		x"1c",	--2696
		x"0e",	--2697
		x"1d",	--2698
		x"10",	--2699
		x"b0",	--2700
		x"bc",	--2701
		x"08",	--2702
		x"09",	--2703
		x"2c",	--2704
		x"1d",	--2705
		x"02",	--2706
		x"0e",	--2707
		x"0f",	--2708
		x"b0",	--2709
		x"c4",	--2710
		x"0a",	--2711
		x"0b",	--2712
		x"87",	--2713
		x"12",	--2714
		x"87",	--2715
		x"14",	--2716
		x"b0",	--2717
		x"e4",	--2718
		x"0c",	--2719
		x"0d",	--2720
		x"b0",	--2721
		x"58",	--2722
		x"1c",	--2723
		x"08",	--2724
		x"1d",	--2725
		x"0a",	--2726
		x"b0",	--2727
		x"bc",	--2728
		x"87",	--2729
		x"0a",	--2730
		x"87",	--2731
		x"0c",	--2732
		x"0e",	--2733
		x"0f",	--2734
		x"b0",	--2735
		x"be",	--2736
		x"0c",	--2737
		x"0d",	--2738
		x"b0",	--2739
		x"58",	--2740
		x"0c",	--2741
		x"0d",	--2742
		x"0e",	--2743
		x"0f",	--2744
		x"b0",	--2745
		x"08",	--2746
		x"87",	--2747
		x"0e",	--2748
		x"87",	--2749
		x"10",	--2750
		x"97",	--2751
		x"04",	--2752
		x"16",	--2753
		x"97",	--2754
		x"06",	--2755
		x"18",	--2756
		x"97",	--2757
		x"1c",	--2758
		x"1a",	--2759
		x"97",	--2760
		x"1e",	--2761
		x"1c",	--2762
		x"31",	--2763
		x"0c",	--2764
		x"34",	--2765
		x"35",	--2766
		x"37",	--2767
		x"38",	--2768
		x"39",	--2769
		x"3a",	--2770
		x"3b",	--2771
		x"30",	--2772
		x"08",	--2773
		x"64",	--2774
		x"09",	--2775
		x"62",	--2776
		x"0c",	--2777
		x"3d",	--2778
		x"00",	--2779
		x"1e",	--2780
		x"08",	--2781
		x"1f",	--2782
		x"0a",	--2783
		x"b0",	--2784
		x"58",	--2785
		x"0a",	--2786
		x"0b",	--2787
		x"18",	--2788
		x"12",	--2789
		x"19",	--2790
		x"14",	--2791
		x"0e",	--2792
		x"0f",	--2793
		x"b0",	--2794
		x"be",	--2795
		x"0c",	--2796
		x"0d",	--2797
		x"b0",	--2798
		x"58",	--2799
		x"0c",	--2800
		x"0d",	--2801
		x"1e",	--2802
		x"0a",	--2803
		x"1f",	--2804
		x"0c",	--2805
		x"b0",	--2806
		x"bc",	--2807
		x"87",	--2808
		x"0a",	--2809
		x"87",	--2810
		x"0c",	--2811
		x"0e",	--2812
		x"0f",	--2813
		x"b0",	--2814
		x"e4",	--2815
		x"0c",	--2816
		x"0d",	--2817
		x"b0",	--2818
		x"58",	--2819
		x"0c",	--2820
		x"0d",	--2821
		x"1e",	--2822
		x"0e",	--2823
		x"1f",	--2824
		x"10",	--2825
		x"b0",	--2826
		x"bc",	--2827
		x"87",	--2828
		x"0e",	--2829
		x"87",	--2830
		x"10",	--2831
		x"ae",	--2832
		x"05",	--2833
		x"ac",	--2834
		x"30",	--2835
		x"76",	--2836
		x"0b",	--2837
		x"0a",	--2838
		x"09",	--2839
		x"09",	--2840
		x"1f",	--2841
		x"20",	--2842
		x"b0",	--2843
		x"24",	--2844
		x"0a",	--2845
		x"0b",	--2846
		x"1f",	--2847
		x"1e",	--2848
		x"b0",	--2849
		x"24",	--2850
		x"0c",	--2851
		x"0d",	--2852
		x"3c",	--2853
		x"3d",	--2854
		x"1c",	--2855
		x"0d",	--2856
		x"0d",	--2857
		x"0c",	--2858
		x"0d",	--2859
		x"0e",	--2860
		x"0f",	--2861
		x"b0",	--2862
		x"b0",	--2863
		x"21",	--2864
		x"39",	--2865
		x"3a",	--2866
		x"3b",	--2867
		x"30",	--2868
		x"0d",	--2869
		x"1f",	--2870
		x"22",	--2871
		x"b0",	--2872
		x"48",	--2873
		x"30",	--2874
		x"1f",	--2875
		x"22",	--2876
		x"b0",	--2877
		x"70",	--2878
		x"30",	--2879
		x"0b",	--2880
		x"0a",	--2881
		x"0b",	--2882
		x"0a",	--2883
		x"8f",	--2884
		x"00",	--2885
		x"8f",	--2886
		x"02",	--2887
		x"8f",	--2888
		x"04",	--2889
		x"0c",	--2890
		x"0d",	--2891
		x"3e",	--2892
		x"00",	--2893
		x"3f",	--2894
		x"6e",	--2895
		x"b0",	--2896
		x"f8",	--2897
		x"8b",	--2898
		x"02",	--2899
		x"02",	--2900
		x"32",	--2901
		x"03",	--2902
		x"82",	--2903
		x"32",	--2904
		x"b2",	--2905
		x"18",	--2906
		x"38",	--2907
		x"9b",	--2908
		x"3a",	--2909
		x"06",	--2910
		x"32",	--2911
		x"0f",	--2912
		x"3a",	--2913
		x"3b",	--2914
		x"30",	--2915
		x"0b",	--2916
		x"09",	--2917
		x"08",	--2918
		x"8f",	--2919
		x"06",	--2920
		x"bf",	--2921
		x"00",	--2922
		x"08",	--2923
		x"2b",	--2924
		x"1e",	--2925
		x"02",	--2926
		x"0f",	--2927
		x"b0",	--2928
		x"92",	--2929
		x"0c",	--2930
		x"3d",	--2931
		x"00",	--2932
		x"b0",	--2933
		x"58",	--2934
		x"08",	--2935
		x"09",	--2936
		x"1e",	--2937
		x"06",	--2938
		x"0f",	--2939
		x"b0",	--2940
		x"92",	--2941
		x"0c",	--2942
		x"0d",	--2943
		x"0e",	--2944
		x"0f",	--2945
		x"b0",	--2946
		x"08",	--2947
		x"b0",	--2948
		x"e8",	--2949
		x"8b",	--2950
		x"04",	--2951
		x"9b",	--2952
		x"00",	--2953
		x"38",	--2954
		x"39",	--2955
		x"3b",	--2956
		x"30",	--2957
		x"0b",	--2958
		x"0a",	--2959
		x"09",	--2960
		x"0a",	--2961
		x"0b",	--2962
		x"8f",	--2963
		x"06",	--2964
		x"8f",	--2965
		x"08",	--2966
		x"29",	--2967
		x"1e",	--2968
		x"02",	--2969
		x"0f",	--2970
		x"b0",	--2971
		x"92",	--2972
		x"0c",	--2973
		x"0d",	--2974
		x"0e",	--2975
		x"0f",	--2976
		x"b0",	--2977
		x"58",	--2978
		x"0a",	--2979
		x"0b",	--2980
		x"1e",	--2981
		x"06",	--2982
		x"0f",	--2983
		x"b0",	--2984
		x"92",	--2985
		x"0c",	--2986
		x"0d",	--2987
		x"0e",	--2988
		x"0f",	--2989
		x"b0",	--2990
		x"08",	--2991
		x"b0",	--2992
		x"e8",	--2993
		x"89",	--2994
		x"04",	--2995
		x"39",	--2996
		x"3a",	--2997
		x"3b",	--2998
		x"30",	--2999
		x"2f",	--3000
		x"8f",	--3001
		x"04",	--3002
		x"30",	--3003
		x"0b",	--3004
		x"0a",	--3005
		x"92",	--3006
		x"40",	--3007
		x"14",	--3008
		x"3b",	--3009
		x"90",	--3010
		x"0a",	--3011
		x"2b",	--3012
		x"5f",	--3013
		x"fc",	--3014
		x"8f",	--3015
		x"0f",	--3016
		x"30",	--3017
		x"7c",	--3018
		x"b0",	--3019
		x"3a",	--3020
		x"31",	--3021
		x"06",	--3022
		x"1a",	--3023
		x"3b",	--3024
		x"06",	--3025
		x"1a",	--3026
		x"40",	--3027
		x"ef",	--3028
		x"0f",	--3029
		x"3a",	--3030
		x"3b",	--3031
		x"30",	--3032
		x"1e",	--3033
		x"40",	--3034
		x"3e",	--3035
		x"20",	--3036
		x"12",	--3037
		x"0f",	--3038
		x"0f",	--3039
		x"0f",	--3040
		x"0f",	--3041
		x"3f",	--3042
		x"8c",	--3043
		x"ff",	--3044
		x"68",	--3045
		x"00",	--3046
		x"bf",	--3047
		x"78",	--3048
		x"02",	--3049
		x"bf",	--3050
		x"08",	--3051
		x"04",	--3052
		x"1e",	--3053
		x"82",	--3054
		x"40",	--3055
		x"30",	--3056
		x"0b",	--3057
		x"1b",	--3058
		x"40",	--3059
		x"3b",	--3060
		x"20",	--3061
		x"12",	--3062
		x"0c",	--3063
		x"0c",	--3064
		x"0c",	--3065
		x"0c",	--3066
		x"3c",	--3067
		x"8c",	--3068
		x"cc",	--3069
		x"00",	--3070
		x"8c",	--3071
		x"02",	--3072
		x"8c",	--3073
		x"04",	--3074
		x"1b",	--3075
		x"82",	--3076
		x"40",	--3077
		x"0f",	--3078
		x"3b",	--3079
		x"30",	--3080
		x"3f",	--3081
		x"fc",	--3082
		x"0b",	--3083
		x"31",	--3084
		x"f0",	--3085
		x"1b",	--3086
		x"40",	--3087
		x"1b",	--3088
		x"0f",	--3089
		x"5f",	--3090
		x"8c",	--3091
		x"16",	--3092
		x"3d",	--3093
		x"92",	--3094
		x"0c",	--3095
		x"05",	--3096
		x"3d",	--3097
		x"06",	--3098
		x"cd",	--3099
		x"fa",	--3100
		x"0e",	--3101
		x"1c",	--3102
		x"0c",	--3103
		x"f8",	--3104
		x"30",	--3105
		x"84",	--3106
		x"b0",	--3107
		x"3a",	--3108
		x"21",	--3109
		x"3f",	--3110
		x"31",	--3111
		x"10",	--3112
		x"3b",	--3113
		x"30",	--3114
		x"0c",	--3115
		x"81",	--3116
		x"00",	--3117
		x"6d",	--3118
		x"4d",	--3119
		x"24",	--3120
		x"1e",	--3121
		x"1f",	--3122
		x"06",	--3123
		x"6d",	--3124
		x"4d",	--3125
		x"11",	--3126
		x"1e",	--3127
		x"3f",	--3128
		x"0e",	--3129
		x"7d",	--3130
		x"20",	--3131
		x"f7",	--3132
		x"ce",	--3133
		x"ff",	--3134
		x"0d",	--3135
		x"0d",	--3136
		x"0d",	--3137
		x"8d",	--3138
		x"00",	--3139
		x"1f",	--3140
		x"6d",	--3141
		x"4d",	--3142
		x"ef",	--3143
		x"0e",	--3144
		x"0e",	--3145
		x"0c",	--3146
		x"0c",	--3147
		x"3c",	--3148
		x"8c",	--3149
		x"0e",	--3150
		x"9c",	--3151
		x"02",	--3152
		x"31",	--3153
		x"10",	--3154
		x"3b",	--3155
		x"30",	--3156
		x"1f",	--3157
		x"f1",	--3158
		x"8f",	--3159
		x"00",	--3160
		x"0f",	--3161
		x"30",	--3162
		x"0e",	--3163
		x"2e",	--3164
		x"2f",	--3165
		x"30",	--3166
		x"0b",	--3167
		x"0a",	--3168
		x"0e",	--3169
		x"2e",	--3170
		x"2c",	--3171
		x"0d",	--3172
		x"0e",	--3173
		x"0f",	--3174
		x"0e",	--3175
		x"0f",	--3176
		x"0a",	--3177
		x"0b",	--3178
		x"0a",	--3179
		x"0b",	--3180
		x"0a",	--3181
		x"0b",	--3182
		x"3c",	--3183
		x"3a",	--3184
		x"0d",	--3185
		x"0e",	--3186
		x"0f",	--3187
		x"b0",	--3188
		x"b8",	--3189
		x"0f",	--3190
		x"3a",	--3191
		x"3b",	--3192
		x"30",	--3193
		x"b2",	--3194
		x"d2",	--3195
		x"60",	--3196
		x"b2",	--3197
		x"b8",	--3198
		x"72",	--3199
		x"0f",	--3200
		x"30",	--3201
		x"0b",	--3202
		x"0b",	--3203
		x"1f",	--3204
		x"42",	--3205
		x"3f",	--3206
		x"20",	--3207
		x"19",	--3208
		x"0c",	--3209
		x"0c",	--3210
		x"0d",	--3211
		x"0d",	--3212
		x"0d",	--3213
		x"0d",	--3214
		x"0d",	--3215
		x"3d",	--3216
		x"4c",	--3217
		x"8d",	--3218
		x"00",	--3219
		x"8d",	--3220
		x"02",	--3221
		x"8d",	--3222
		x"08",	--3223
		x"8d",	--3224
		x"0a",	--3225
		x"8d",	--3226
		x"0c",	--3227
		x"0e",	--3228
		x"1e",	--3229
		x"82",	--3230
		x"42",	--3231
		x"3b",	--3232
		x"30",	--3233
		x"3f",	--3234
		x"fc",	--3235
		x"0f",	--3236
		x"0c",	--3237
		x"0c",	--3238
		x"0c",	--3239
		x"0c",	--3240
		x"0c",	--3241
		x"3c",	--3242
		x"4c",	--3243
		x"8c",	--3244
		x"02",	--3245
		x"8c",	--3246
		x"04",	--3247
		x"8c",	--3248
		x"06",	--3249
		x"8c",	--3250
		x"08",	--3251
		x"9c",	--3252
		x"00",	--3253
		x"0f",	--3254
		x"30",	--3255
		x"0f",	--3256
		x"0e",	--3257
		x"0e",	--3258
		x"0e",	--3259
		x"0e",	--3260
		x"0e",	--3261
		x"8e",	--3262
		x"4c",	--3263
		x"0f",	--3264
		x"30",	--3265
		x"0f",	--3266
		x"0e",	--3267
		x"0d",	--3268
		x"0c",	--3269
		x"0b",	--3270
		x"0a",	--3271
		x"09",	--3272
		x"08",	--3273
		x"07",	--3274
		x"92",	--3275
		x"42",	--3276
		x"33",	--3277
		x"3a",	--3278
		x"4c",	--3279
		x"0b",	--3280
		x"2b",	--3281
		x"08",	--3282
		x"38",	--3283
		x"07",	--3284
		x"37",	--3285
		x"06",	--3286
		x"09",	--3287
		x"0f",	--3288
		x"1f",	--3289
		x"8b",	--3290
		x"00",	--3291
		x"19",	--3292
		x"3a",	--3293
		x"0e",	--3294
		x"3b",	--3295
		x"0e",	--3296
		x"38",	--3297
		x"0e",	--3298
		x"37",	--3299
		x"0e",	--3300
		x"19",	--3301
		x"42",	--3302
		x"19",	--3303
		x"8a",	--3304
		x"00",	--3305
		x"f1",	--3306
		x"2f",	--3307
		x"1f",	--3308
		x"02",	--3309
		x"ea",	--3310
		x"8b",	--3311
		x"00",	--3312
		x"1f",	--3313
		x"0a",	--3314
		x"9b",	--3315
		x"08",	--3316
		x"88",	--3317
		x"00",	--3318
		x"e4",	--3319
		x"2f",	--3320
		x"1f",	--3321
		x"87",	--3322
		x"00",	--3323
		x"2f",	--3324
		x"de",	--3325
		x"8a",	--3326
		x"00",	--3327
		x"db",	--3328
		x"b2",	--3329
		x"fe",	--3330
		x"60",	--3331
		x"37",	--3332
		x"38",	--3333
		x"39",	--3334
		x"3a",	--3335
		x"3b",	--3336
		x"3c",	--3337
		x"3d",	--3338
		x"3e",	--3339
		x"3f",	--3340
		x"00",	--3341
		x"8f",	--3342
		x"00",	--3343
		x"0f",	--3344
		x"30",	--3345
		x"2f",	--3346
		x"2e",	--3347
		x"1f",	--3348
		x"02",	--3349
		x"30",	--3350
		x"8f",	--3351
		x"00",	--3352
		x"30",	--3353
		x"8f",	--3354
		x"00",	--3355
		x"3f",	--3356
		x"2e",	--3357
		x"b0",	--3358
		x"04",	--3359
		x"82",	--3360
		x"0e",	--3361
		x"0f",	--3362
		x"30",	--3363
		x"0c",	--3364
		x"2f",	--3365
		x"8f",	--3366
		x"00",	--3367
		x"1d",	--3368
		x"0e",	--3369
		x"1f",	--3370
		x"0e",	--3371
		x"b0",	--3372
		x"48",	--3373
		x"30",	--3374
		x"5e",	--3375
		x"81",	--3376
		x"3e",	--3377
		x"fc",	--3378
		x"c2",	--3379
		x"84",	--3380
		x"0f",	--3381
		x"30",	--3382
		x"3f",	--3383
		x"0f",	--3384
		x"5f",	--3385
		x"42",	--3386
		x"8f",	--3387
		x"b0",	--3388
		x"5e",	--3389
		x"30",	--3390
		x"0b",	--3391
		x"0b",	--3392
		x"0e",	--3393
		x"0e",	--3394
		x"0e",	--3395
		x"0e",	--3396
		x"0e",	--3397
		x"0f",	--3398
		x"b0",	--3399
		x"6e",	--3400
		x"0f",	--3401
		x"b0",	--3402
		x"6e",	--3403
		x"3b",	--3404
		x"30",	--3405
		x"0b",	--3406
		x"0a",	--3407
		x"0a",	--3408
		x"3b",	--3409
		x"07",	--3410
		x"0e",	--3411
		x"4d",	--3412
		x"7d",	--3413
		x"0f",	--3414
		x"03",	--3415
		x"0e",	--3416
		x"7d",	--3417
		x"fd",	--3418
		x"1e",	--3419
		x"0a",	--3420
		x"3f",	--3421
		x"31",	--3422
		x"b0",	--3423
		x"5e",	--3424
		x"3b",	--3425
		x"3b",	--3426
		x"ef",	--3427
		x"3a",	--3428
		x"3b",	--3429
		x"30",	--3430
		x"3f",	--3431
		x"30",	--3432
		x"f5",	--3433
		x"0b",	--3434
		x"0b",	--3435
		x"0e",	--3436
		x"8e",	--3437
		x"8e",	--3438
		x"0f",	--3439
		x"b0",	--3440
		x"7e",	--3441
		x"0f",	--3442
		x"b0",	--3443
		x"7e",	--3444
		x"3b",	--3445
		x"30",	--3446
		x"0b",	--3447
		x"0a",	--3448
		x"0a",	--3449
		x"0b",	--3450
		x"0d",	--3451
		x"8d",	--3452
		x"8d",	--3453
		x"0f",	--3454
		x"b0",	--3455
		x"7e",	--3456
		x"0f",	--3457
		x"b0",	--3458
		x"7e",	--3459
		x"0c",	--3460
		x"0d",	--3461
		x"8d",	--3462
		x"8c",	--3463
		x"4d",	--3464
		x"0d",	--3465
		x"0f",	--3466
		x"b0",	--3467
		x"7e",	--3468
		x"0f",	--3469
		x"b0",	--3470
		x"7e",	--3471
		x"3a",	--3472
		x"3b",	--3473
		x"30",	--3474
		x"0b",	--3475
		x"0a",	--3476
		x"09",	--3477
		x"0a",	--3478
		x"0e",	--3479
		x"19",	--3480
		x"09",	--3481
		x"39",	--3482
		x"0b",	--3483
		x"0d",	--3484
		x"0d",	--3485
		x"6f",	--3486
		x"8f",	--3487
		x"b0",	--3488
		x"7e",	--3489
		x"0b",	--3490
		x"0e",	--3491
		x"1b",	--3492
		x"3b",	--3493
		x"07",	--3494
		x"05",	--3495
		x"3f",	--3496
		x"20",	--3497
		x"b0",	--3498
		x"5e",	--3499
		x"ef",	--3500
		x"3f",	--3501
		x"3a",	--3502
		x"b0",	--3503
		x"5e",	--3504
		x"ea",	--3505
		x"39",	--3506
		x"3a",	--3507
		x"3b",	--3508
		x"30",	--3509
		x"0b",	--3510
		x"0a",	--3511
		x"09",	--3512
		x"0a",	--3513
		x"0e",	--3514
		x"17",	--3515
		x"09",	--3516
		x"39",	--3517
		x"0b",	--3518
		x"6f",	--3519
		x"8f",	--3520
		x"b0",	--3521
		x"6e",	--3522
		x"0b",	--3523
		x"0e",	--3524
		x"1b",	--3525
		x"3b",	--3526
		x"07",	--3527
		x"f6",	--3528
		x"3f",	--3529
		x"20",	--3530
		x"b0",	--3531
		x"5e",	--3532
		x"6f",	--3533
		x"8f",	--3534
		x"b0",	--3535
		x"6e",	--3536
		x"0b",	--3537
		x"f2",	--3538
		x"39",	--3539
		x"3a",	--3540
		x"3b",	--3541
		x"30",	--3542
		x"0b",	--3543
		x"0a",	--3544
		x"09",	--3545
		x"31",	--3546
		x"ec",	--3547
		x"0b",	--3548
		x"0f",	--3549
		x"34",	--3550
		x"3b",	--3551
		x"0a",	--3552
		x"38",	--3553
		x"09",	--3554
		x"0a",	--3555
		x"0a",	--3556
		x"3e",	--3557
		x"0a",	--3558
		x"0f",	--3559
		x"b0",	--3560
		x"b0",	--3561
		x"7f",	--3562
		x"30",	--3563
		x"ca",	--3564
		x"00",	--3565
		x"19",	--3566
		x"3e",	--3567
		x"0a",	--3568
		x"0f",	--3569
		x"b0",	--3570
		x"7e",	--3571
		x"0b",	--3572
		x"3f",	--3573
		x"0a",	--3574
		x"eb",	--3575
		x"0a",	--3576
		x"1a",	--3577
		x"09",	--3578
		x"3e",	--3579
		x"0a",	--3580
		x"0f",	--3581
		x"b0",	--3582
		x"b0",	--3583
		x"7f",	--3584
		x"30",	--3585
		x"c9",	--3586
		x"00",	--3587
		x"3a",	--3588
		x"0f",	--3589
		x"0f",	--3590
		x"6f",	--3591
		x"8f",	--3592
		x"b0",	--3593
		x"5e",	--3594
		x"0a",	--3595
		x"f7",	--3596
		x"31",	--3597
		x"14",	--3598
		x"39",	--3599
		x"3a",	--3600
		x"3b",	--3601
		x"30",	--3602
		x"3f",	--3603
		x"2d",	--3604
		x"b0",	--3605
		x"5e",	--3606
		x"3b",	--3607
		x"1b",	--3608
		x"c5",	--3609
		x"1a",	--3610
		x"09",	--3611
		x"dd",	--3612
		x"0b",	--3613
		x"0a",	--3614
		x"09",	--3615
		x"0b",	--3616
		x"3b",	--3617
		x"39",	--3618
		x"6f",	--3619
		x"4f",	--3620
		x"0b",	--3621
		x"1a",	--3622
		x"8f",	--3623
		x"b0",	--3624
		x"5e",	--3625
		x"0a",	--3626
		x"09",	--3627
		x"19",	--3628
		x"5f",	--3629
		x"01",	--3630
		x"4f",	--3631
		x"10",	--3632
		x"7f",	--3633
		x"25",	--3634
		x"f3",	--3635
		x"0a",	--3636
		x"1a",	--3637
		x"5f",	--3638
		x"01",	--3639
		x"7f",	--3640
		x"db",	--3641
		x"7f",	--3642
		x"54",	--3643
		x"ee",	--3644
		x"4f",	--3645
		x"0f",	--3646
		x"10",	--3647
		x"9a",	--3648
		x"39",	--3649
		x"3a",	--3650
		x"3b",	--3651
		x"30",	--3652
		x"09",	--3653
		x"29",	--3654
		x"1e",	--3655
		x"02",	--3656
		x"2f",	--3657
		x"b0",	--3658
		x"26",	--3659
		x"0b",	--3660
		x"dd",	--3661
		x"09",	--3662
		x"29",	--3663
		x"2f",	--3664
		x"b0",	--3665
		x"d4",	--3666
		x"0b",	--3667
		x"d6",	--3668
		x"0f",	--3669
		x"2b",	--3670
		x"29",	--3671
		x"6f",	--3672
		x"4f",	--3673
		x"d0",	--3674
		x"19",	--3675
		x"8f",	--3676
		x"b0",	--3677
		x"5e",	--3678
		x"7f",	--3679
		x"4f",	--3680
		x"fa",	--3681
		x"c8",	--3682
		x"09",	--3683
		x"29",	--3684
		x"1e",	--3685
		x"02",	--3686
		x"2f",	--3687
		x"b0",	--3688
		x"6c",	--3689
		x"0b",	--3690
		x"bf",	--3691
		x"09",	--3692
		x"29",	--3693
		x"2e",	--3694
		x"0f",	--3695
		x"8f",	--3696
		x"8f",	--3697
		x"8f",	--3698
		x"8f",	--3699
		x"b0",	--3700
		x"ee",	--3701
		x"0b",	--3702
		x"b3",	--3703
		x"09",	--3704
		x"29",	--3705
		x"2f",	--3706
		x"b0",	--3707
		x"ae",	--3708
		x"0b",	--3709
		x"ac",	--3710
		x"09",	--3711
		x"29",	--3712
		x"2f",	--3713
		x"b0",	--3714
		x"5e",	--3715
		x"0b",	--3716
		x"a5",	--3717
		x"09",	--3718
		x"29",	--3719
		x"2f",	--3720
		x"b0",	--3721
		x"7e",	--3722
		x"0b",	--3723
		x"9e",	--3724
		x"09",	--3725
		x"29",	--3726
		x"2f",	--3727
		x"b0",	--3728
		x"9c",	--3729
		x"0b",	--3730
		x"97",	--3731
		x"3f",	--3732
		x"25",	--3733
		x"b0",	--3734
		x"5e",	--3735
		x"92",	--3736
		x"0f",	--3737
		x"0e",	--3738
		x"1f",	--3739
		x"44",	--3740
		x"df",	--3741
		x"85",	--3742
		x"0c",	--3743
		x"1f",	--3744
		x"44",	--3745
		x"3f",	--3746
		x"3f",	--3747
		x"13",	--3748
		x"92",	--3749
		x"44",	--3750
		x"1e",	--3751
		x"44",	--3752
		x"1f",	--3753
		x"46",	--3754
		x"0e",	--3755
		x"02",	--3756
		x"92",	--3757
		x"46",	--3758
		x"f2",	--3759
		x"10",	--3760
		x"81",	--3761
		x"3e",	--3762
		x"3f",	--3763
		x"b1",	--3764
		x"f0",	--3765
		x"00",	--3766
		x"00",	--3767
		x"82",	--3768
		x"44",	--3769
		x"ec",	--3770
		x"0c",	--3771
		x"0d",	--3772
		x"3e",	--3773
		x"00",	--3774
		x"3f",	--3775
		x"6e",	--3776
		x"b0",	--3777
		x"b8",	--3778
		x"3e",	--3779
		x"82",	--3780
		x"82",	--3781
		x"f2",	--3782
		x"11",	--3783
		x"80",	--3784
		x"30",	--3785
		x"1e",	--3786
		x"44",	--3787
		x"1f",	--3788
		x"46",	--3789
		x"0e",	--3790
		x"05",	--3791
		x"1f",	--3792
		x"44",	--3793
		x"1f",	--3794
		x"46",	--3795
		x"30",	--3796
		x"1d",	--3797
		x"44",	--3798
		x"1e",	--3799
		x"46",	--3800
		x"3f",	--3801
		x"40",	--3802
		x"0f",	--3803
		x"0f",	--3804
		x"30",	--3805
		x"1f",	--3806
		x"46",	--3807
		x"5f",	--3808
		x"0c",	--3809
		x"1d",	--3810
		x"46",	--3811
		x"1e",	--3812
		x"44",	--3813
		x"0d",	--3814
		x"0b",	--3815
		x"1e",	--3816
		x"46",	--3817
		x"3e",	--3818
		x"3f",	--3819
		x"03",	--3820
		x"82",	--3821
		x"46",	--3822
		x"30",	--3823
		x"92",	--3824
		x"46",	--3825
		x"30",	--3826
		x"4f",	--3827
		x"30",	--3828
		x"0b",	--3829
		x"0a",	--3830
		x"09",	--3831
		x"08",	--3832
		x"07",	--3833
		x"06",	--3834
		x"05",	--3835
		x"04",	--3836
		x"31",	--3837
		x"04",	--3838
		x"05",	--3839
		x"81",	--3840
		x"00",	--3841
		x"81",	--3842
		x"02",	--3843
		x"08",	--3844
		x"09",	--3845
		x"38",	--3846
		x"39",	--3847
		x"ff",	--3848
		x"39",	--3849
		x"80",	--3850
		x"1f",	--3851
		x"39",	--3852
		x"80",	--3853
		x"0b",	--3854
		x"02",	--3855
		x"18",	--3856
		x"08",	--3857
		x"0c",	--3858
		x"0d",	--3859
		x"0e",	--3860
		x"0f",	--3861
		x"b0",	--3862
		x"bc",	--3863
		x"30",	--3864
		x"be",	--3865
		x"81",	--3866
		x"02",	--3867
		x"02",	--3868
		x"30",	--3869
		x"1e",	--3870
		x"05",	--3871
		x"91",	--3872
		x"00",	--3873
		x"02",	--3874
		x"30",	--3875
		x"1e",	--3876
		x"34",	--3877
		x"db",	--3878
		x"35",	--3879
		x"c9",	--3880
		x"30",	--3881
		x"26",	--3882
		x"39",	--3883
		x"e0",	--3884
		x"08",	--3885
		x"0a",	--3886
		x"0b",	--3887
		x"3b",	--3888
		x"ff",	--3889
		x"39",	--3890
		x"98",	--3891
		x"1b",	--3892
		x"16",	--3893
		x"39",	--3894
		x"00",	--3895
		x"10",	--3896
		x"3c",	--3897
		x"ca",	--3898
		x"3d",	--3899
		x"49",	--3900
		x"b0",	--3901
		x"bc",	--3902
		x"0c",	--3903
		x"3d",	--3904
		x"80",	--3905
		x"b0",	--3906
		x"1c",	--3907
		x"0f",	--3908
		x"03",	--3909
		x"02",	--3910
		x"30",	--3911
		x"26",	--3912
		x"36",	--3913
		x"37",	--3914
		x"6d",	--3915
		x"39",	--3916
		x"1c",	--3917
		x"4b",	--3918
		x"3d",	--3919
		x"39",	--3920
		x"30",	--3921
		x"1b",	--3922
		x"0c",	--3923
		x"3d",	--3924
		x"80",	--3925
		x"0e",	--3926
		x"0f",	--3927
		x"b0",	--3928
		x"08",	--3929
		x"08",	--3930
		x"09",	--3931
		x"0c",	--3932
		x"3d",	--3933
		x"80",	--3934
		x"0e",	--3935
		x"0f",	--3936
		x"b0",	--3937
		x"bc",	--3938
		x"0c",	--3939
		x"0d",	--3940
		x"0e",	--3941
		x"0f",	--3942
		x"b0",	--3943
		x"7c",	--3944
		x"04",	--3945
		x"05",	--3946
		x"16",	--3947
		x"07",	--3948
		x"4b",	--3949
		x"0c",	--3950
		x"0d",	--3951
		x"0e",	--3952
		x"0f",	--3953
		x"b0",	--3954
		x"bc",	--3955
		x"0c",	--3956
		x"3d",	--3957
		x"80",	--3958
		x"b0",	--3959
		x"08",	--3960
		x"08",	--3961
		x"09",	--3962
		x"0c",	--3963
		x"3d",	--3964
		x"00",	--3965
		x"0e",	--3966
		x"0f",	--3967
		x"b0",	--3968
		x"bc",	--3969
		x"0c",	--3970
		x"0d",	--3971
		x"0e",	--3972
		x"0f",	--3973
		x"b0",	--3974
		x"7c",	--3975
		x"04",	--3976
		x"05",	--3977
		x"06",	--3978
		x"07",	--3979
		x"2c",	--3980
		x"0c",	--3981
		x"0d",	--3982
		x"0e",	--3983
		x"3f",	--3984
		x"80",	--3985
		x"b0",	--3986
		x"7c",	--3987
		x"04",	--3988
		x"05",	--3989
		x"36",	--3990
		x"03",	--3991
		x"07",	--3992
		x"1f",	--3993
		x"0c",	--3994
		x"3d",	--3995
		x"c0",	--3996
		x"0e",	--3997
		x"0f",	--3998
		x"b0",	--3999
		x"08",	--4000
		x"08",	--4001
		x"09",	--4002
		x"0c",	--4003
		x"3d",	--4004
		x"c0",	--4005
		x"0e",	--4006
		x"0f",	--4007
		x"b0",	--4008
		x"58",	--4009
		x"0c",	--4010
		x"3d",	--4011
		x"80",	--4012
		x"b0",	--4013
		x"bc",	--4014
		x"0c",	--4015
		x"0d",	--4016
		x"0e",	--4017
		x"0f",	--4018
		x"b0",	--4019
		x"7c",	--4020
		x"04",	--4021
		x"05",	--4022
		x"26",	--4023
		x"07",	--4024
		x"0c",	--4025
		x"0d",	--4026
		x"0e",	--4027
		x"0f",	--4028
		x"b0",	--4029
		x"58",	--4030
		x"08",	--4031
		x"09",	--4032
		x"0c",	--4033
		x"0d",	--4034
		x"b0",	--4035
		x"58",	--4036
		x"0a",	--4037
		x"0b",	--4038
		x"3c",	--4039
		x"d7",	--4040
		x"3d",	--4041
		x"85",	--4042
		x"b0",	--4043
		x"58",	--4044
		x"3c",	--4045
		x"59",	--4046
		x"3d",	--4047
		x"4b",	--4048
		x"b0",	--4049
		x"bc",	--4050
		x"0c",	--4051
		x"0d",	--4052
		x"0e",	--4053
		x"0f",	--4054
		x"b0",	--4055
		x"58",	--4056
		x"3c",	--4057
		x"35",	--4058
		x"3d",	--4059
		x"88",	--4060
		x"b0",	--4061
		x"bc",	--4062
		x"0c",	--4063
		x"0d",	--4064
		x"0e",	--4065
		x"0f",	--4066
		x"b0",	--4067
		x"58",	--4068
		x"3c",	--4069
		x"6e",	--4070
		x"3d",	--4071
		x"ba",	--4072
		x"b0",	--4073
		x"bc",	--4074
		x"0c",	--4075
		x"0d",	--4076
		x"0e",	--4077
		x"0f",	--4078
		x"b0",	--4079
		x"58",	--4080
		x"3c",	--4081
		x"25",	--4082
		x"3d",	--4083
		x"12",	--4084
		x"b0",	--4085
		x"bc",	--4086
		x"0c",	--4087
		x"0d",	--4088
		x"0e",	--4089
		x"0f",	--4090
		x"b0",	--4091
		x"58",	--4092
		x"3c",	--4093
		x"ab",	--4094
		x"3d",	--4095
		x"aa",	--4096
		x"b0",	--4097
		x"bc",	--4098
		x"0c",	--4099
		x"0d",	--4100
		x"0e",	--4101
		x"0f",	--4102
		x"b0",	--4103
		x"58",	--4104
		x"81",	--4105
		x"04",	--4106
		x"81",	--4107
		x"06",	--4108
		x"3c",	--4109
		x"21",	--4110
		x"3d",	--4111
		x"15",	--4112
		x"0e",	--4113
		x"0f",	--4114
		x"b0",	--4115
		x"58",	--4116
		x"3c",	--4117
		x"6b",	--4118
		x"3d",	--4119
		x"6e",	--4120
		x"b0",	--4121
		x"08",	--4122
		x"0c",	--4123
		x"0d",	--4124
		x"0e",	--4125
		x"0f",	--4126
		x"b0",	--4127
		x"58",	--4128
		x"3c",	--4129
		x"95",	--4130
		x"3d",	--4131
		x"9d",	--4132
		x"b0",	--4133
		x"08",	--4134
		x"0c",	--4135
		x"0d",	--4136
		x"0e",	--4137
		x"0f",	--4138
		x"b0",	--4139
		x"58",	--4140
		x"3c",	--4141
		x"38",	--4142
		x"3d",	--4143
		x"e3",	--4144
		x"b0",	--4145
		x"08",	--4146
		x"0c",	--4147
		x"0d",	--4148
		x"0e",	--4149
		x"0f",	--4150
		x"b0",	--4151
		x"58",	--4152
		x"3c",	--4153
		x"cd",	--4154
		x"3d",	--4155
		x"4c",	--4156
		x"b0",	--4157
		x"08",	--4158
		x"0c",	--4159
		x"0d",	--4160
		x"0e",	--4161
		x"0f",	--4162
		x"b0",	--4163
		x"58",	--4164
		x"08",	--4165
		x"09",	--4166
		x"36",	--4167
		x"19",	--4168
		x"37",	--4169
		x"17",	--4170
		x"0c",	--4171
		x"0d",	--4172
		x"1e",	--4173
		x"04",	--4174
		x"1f",	--4175
		x"06",	--4176
		x"b0",	--4177
		x"bc",	--4178
		x"0c",	--4179
		x"0d",	--4180
		x"0e",	--4181
		x"0f",	--4182
		x"b0",	--4183
		x"58",	--4184
		x"0c",	--4185
		x"0d",	--4186
		x"0e",	--4187
		x"0f",	--4188
		x"b0",	--4189
		x"08",	--4190
		x"04",	--4191
		x"05",	--4192
		x"31",	--4193
		x"0b",	--4194
		x"0b",	--4195
		x"0b",	--4196
		x"07",	--4197
		x"37",	--4198
		x"54",	--4199
		x"0c",	--4200
		x"0d",	--4201
		x"1e",	--4202
		x"04",	--4203
		x"1f",	--4204
		x"06",	--4205
		x"b0",	--4206
		x"bc",	--4207
		x"0c",	--4208
		x"0d",	--4209
		x"0e",	--4210
		x"0f",	--4211
		x"b0",	--4212
		x"58",	--4213
		x"1c",	--4214
		x"64",	--4215
		x"1d",	--4216
		x"66",	--4217
		x"b0",	--4218
		x"08",	--4219
		x"0c",	--4220
		x"0d",	--4221
		x"b0",	--4222
		x"08",	--4223
		x"0c",	--4224
		x"0d",	--4225
		x"2e",	--4226
		x"1f",	--4227
		x"02",	--4228
		x"b0",	--4229
		x"08",	--4230
		x"04",	--4231
		x"05",	--4232
		x"81",	--4233
		x"02",	--4234
		x"07",	--4235
		x"35",	--4236
		x"00",	--4237
		x"04",	--4238
		x"34",	--4239
		x"db",	--4240
		x"35",	--4241
		x"c9",	--4242
		x"0e",	--4243
		x"0f",	--4244
		x"31",	--4245
		x"34",	--4246
		x"35",	--4247
		x"36",	--4248
		x"37",	--4249
		x"38",	--4250
		x"39",	--4251
		x"3a",	--4252
		x"3b",	--4253
		x"30",	--4254
		x"b0",	--4255
		x"ea",	--4256
		x"30",	--4257
		x"0b",	--4258
		x"0a",	--4259
		x"31",	--4260
		x"0c",	--4261
		x"0d",	--4262
		x"3c",	--4263
		x"3d",	--4264
		x"ff",	--4265
		x"3d",	--4266
		x"49",	--4267
		x"06",	--4268
		x"3d",	--4269
		x"4a",	--4270
		x"07",	--4271
		x"3c",	--4272
		x"d9",	--4273
		x"04",	--4274
		x"03",	--4275
		x"0c",	--4276
		x"0d",	--4277
		x"27",	--4278
		x"3d",	--4279
		x"80",	--4280
		x"05",	--4281
		x"0c",	--4282
		x"0d",	--4283
		x"b0",	--4284
		x"08",	--4285
		x"2f",	--4286
		x"0d",	--4287
		x"b0",	--4288
		x"ce",	--4289
		x"0a",	--4290
		x"0b",	--4291
		x"3a",	--4292
		x"03",	--4293
		x"0b",	--4294
		x"1c",	--4295
		x"04",	--4296
		x"1d",	--4297
		x"06",	--4298
		x"2e",	--4299
		x"1f",	--4300
		x"02",	--4301
		x"1a",	--4302
		x"02",	--4303
		x"0b",	--4304
		x"10",	--4305
		x"2a",	--4306
		x"02",	--4307
		x"0b",	--4308
		x"0f",	--4309
		x"2e",	--4310
		x"1f",	--4311
		x"02",	--4312
		x"0a",	--4313
		x"0f",	--4314
		x"0b",	--4315
		x"0d",	--4316
		x"13",	--4317
		x"b0",	--4318
		x"c4",	--4319
		x"21",	--4320
		x"0c",	--4321
		x"b0",	--4322
		x"ea",	--4323
		x"09",	--4324
		x"13",	--4325
		x"b0",	--4326
		x"c4",	--4327
		x"21",	--4328
		x"02",	--4329
		x"b0",	--4330
		x"ea",	--4331
		x"3f",	--4332
		x"00",	--4333
		x"31",	--4334
		x"3a",	--4335
		x"3b",	--4336
		x"30",	--4337
		x"b0",	--4338
		x"44",	--4339
		x"30",	--4340
		x"0b",	--4341
		x"0a",	--4342
		x"09",	--4343
		x"08",	--4344
		x"07",	--4345
		x"06",	--4346
		x"05",	--4347
		x"04",	--4348
		x"31",	--4349
		x"06",	--4350
		x"07",	--4351
		x"04",	--4352
		x"05",	--4353
		x"0a",	--4354
		x"0b",	--4355
		x"3a",	--4356
		x"3b",	--4357
		x"ff",	--4358
		x"3b",	--4359
		x"00",	--4360
		x"04",	--4361
		x"b0",	--4362
		x"02",	--4363
		x"0e",	--4364
		x"cc",	--4365
		x"0c",	--4366
		x"0d",	--4367
		x"0e",	--4368
		x"0f",	--4369
		x"b0",	--4370
		x"58",	--4371
		x"08",	--4372
		x"09",	--4373
		x"3c",	--4374
		x"4e",	--4375
		x"3d",	--4376
		x"47",	--4377
		x"b0",	--4378
		x"58",	--4379
		x"3c",	--4380
		x"f6",	--4381
		x"3d",	--4382
		x"0f",	--4383
		x"b0",	--4384
		x"bc",	--4385
		x"0c",	--4386
		x"0d",	--4387
		x"0e",	--4388
		x"0f",	--4389
		x"b0",	--4390
		x"58",	--4391
		x"3c",	--4392
		x"7c",	--4393
		x"3d",	--4394
		x"93",	--4395
		x"b0",	--4396
		x"08",	--4397
		x"0c",	--4398
		x"0d",	--4399
		x"0e",	--4400
		x"0f",	--4401
		x"b0",	--4402
		x"58",	--4403
		x"3c",	--4404
		x"01",	--4405
		x"3d",	--4406
		x"d0",	--4407
		x"b0",	--4408
		x"bc",	--4409
		x"0c",	--4410
		x"0d",	--4411
		x"0e",	--4412
		x"0f",	--4413
		x"b0",	--4414
		x"58",	--4415
		x"3c",	--4416
		x"61",	--4417
		x"3d",	--4418
		x"b6",	--4419
		x"b0",	--4420
		x"08",	--4421
		x"0c",	--4422
		x"0d",	--4423
		x"0e",	--4424
		x"0f",	--4425
		x"b0",	--4426
		x"58",	--4427
		x"3c",	--4428
		x"ab",	--4429
		x"3d",	--4430
		x"2a",	--4431
		x"b0",	--4432
		x"bc",	--4433
		x"0c",	--4434
		x"0d",	--4435
		x"0e",	--4436
		x"0f",	--4437
		x"b0",	--4438
		x"58",	--4439
		x"81",	--4440
		x"00",	--4441
		x"81",	--4442
		x"02",	--4443
		x"3b",	--4444
		x"99",	--4445
		x"06",	--4446
		x"3b",	--4447
		x"9a",	--4448
		x"2d",	--4449
		x"3a",	--4450
		x"9a",	--4451
		x"2a",	--4452
		x"0c",	--4453
		x"3d",	--4454
		x"00",	--4455
		x"0e",	--4456
		x"0f",	--4457
		x"b0",	--4458
		x"58",	--4459
		x"0a",	--4460
		x"0b",	--4461
		x"2c",	--4462
		x"1d",	--4463
		x"02",	--4464
		x"0e",	--4465
		x"0f",	--4466
		x"b0",	--4467
		x"58",	--4468
		x"08",	--4469
		x"09",	--4470
		x"0c",	--4471
		x"0d",	--4472
		x"0e",	--4473
		x"0f",	--4474
		x"b0",	--4475
		x"58",	--4476
		x"0c",	--4477
		x"0d",	--4478
		x"0e",	--4479
		x"0f",	--4480
		x"b0",	--4481
		x"08",	--4482
		x"0c",	--4483
		x"0d",	--4484
		x"0e",	--4485
		x"0f",	--4486
		x"b0",	--4487
		x"08",	--4488
		x"0c",	--4489
		x"0d",	--4490
		x"0e",	--4491
		x"3f",	--4492
		x"80",	--4493
		x"48",	--4494
		x"3b",	--4495
		x"48",	--4496
		x"05",	--4497
		x"3b",	--4498
		x"49",	--4499
		x"06",	--4500
		x"1a",	--4501
		x"04",	--4502
		x"0a",	--4503
		x"3b",	--4504
		x"00",	--4505
		x"03",	--4506
		x"0a",	--4507
		x"3b",	--4508
		x"90",	--4509
		x"0c",	--4510
		x"0d",	--4511
		x"0e",	--4512
		x"3f",	--4513
		x"80",	--4514
		x"b0",	--4515
		x"08",	--4516
		x"81",	--4517
		x"04",	--4518
		x"81",	--4519
		x"06",	--4520
		x"0c",	--4521
		x"3d",	--4522
		x"00",	--4523
		x"0e",	--4524
		x"0f",	--4525
		x"b0",	--4526
		x"58",	--4527
		x"0c",	--4528
		x"0d",	--4529
		x"b0",	--4530
		x"08",	--4531
		x"0a",	--4532
		x"0b",	--4533
		x"2c",	--4534
		x"1d",	--4535
		x"02",	--4536
		x"0e",	--4537
		x"0f",	--4538
		x"b0",	--4539
		x"58",	--4540
		x"08",	--4541
		x"09",	--4542
		x"0c",	--4543
		x"0d",	--4544
		x"0e",	--4545
		x"0f",	--4546
		x"b0",	--4547
		x"58",	--4548
		x"0c",	--4549
		x"0d",	--4550
		x"0e",	--4551
		x"0f",	--4552
		x"b0",	--4553
		x"08",	--4554
		x"0c",	--4555
		x"0d",	--4556
		x"0e",	--4557
		x"0f",	--4558
		x"b0",	--4559
		x"08",	--4560
		x"0c",	--4561
		x"0d",	--4562
		x"1e",	--4563
		x"04",	--4564
		x"1f",	--4565
		x"06",	--4566
		x"b0",	--4567
		x"08",	--4568
		x"03",	--4569
		x"0e",	--4570
		x"3f",	--4571
		x"80",	--4572
		x"31",	--4573
		x"34",	--4574
		x"35",	--4575
		x"36",	--4576
		x"37",	--4577
		x"38",	--4578
		x"39",	--4579
		x"3a",	--4580
		x"3b",	--4581
		x"30",	--4582
		x"0b",	--4583
		x"0a",	--4584
		x"09",	--4585
		x"08",	--4586
		x"07",	--4587
		x"06",	--4588
		x"05",	--4589
		x"04",	--4590
		x"31",	--4591
		x"de",	--4592
		x"81",	--4593
		x"0c",	--4594
		x"81",	--4595
		x"12",	--4596
		x"81",	--4597
		x"14",	--4598
		x"0a",	--4599
		x"0b",	--4600
		x"3a",	--4601
		x"3b",	--4602
		x"ff",	--4603
		x"3b",	--4604
		x"49",	--4605
		x"06",	--4606
		x"3b",	--4607
		x"4a",	--4608
		x"0f",	--4609
		x"3a",	--4610
		x"d9",	--4611
		x"0c",	--4612
		x"1d",	--4613
		x"0c",	--4614
		x"8d",	--4615
		x"00",	--4616
		x"8d",	--4617
		x"02",	--4618
		x"8d",	--4619
		x"04",	--4620
		x"8d",	--4621
		x"06",	--4622
		x"30",	--4623
		x"9a",	--4624
		x"3b",	--4625
		x"16",	--4626
		x"06",	--4627
		x"3b",	--4628
		x"17",	--4629
		x"b2",	--4630
		x"3a",	--4631
		x"e4",	--4632
		x"af",	--4633
		x"81",	--4634
		x"14",	--4635
		x"58",	--4636
		x"03",	--4637
		x"91",	--4638
		x"12",	--4639
		x"54",	--4640
		x"3c",	--4641
		x"80",	--4642
		x"3d",	--4643
		x"c9",	--4644
		x"b0",	--4645
		x"08",	--4646
		x"08",	--4647
		x"09",	--4648
		x"3a",	--4649
		x"f0",	--4650
		x"3b",	--4651
		x"3a",	--4652
		x"d0",	--4653
		x"03",	--4654
		x"3b",	--4655
		x"c9",	--4656
		x"19",	--4657
		x"3c",	--4658
		x"43",	--4659
		x"3d",	--4660
		x"35",	--4661
		x"0e",	--4662
		x"0f",	--4663
		x"b0",	--4664
		x"08",	--4665
		x"0c",	--4666
		x"0d",	--4667
		x"1f",	--4668
		x"0c",	--4669
		x"8f",	--4670
		x"00",	--4671
		x"8f",	--4672
		x"02",	--4673
		x"0e",	--4674
		x"0f",	--4675
		x"b0",	--4676
		x"08",	--4677
		x"3c",	--4678
		x"43",	--4679
		x"3d",	--4680
		x"35",	--4681
		x"1e",	--4682
		x"3c",	--4683
		x"00",	--4684
		x"3d",	--4685
		x"35",	--4686
		x"b0",	--4687
		x"08",	--4688
		x"0a",	--4689
		x"0b",	--4690
		x"3c",	--4691
		x"08",	--4692
		x"3d",	--4693
		x"85",	--4694
		x"b0",	--4695
		x"08",	--4696
		x"0c",	--4697
		x"0d",	--4698
		x"1e",	--4699
		x"0c",	--4700
		x"8e",	--4701
		x"00",	--4702
		x"8e",	--4703
		x"02",	--4704
		x"0e",	--4705
		x"0f",	--4706
		x"b0",	--4707
		x"08",	--4708
		x"3c",	--4709
		x"08",	--4710
		x"3d",	--4711
		x"85",	--4712
		x"b0",	--4713
		x"08",	--4714
		x"1d",	--4715
		x"0c",	--4716
		x"8d",	--4717
		x"04",	--4718
		x"8d",	--4719
		x"06",	--4720
		x"16",	--4721
		x"07",	--4722
		x"30",	--4723
		x"94",	--4724
		x"3c",	--4725
		x"80",	--4726
		x"3d",	--4727
		x"c9",	--4728
		x"b0",	--4729
		x"bc",	--4730
		x"08",	--4731
		x"09",	--4732
		x"3a",	--4733
		x"f0",	--4734
		x"3b",	--4735
		x"3a",	--4736
		x"d0",	--4737
		x"03",	--4738
		x"3b",	--4739
		x"c9",	--4740
		x"19",	--4741
		x"3c",	--4742
		x"43",	--4743
		x"3d",	--4744
		x"35",	--4745
		x"0e",	--4746
		x"0f",	--4747
		x"b0",	--4748
		x"bc",	--4749
		x"0c",	--4750
		x"0d",	--4751
		x"1e",	--4752
		x"0c",	--4753
		x"8e",	--4754
		x"00",	--4755
		x"8e",	--4756
		x"02",	--4757
		x"0e",	--4758
		x"0f",	--4759
		x"b0",	--4760
		x"08",	--4761
		x"3c",	--4762
		x"43",	--4763
		x"3d",	--4764
		x"35",	--4765
		x"1e",	--4766
		x"3c",	--4767
		x"00",	--4768
		x"3d",	--4769
		x"35",	--4770
		x"b0",	--4771
		x"bc",	--4772
		x"0a",	--4773
		x"0b",	--4774
		x"3c",	--4775
		x"08",	--4776
		x"3d",	--4777
		x"85",	--4778
		x"b0",	--4779
		x"bc",	--4780
		x"0c",	--4781
		x"0d",	--4782
		x"1e",	--4783
		x"0c",	--4784
		x"8e",	--4785
		x"00",	--4786
		x"8e",	--4787
		x"02",	--4788
		x"0e",	--4789
		x"0f",	--4790
		x"b0",	--4791
		x"08",	--4792
		x"3c",	--4793
		x"08",	--4794
		x"3d",	--4795
		x"85",	--4796
		x"b0",	--4797
		x"bc",	--4798
		x"1d",	--4799
		x"0c",	--4800
		x"8d",	--4801
		x"04",	--4802
		x"8d",	--4803
		x"06",	--4804
		x"36",	--4805
		x"37",	--4806
		x"30",	--4807
		x"94",	--4808
		x"3b",	--4809
		x"49",	--4810
		x"0a",	--4811
		x"3b",	--4812
		x"4a",	--4813
		x"02",	--4814
		x"30",	--4815
		x"78",	--4816
		x"3a",	--4817
		x"81",	--4818
		x"02",	--4819
		x"30",	--4820
		x"78",	--4821
		x"08",	--4822
		x"09",	--4823
		x"39",	--4824
		x"ff",	--4825
		x"3c",	--4826
		x"84",	--4827
		x"3d",	--4828
		x"22",	--4829
		x"0e",	--4830
		x"0f",	--4831
		x"b0",	--4832
		x"58",	--4833
		x"0c",	--4834
		x"3d",	--4835
		x"00",	--4836
		x"b0",	--4837
		x"bc",	--4838
		x"b0",	--4839
		x"02",	--4840
		x"06",	--4841
		x"07",	--4842
		x"b0",	--4843
		x"5c",	--4844
		x"81",	--4845
		x"1a",	--4846
		x"81",	--4847
		x"1c",	--4848
		x"3c",	--4849
		x"80",	--4850
		x"3d",	--4851
		x"c9",	--4852
		x"b0",	--4853
		x"58",	--4854
		x"0c",	--4855
		x"0d",	--4856
		x"0e",	--4857
		x"0f",	--4858
		x"b0",	--4859
		x"08",	--4860
		x"04",	--4861
		x"05",	--4862
		x"3c",	--4863
		x"43",	--4864
		x"3d",	--4865
		x"35",	--4866
		x"1e",	--4867
		x"1a",	--4868
		x"1f",	--4869
		x"1c",	--4870
		x"b0",	--4871
		x"58",	--4872
		x"81",	--4873
		x"0e",	--4874
		x"81",	--4875
		x"10",	--4876
		x"07",	--4877
		x"05",	--4878
		x"17",	--4879
		x"19",	--4880
		x"36",	--4881
		x"20",	--4882
		x"16",	--4883
		x"08",	--4884
		x"09",	--4885
		x"38",	--4886
		x"00",	--4887
		x"39",	--4888
		x"0f",	--4889
		x"3f",	--4890
		x"0f",	--4891
		x"0f",	--4892
		x"3f",	--4893
		x"74",	--4894
		x"28",	--4895
		x"03",	--4896
		x"19",	--4897
		x"02",	--4898
		x"06",	--4899
		x"1c",	--4900
		x"0e",	--4901
		x"1d",	--4902
		x"10",	--4903
		x"30",	--4904
		x"00",	--4905
		x"1c",	--4906
		x"0e",	--4907
		x"1d",	--4908
		x"10",	--4909
		x"0e",	--4910
		x"0f",	--4911
		x"b0",	--4912
		x"08",	--4913
		x"08",	--4914
		x"09",	--4915
		x"1e",	--4916
		x"0c",	--4917
		x"8e",	--4918
		x"00",	--4919
		x"8e",	--4920
		x"02",	--4921
		x"81",	--4922
		x"16",	--4923
		x"0d",	--4924
		x"8d",	--4925
		x"8d",	--4926
		x"8d",	--4927
		x"8d",	--4928
		x"81",	--4929
		x"18",	--4930
		x"7d",	--4931
		x"07",	--4932
		x"0c",	--4933
		x"1e",	--4934
		x"16",	--4935
		x"1f",	--4936
		x"18",	--4937
		x"0f",	--4938
		x"0e",	--4939
		x"7d",	--4940
		x"fc",	--4941
		x"81",	--4942
		x"16",	--4943
		x"81",	--4944
		x"18",	--4945
		x"0a",	--4946
		x"0b",	--4947
		x"7f",	--4948
		x"07",	--4949
		x"12",	--4950
		x"0b",	--4951
		x"0a",	--4952
		x"7f",	--4953
		x"fb",	--4954
		x"3a",	--4955
		x"ff",	--4956
		x"0b",	--4957
		x"18",	--4958
		x"16",	--4959
		x"19",	--4960
		x"18",	--4961
		x"08",	--4962
		x"09",	--4963
		x"09",	--4964
		x"a9",	--4965
		x"03",	--4966
		x"38",	--4967
		x"09",	--4968
		x"a5",	--4969
		x"3c",	--4970
		x"00",	--4971
		x"3d",	--4972
		x"35",	--4973
		x"1e",	--4974
		x"1a",	--4975
		x"1f",	--4976
		x"1c",	--4977
		x"b0",	--4978
		x"58",	--4979
		x"08",	--4980
		x"09",	--4981
		x"0c",	--4982
		x"0d",	--4983
		x"0e",	--4984
		x"0f",	--4985
		x"b0",	--4986
		x"08",	--4987
		x"81",	--4988
		x"1e",	--4989
		x"81",	--4990
		x"20",	--4991
		x"0c",	--4992
		x"0d",	--4993
		x"0e",	--4994
		x"0f",	--4995
		x"b0",	--4996
		x"08",	--4997
		x"0c",	--4998
		x"0d",	--4999
		x"b0",	--5000
		x"08",	--5001
		x"08",	--5002
		x"09",	--5003
		x"3c",	--5004
		x"08",	--5005
		x"3d",	--5006
		x"85",	--5007
		x"1e",	--5008
		x"1a",	--5009
		x"1f",	--5010
		x"1c",	--5011
		x"b0",	--5012
		x"58",	--5013
		x"0c",	--5014
		x"0d",	--5015
		x"b0",	--5016
		x"08",	--5017
		x"81",	--5018
		x"0e",	--5019
		x"81",	--5020
		x"10",	--5021
		x"0c",	--5022
		x"0d",	--5023
		x"1e",	--5024
		x"1e",	--5025
		x"1f",	--5026
		x"20",	--5027
		x"b0",	--5028
		x"08",	--5029
		x"0a",	--5030
		x"0b",	--5031
		x"1e",	--5032
		x"0c",	--5033
		x"8e",	--5034
		x"00",	--5035
		x"8e",	--5036
		x"02",	--5037
		x"0a",	--5038
		x"0b",	--5039
		x"7f",	--5040
		x"07",	--5041
		x"12",	--5042
		x"0b",	--5043
		x"0a",	--5044
		x"7f",	--5045
		x"fb",	--5046
		x"3a",	--5047
		x"ff",	--5048
		x"0b",	--5049
		x"1d",	--5050
		x"16",	--5051
		x"1e",	--5052
		x"18",	--5053
		x"0d",	--5054
		x"0e",	--5055
		x"0a",	--5056
		x"0b",	--5057
		x"0b",	--5058
		x"47",	--5059
		x"03",	--5060
		x"3d",	--5061
		x"1a",	--5062
		x"43",	--5063
		x"3c",	--5064
		x"00",	--5065
		x"3d",	--5066
		x"85",	--5067
		x"1e",	--5068
		x"1a",	--5069
		x"1f",	--5070
		x"1c",	--5071
		x"b0",	--5072
		x"58",	--5073
		x"0a",	--5074
		x"0b",	--5075
		x"0c",	--5076
		x"0d",	--5077
		x"1e",	--5078
		x"1e",	--5079
		x"1f",	--5080
		x"20",	--5081
		x"b0",	--5082
		x"08",	--5083
		x"04",	--5084
		x"05",	--5085
		x"0c",	--5086
		x"0d",	--5087
		x"1e",	--5088
		x"1e",	--5089
		x"1f",	--5090
		x"20",	--5091
		x"b0",	--5092
		x"08",	--5093
		x"0c",	--5094
		x"0d",	--5095
		x"b0",	--5096
		x"08",	--5097
		x"0a",	--5098
		x"0b",	--5099
		x"3c",	--5100
		x"32",	--5101
		x"3d",	--5102
		x"8d",	--5103
		x"1e",	--5104
		x"1a",	--5105
		x"1f",	--5106
		x"1c",	--5107
		x"b0",	--5108
		x"58",	--5109
		x"0c",	--5110
		x"0d",	--5111
		x"b0",	--5112
		x"08",	--5113
		x"81",	--5114
		x"0e",	--5115
		x"81",	--5116
		x"10",	--5117
		x"0c",	--5118
		x"0d",	--5119
		x"0e",	--5120
		x"0f",	--5121
		x"b0",	--5122
		x"08",	--5123
		x"1d",	--5124
		x"0c",	--5125
		x"8d",	--5126
		x"00",	--5127
		x"8d",	--5128
		x"02",	--5129
		x"04",	--5130
		x"14",	--5131
		x"1e",	--5132
		x"15",	--5133
		x"20",	--5134
		x"1e",	--5135
		x"0c",	--5136
		x"28",	--5137
		x"19",	--5138
		x"02",	--5139
		x"0c",	--5140
		x"0d",	--5141
		x"0e",	--5142
		x"0f",	--5143
		x"b0",	--5144
		x"08",	--5145
		x"1c",	--5146
		x"0e",	--5147
		x"1d",	--5148
		x"10",	--5149
		x"b0",	--5150
		x"08",	--5151
		x"0a",	--5152
		x"0b",	--5153
		x"1f",	--5154
		x"0c",	--5155
		x"8f",	--5156
		x"04",	--5157
		x"8f",	--5158
		x"06",	--5159
		x"81",	--5160
		x"14",	--5161
		x"9f",	--5162
		x"0d",	--5163
		x"0e",	--5164
		x"3e",	--5165
		x"00",	--5166
		x"8f",	--5167
		x"00",	--5168
		x"8f",	--5169
		x"02",	--5170
		x"0d",	--5171
		x"0e",	--5172
		x"3e",	--5173
		x"00",	--5174
		x"8f",	--5175
		x"04",	--5176
		x"8f",	--5177
		x"06",	--5178
		x"8a",	--5179
		x"3b",	--5180
		x"80",	--5181
		x"11",	--5182
		x"0c",	--5183
		x"0d",	--5184
		x"b0",	--5185
		x"08",	--5186
		x"1d",	--5187
		x"0c",	--5188
		x"8d",	--5189
		x"04",	--5190
		x"8d",	--5191
		x"06",	--5192
		x"8d",	--5193
		x"00",	--5194
		x"8d",	--5195
		x"02",	--5196
		x"06",	--5197
		x"07",	--5198
		x"7a",	--5199
		x"0c",	--5200
		x"0d",	--5201
		x"8d",	--5202
		x"8d",	--5203
		x"8d",	--5204
		x"8d",	--5205
		x"7f",	--5206
		x"07",	--5207
		x"0d",	--5208
		x"0c",	--5209
		x"7f",	--5210
		x"fc",	--5211
		x"09",	--5212
		x"39",	--5213
		x"7a",	--5214
		x"0c",	--5215
		x"0d",	--5216
		x"0d",	--5217
		x"7f",	--5218
		x"07",	--5219
		x"0c",	--5220
		x"0d",	--5221
		x"7f",	--5222
		x"fc",	--5223
		x"0a",	--5224
		x"0b",	--5225
		x"0e",	--5226
		x"0f",	--5227
		x"b0",	--5228
		x"02",	--5229
		x"b0",	--5230
		x"5c",	--5231
		x"0c",	--5232
		x"0d",	--5233
		x"81",	--5234
		x"00",	--5235
		x"81",	--5236
		x"02",	--5237
		x"0e",	--5238
		x"0f",	--5239
		x"b0",	--5240
		x"08",	--5241
		x"0c",	--5242
		x"3d",	--5243
		x"80",	--5244
		x"b0",	--5245
		x"58",	--5246
		x"0a",	--5247
		x"0b",	--5248
		x"b0",	--5249
		x"02",	--5250
		x"b0",	--5251
		x"5c",	--5252
		x"0c",	--5253
		x"0d",	--5254
		x"81",	--5255
		x"04",	--5256
		x"81",	--5257
		x"06",	--5258
		x"0e",	--5259
		x"0f",	--5260
		x"b0",	--5261
		x"08",	--5262
		x"0c",	--5263
		x"3d",	--5264
		x"80",	--5265
		x"b0",	--5266
		x"58",	--5267
		x"81",	--5268
		x"08",	--5269
		x"81",	--5270
		x"0a",	--5271
		x"08",	--5272
		x"38",	--5273
		x"3a",	--5274
		x"03",	--5275
		x"01",	--5276
		x"3a",	--5277
		x"28",	--5278
		x"0c",	--5279
		x"0d",	--5280
		x"1e",	--5281
		x"04",	--5282
		x"1f",	--5283
		x"06",	--5284
		x"b0",	--5285
		x"cc",	--5286
		x"0f",	--5287
		x"f4",	--5288
		x"30",	--5289
		x"f4",	--5290
		x"23",	--5291
		x"0c",	--5292
		x"0d",	--5293
		x"1e",	--5294
		x"10",	--5295
		x"0f",	--5296
		x"2f",	--5297
		x"b0",	--5298
		x"ae",	--5299
		x"21",	--5300
		x"06",	--5301
		x"8f",	--5302
		x"8f",	--5303
		x"8f",	--5304
		x"8f",	--5305
		x"07",	--5306
		x"81",	--5307
		x"14",	--5308
		x"0c",	--5309
		x"1e",	--5310
		x"0c",	--5311
		x"be",	--5312
		x"00",	--5313
		x"02",	--5314
		x"be",	--5315
		x"00",	--5316
		x"06",	--5317
		x"36",	--5318
		x"37",	--5319
		x"16",	--5320
		x"07",	--5321
		x"0e",	--5322
		x"0f",	--5323
		x"31",	--5324
		x"22",	--5325
		x"34",	--5326
		x"35",	--5327
		x"36",	--5328
		x"37",	--5329
		x"38",	--5330
		x"39",	--5331
		x"3a",	--5332
		x"3b",	--5333
		x"30",	--5334
		x"0b",	--5335
		x"0a",	--5336
		x"09",	--5337
		x"08",	--5338
		x"07",	--5339
		x"06",	--5340
		x"05",	--5341
		x"04",	--5342
		x"31",	--5343
		x"8c",	--5344
		x"81",	--5345
		x"66",	--5346
		x"81",	--5347
		x"60",	--5348
		x"81",	--5349
		x"48",	--5350
		x"1a",	--5351
		x"86",	--5352
		x"0a",	--5353
		x"81",	--5354
		x"4c",	--5355
		x"81",	--5356
		x"4e",	--5357
		x"91",	--5358
		x"0c",	--5359
		x"4c",	--5360
		x"1a",	--5361
		x"4c",	--5362
		x"8a",	--5363
		x"8a",	--5364
		x"8a",	--5365
		x"8a",	--5366
		x"81",	--5367
		x"4e",	--5368
		x"0a",	--5369
		x"3a",	--5370
		x"81",	--5371
		x"50",	--5372
		x"8a",	--5373
		x"8a",	--5374
		x"8a",	--5375
		x"8a",	--5376
		x"81",	--5377
		x"52",	--5378
		x"0a",	--5379
		x"3a",	--5380
		x"fd",	--5381
		x"0a",	--5382
		x"02",	--5383
		x"3a",	--5384
		x"07",	--5385
		x"0a",	--5386
		x"0a",	--5387
		x"0a",	--5388
		x"08",	--5389
		x"88",	--5390
		x"88",	--5391
		x"88",	--5392
		x"88",	--5393
		x"81",	--5394
		x"54",	--5395
		x"81",	--5396
		x"56",	--5397
		x"04",	--5398
		x"81",	--5399
		x"54",	--5400
		x"81",	--5401
		x"56",	--5402
		x"08",	--5403
		x"8d",	--5404
		x"8d",	--5405
		x"8d",	--5406
		x"8d",	--5407
		x"09",	--5408
		x"1a",	--5409
		x"54",	--5410
		x"1b",	--5411
		x"56",	--5412
		x"3a",	--5413
		x"3b",	--5414
		x"0a",	--5415
		x"0b",	--5416
		x"0a",	--5417
		x"0b",	--5418
		x"0a",	--5419
		x"0b",	--5420
		x"0d",	--5421
		x"0e",	--5422
		x"0d",	--5423
		x"0e",	--5424
		x"81",	--5425
		x"44",	--5426
		x"81",	--5427
		x"46",	--5428
		x"18",	--5429
		x"54",	--5430
		x"19",	--5431
		x"56",	--5432
		x"18",	--5433
		x"50",	--5434
		x"19",	--5435
		x"52",	--5436
		x"81",	--5437
		x"40",	--5438
		x"81",	--5439
		x"42",	--5440
		x"14",	--5441
		x"50",	--5442
		x"15",	--5443
		x"52",	--5444
		x"14",	--5445
		x"4c",	--5446
		x"15",	--5447
		x"4e",	--5448
		x"09",	--5449
		x"06",	--5450
		x"07",	--5451
		x"22",	--5452
		x"1e",	--5453
		x"40",	--5454
		x"1f",	--5455
		x"42",	--5456
		x"0e",	--5457
		x"0f",	--5458
		x"0f",	--5459
		x"0d",	--5460
		x"1f",	--5461
		x"40",	--5462
		x"0f",	--5463
		x"0f",	--5464
		x"1f",	--5465
		x"88",	--5466
		x"0f",	--5467
		x"2e",	--5468
		x"1f",	--5469
		x"02",	--5470
		x"b0",	--5471
		x"5c",	--5472
		x"02",	--5473
		x"0e",	--5474
		x"0f",	--5475
		x"3d",	--5476
		x"a0",	--5477
		x"0d",	--5478
		x"0d",	--5479
		x"8d",	--5480
		x"00",	--5481
		x"8d",	--5482
		x"02",	--5483
		x"16",	--5484
		x"07",	--5485
		x"29",	--5486
		x"05",	--5487
		x"04",	--5488
		x"07",	--5489
		x"da",	--5490
		x"04",	--5491
		x"d8",	--5492
		x"81",	--5493
		x"40",	--5494
		x"81",	--5495
		x"42",	--5496
		x"04",	--5497
		x"2d",	--5498
		x"1f",	--5499
		x"48",	--5500
		x"3f",	--5501
		x"0f",	--5502
		x"0f",	--5503
		x"3f",	--5504
		x"a0",	--5505
		x"0f",	--5506
		x"0f",	--5507
		x"2c",	--5508
		x"1d",	--5509
		x"02",	--5510
		x"3e",	--5511
		x"3f",	--5512
		x"b0",	--5513
		x"58",	--5514
		x"0c",	--5515
		x"0d",	--5516
		x"0e",	--5517
		x"0f",	--5518
		x"b0",	--5519
		x"bc",	--5520
		x"0a",	--5521
		x"0b",	--5522
		x"18",	--5523
		x"09",	--5524
		x"25",	--5525
		x"81",	--5526
		x"52",	--5527
		x"06",	--5528
		x"19",	--5529
		x"52",	--5530
		x"df",	--5531
		x"81",	--5532
		x"50",	--5533
		x"dc",	--5534
		x"84",	--5535
		x"00",	--5536
		x"84",	--5537
		x"02",	--5538
		x"91",	--5539
		x"40",	--5540
		x"81",	--5541
		x"42",	--5542
		x"24",	--5543
		x"91",	--5544
		x"42",	--5545
		x"4e",	--5546
		x"08",	--5547
		x"91",	--5548
		x"4e",	--5549
		x"42",	--5550
		x"15",	--5551
		x"91",	--5552
		x"40",	--5553
		x"4c",	--5554
		x"11",	--5555
		x"91",	--5556
		x"4c",	--5557
		x"40",	--5558
		x"91",	--5559
		x"4e",	--5560
		x"42",	--5561
		x"19",	--5562
		x"4c",	--5563
		x"1a",	--5564
		x"4e",	--5565
		x"39",	--5566
		x"3a",	--5567
		x"81",	--5568
		x"70",	--5569
		x"81",	--5570
		x"72",	--5571
		x"08",	--5572
		x"17",	--5573
		x"66",	--5574
		x"05",	--5575
		x"0a",	--5576
		x"0b",	--5577
		x"08",	--5578
		x"09",	--5579
		x"c9",	--5580
		x"1f",	--5581
		x"40",	--5582
		x"0f",	--5583
		x"0f",	--5584
		x"0f",	--5585
		x"28",	--5586
		x"19",	--5587
		x"02",	--5588
		x"0a",	--5589
		x"3a",	--5590
		x"f0",	--5591
		x"81",	--5592
		x"62",	--5593
		x"16",	--5594
		x"40",	--5595
		x"17",	--5596
		x"42",	--5597
		x"81",	--5598
		x"48",	--5599
		x"04",	--5600
		x"05",	--5601
		x"34",	--5602
		x"35",	--5603
		x"81",	--5604
		x"58",	--5605
		x"81",	--5606
		x"5a",	--5607
		x"05",	--5608
		x"32",	--5609
		x"0c",	--5610
		x"3d",	--5611
		x"80",	--5612
		x"0e",	--5613
		x"0f",	--5614
		x"b0",	--5615
		x"58",	--5616
		x"b0",	--5617
		x"02",	--5618
		x"b0",	--5619
		x"5c",	--5620
		x"0a",	--5621
		x"0b",	--5622
		x"0c",	--5623
		x"3d",	--5624
		x"80",	--5625
		x"b0",	--5626
		x"58",	--5627
		x"0c",	--5628
		x"0d",	--5629
		x"0e",	--5630
		x"0f",	--5631
		x"b0",	--5632
		x"08",	--5633
		x"b0",	--5634
		x"02",	--5635
		x"85",	--5636
		x"00",	--5637
		x"85",	--5638
		x"02",	--5639
		x"1f",	--5640
		x"58",	--5641
		x"0f",	--5642
		x"0f",	--5643
		x"0f",	--5644
		x"1f",	--5645
		x"48",	--5646
		x"1c",	--5647
		x"04",	--5648
		x"1d",	--5649
		x"06",	--5650
		x"0e",	--5651
		x"0f",	--5652
		x"b0",	--5653
		x"bc",	--5654
		x"08",	--5655
		x"09",	--5656
		x"36",	--5657
		x"37",	--5658
		x"25",	--5659
		x"a1",	--5660
		x"48",	--5661
		x"07",	--5662
		x"04",	--5663
		x"17",	--5664
		x"c8",	--5665
		x"16",	--5666
		x"c6",	--5667
		x"91",	--5668
		x"44",	--5669
		x"5c",	--5670
		x"1d",	--5671
		x"44",	--5672
		x"0e",	--5673
		x"0f",	--5674
		x"b0",	--5675
		x"48",	--5676
		x"0a",	--5677
		x"0b",	--5678
		x"0c",	--5679
		x"3d",	--5680
		x"00",	--5681
		x"b0",	--5682
		x"58",	--5683
		x"b0",	--5684
		x"cc",	--5685
		x"0c",	--5686
		x"3d",	--5687
		x"00",	--5688
		x"b0",	--5689
		x"58",	--5690
		x"0c",	--5691
		x"0d",	--5692
		x"0e",	--5693
		x"0f",	--5694
		x"b0",	--5695
		x"08",	--5696
		x"0a",	--5697
		x"0b",	--5698
		x"b0",	--5699
		x"02",	--5700
		x"81",	--5701
		x"58",	--5702
		x"81",	--5703
		x"5a",	--5704
		x"b0",	--5705
		x"5c",	--5706
		x"0c",	--5707
		x"0d",	--5708
		x"0e",	--5709
		x"0f",	--5710
		x"b0",	--5711
		x"08",	--5712
		x"81",	--5713
		x"48",	--5714
		x"81",	--5715
		x"4a",	--5716
		x"81",	--5717
		x"46",	--5718
		x"46",	--5719
		x"03",	--5720
		x"91",	--5721
		x"44",	--5722
		x"42",	--5723
		x"1c",	--5724
		x"40",	--5725
		x"1d",	--5726
		x"42",	--5727
		x"3c",	--5728
		x"3d",	--5729
		x"0b",	--5730
		x"0b",	--5731
		x"0b",	--5732
		x"0b",	--5733
		x"16",	--5734
		x"f0",	--5735
		x"17",	--5736
		x"f2",	--5737
		x"1e",	--5738
		x"44",	--5739
		x"39",	--5740
		x"09",	--5741
		x"0a",	--5742
		x"0b",	--5743
		x"48",	--5744
		x"78",	--5745
		x"1f",	--5746
		x"48",	--5747
		x"04",	--5748
		x"0b",	--5749
		x"0a",	--5750
		x"78",	--5751
		x"fa",	--5752
		x"81",	--5753
		x"58",	--5754
		x"81",	--5755
		x"5a",	--5756
		x"79",	--5757
		x"1f",	--5758
		x"49",	--5759
		x"04",	--5760
		x"0a",	--5761
		x"0b",	--5762
		x"79",	--5763
		x"fa",	--5764
		x"08",	--5765
		x"09",	--5766
		x"08",	--5767
		x"09",	--5768
		x"0f",	--5769
		x"0f",	--5770
		x"0f",	--5771
		x"0f",	--5772
		x"8f",	--5773
		x"f0",	--5774
		x"8f",	--5775
		x"f2",	--5776
		x"06",	--5777
		x"07",	--5778
		x"3f",	--5779
		x"07",	--5780
		x"4f",	--5781
		x"7f",	--5782
		x"1f",	--5783
		x"4f",	--5784
		x"28",	--5785
		x"07",	--5786
		x"06",	--5787
		x"7f",	--5788
		x"fa",	--5789
		x"81",	--5790
		x"44",	--5791
		x"13",	--5792
		x"81",	--5793
		x"46",	--5794
		x"10",	--5795
		x"1f",	--5796
		x"40",	--5797
		x"3f",	--5798
		x"0f",	--5799
		x"0f",	--5800
		x"0f",	--5801
		x"16",	--5802
		x"f0",	--5803
		x"17",	--5804
		x"f2",	--5805
		x"86",	--5806
		x"87",	--5807
		x"46",	--5808
		x"06",	--5809
		x"87",	--5810
		x"0e",	--5811
		x"0c",	--5812
		x"3d",	--5813
		x"00",	--5814
		x"1e",	--5815
		x"48",	--5816
		x"1f",	--5817
		x"4a",	--5818
		x"b0",	--5819
		x"6c",	--5820
		x"0f",	--5821
		x"09",	--5822
		x"06",	--5823
		x"07",	--5824
		x"94",	--5825
		x"07",	--5826
		x"92",	--5827
		x"05",	--5828
		x"16",	--5829
		x"8f",	--5830
		x"02",	--5831
		x"26",	--5832
		x"07",	--5833
		x"91",	--5834
		x"58",	--5835
		x"81",	--5836
		x"5a",	--5837
		x"04",	--5838
		x"05",	--5839
		x"08",	--5840
		x"09",	--5841
		x"1b",	--5842
		x"62",	--5843
		x"27",	--5844
		x"2c",	--5845
		x"1d",	--5846
		x"02",	--5847
		x"08",	--5848
		x"12",	--5849
		x"09",	--5850
		x"10",	--5851
		x"0c",	--5852
		x"02",	--5853
		x"0d",	--5854
		x"19",	--5855
		x"3e",	--5856
		x"00",	--5857
		x"0f",	--5858
		x"09",	--5859
		x"0a",	--5860
		x"09",	--5861
		x"0a",	--5862
		x"8b",	--5863
		x"00",	--5864
		x"8b",	--5865
		x"02",	--5866
		x"0b",	--5867
		x"3e",	--5868
		x"ff",	--5869
		x"0f",	--5870
		x"08",	--5871
		x"09",	--5872
		x"08",	--5873
		x"09",	--5874
		x"8b",	--5875
		x"00",	--5876
		x"8b",	--5877
		x"02",	--5878
		x"18",	--5879
		x"09",	--5880
		x"14",	--5881
		x"05",	--5882
		x"2b",	--5883
		x"15",	--5884
		x"42",	--5885
		x"d6",	--5886
		x"03",	--5887
		x"14",	--5888
		x"40",	--5889
		x"d2",	--5890
		x"81",	--5891
		x"46",	--5892
		x"28",	--5893
		x"03",	--5894
		x"91",	--5895
		x"44",	--5896
		x"24",	--5897
		x"91",	--5898
		x"44",	--5899
		x"03",	--5900
		x"81",	--5901
		x"46",	--5902
		x"07",	--5903
		x"a1",	--5904
		x"44",	--5905
		x"1b",	--5906
		x"81",	--5907
		x"46",	--5908
		x"0d",	--5909
		x"17",	--5910
		x"1f",	--5911
		x"40",	--5912
		x"3f",	--5913
		x"0f",	--5914
		x"0f",	--5915
		x"0f",	--5916
		x"bf",	--5917
		x"7f",	--5918
		x"f0",	--5919
		x"8f",	--5920
		x"f2",	--5921
		x"0b",	--5922
		x"1f",	--5923
		x"40",	--5924
		x"3f",	--5925
		x"0f",	--5926
		x"0f",	--5927
		x"0f",	--5928
		x"bf",	--5929
		x"3f",	--5930
		x"f0",	--5931
		x"8f",	--5932
		x"f2",	--5933
		x"26",	--5934
		x"26",	--5935
		x"07",	--5936
		x"24",	--5937
		x"1c",	--5938
		x"48",	--5939
		x"1d",	--5940
		x"4a",	--5941
		x"0e",	--5942
		x"3f",	--5943
		x"80",	--5944
		x"b0",	--5945
		x"08",	--5946
		x"81",	--5947
		x"48",	--5948
		x"81",	--5949
		x"4a",	--5950
		x"08",	--5951
		x"02",	--5952
		x"09",	--5953
		x"13",	--5954
		x"1d",	--5955
		x"5c",	--5956
		x"0e",	--5957
		x"3f",	--5958
		x"80",	--5959
		x"b0",	--5960
		x"48",	--5961
		x"0c",	--5962
		x"0d",	--5963
		x"1e",	--5964
		x"48",	--5965
		x"1f",	--5966
		x"4a",	--5967
		x"b0",	--5968
		x"08",	--5969
		x"81",	--5970
		x"48",	--5971
		x"81",	--5972
		x"4a",	--5973
		x"0c",	--5974
		x"0d",	--5975
		x"1e",	--5976
		x"48",	--5977
		x"1f",	--5978
		x"4a",	--5979
		x"b0",	--5980
		x"cc",	--5981
		x"0f",	--5982
		x"d7",	--5983
		x"1a",	--5984
		x"40",	--5985
		x"1b",	--5986
		x"42",	--5987
		x"3a",	--5988
		x"3b",	--5989
		x"1c",	--5990
		x"40",	--5991
		x"1d",	--5992
		x"42",	--5993
		x"09",	--5994
		x"81",	--5995
		x"5c",	--5996
		x"81",	--5997
		x"5e",	--5998
		x"0e",	--5999
		x"0f",	--6000
		x"0f",	--6001
		x"0f",	--6002
		x"3e",	--6003
		x"f0",	--6004
		x"0e",	--6005
		x"0f",	--6006
		x"0f",	--6007
		x"91",	--6008
		x"04",	--6009
		x"5c",	--6010
		x"91",	--6011
		x"06",	--6012
		x"5e",	--6013
		x"3c",	--6014
		x"3d",	--6015
		x"29",	--6016
		x"1d",	--6017
		x"4e",	--6018
		x"06",	--6019
		x"81",	--6020
		x"4e",	--6021
		x"e9",	--6022
		x"1c",	--6023
		x"4c",	--6024
		x"e6",	--6025
		x"81",	--6026
		x"5c",	--6027
		x"c3",	--6028
		x"81",	--6029
		x"5e",	--6030
		x"06",	--6031
		x"bf",	--6032
		x"91",	--6033
		x"62",	--6034
		x"81",	--6035
		x"64",	--6036
		x"05",	--6037
		x"0e",	--6038
		x"91",	--6039
		x"62",	--6040
		x"81",	--6041
		x"64",	--6042
		x"2e",	--6043
		x"1f",	--6044
		x"70",	--6045
		x"0f",	--6046
		x"0f",	--6047
		x"38",	--6048
		x"f0",	--6049
		x"08",	--6050
		x"0f",	--6051
		x"0f",	--6052
		x"8f",	--6053
		x"04",	--6054
		x"03",	--6055
		x"8f",	--6056
		x"06",	--6057
		x"e6",	--6058
		x"19",	--6059
		x"40",	--6060
		x"1a",	--6061
		x"42",	--6062
		x"19",	--6063
		x"0a",	--6064
		x"81",	--6065
		x"48",	--6066
		x"81",	--6067
		x"4a",	--6068
		x"81",	--6069
		x"58",	--6070
		x"04",	--6071
		x"81",	--6072
		x"68",	--6073
		x"1d",	--6074
		x"50",	--6075
		x"1e",	--6076
		x"52",	--6077
		x"0d",	--6078
		x"0e",	--6079
		x"81",	--6080
		x"6a",	--6081
		x"81",	--6082
		x"6c",	--6083
		x"08",	--6084
		x"18",	--6085
		x"54",	--6086
		x"81",	--6087
		x"6e",	--6088
		x"06",	--6089
		x"55",	--6090
		x"a1",	--6091
		x"58",	--6092
		x"1f",	--6093
		x"6a",	--6094
		x"0f",	--6095
		x"0f",	--6096
		x"04",	--6097
		x"34",	--6098
		x"a0",	--6099
		x"04",	--6100
		x"1b",	--6101
		x"58",	--6102
		x"0b",	--6103
		x"1f",	--6104
		x"6e",	--6105
		x"0f",	--6106
		x"0f",	--6107
		x"1f",	--6108
		x"88",	--6109
		x"0f",	--6110
		x"2e",	--6111
		x"1f",	--6112
		x"02",	--6113
		x"b0",	--6114
		x"5c",	--6115
		x"8b",	--6116
		x"fc",	--6117
		x"8b",	--6118
		x"fe",	--6119
		x"17",	--6120
		x"66",	--6121
		x"1a",	--6122
		x"5c",	--6123
		x"1b",	--6124
		x"5e",	--6125
		x"05",	--6126
		x"08",	--6127
		x"09",	--6128
		x"04",	--6129
		x"14",	--6130
		x"0f",	--6131
		x"0f",	--6132
		x"2c",	--6133
		x"1d",	--6134
		x"02",	--6135
		x"3e",	--6136
		x"3f",	--6137
		x"b0",	--6138
		x"58",	--6139
		x"0c",	--6140
		x"0d",	--6141
		x"0e",	--6142
		x"0f",	--6143
		x"b0",	--6144
		x"bc",	--6145
		x"08",	--6146
		x"09",	--6147
		x"1a",	--6148
		x"0b",	--6149
		x"25",	--6150
		x"81",	--6151
		x"52",	--6152
		x"06",	--6153
		x"1b",	--6154
		x"52",	--6155
		x"e6",	--6156
		x"81",	--6157
		x"50",	--6158
		x"e3",	--6159
		x"1f",	--6160
		x"68",	--6161
		x"0f",	--6162
		x"0f",	--6163
		x"0f",	--6164
		x"1f",	--6165
		x"58",	--6166
		x"8f",	--6167
		x"fc",	--6168
		x"8f",	--6169
		x"fe",	--6170
		x"91",	--6171
		x"48",	--6172
		x"81",	--6173
		x"4a",	--6174
		x"26",	--6175
		x"1e",	--6176
		x"40",	--6177
		x"1f",	--6178
		x"42",	--6179
		x"1e",	--6180
		x"62",	--6181
		x"1f",	--6182
		x"64",	--6183
		x"1f",	--6184
		x"4a",	--6185
		x"06",	--6186
		x"81",	--6187
		x"4a",	--6188
		x"9d",	--6189
		x"1e",	--6190
		x"48",	--6191
		x"9a",	--6192
		x"81",	--6193
		x"40",	--6194
		x"81",	--6195
		x"42",	--6196
		x"30",	--6197
		x"9a",	--6198
		x"81",	--6199
		x"50",	--6200
		x"81",	--6201
		x"52",	--6202
		x"17",	--6203
		x"5c",	--6204
		x"37",	--6205
		x"0d",	--6206
		x"1d",	--6207
		x"1e",	--6208
		x"48",	--6209
		x"1f",	--6210
		x"4a",	--6211
		x"b0",	--6212
		x"48",	--6213
		x"06",	--6214
		x"07",	--6215
		x"0c",	--6216
		x"3d",	--6217
		x"80",	--6218
		x"b0",	--6219
		x"6c",	--6220
		x"0f",	--6221
		x"2d",	--6222
		x"6b",	--6223
		x"81",	--6224
		x"50",	--6225
		x"81",	--6226
		x"52",	--6227
		x"16",	--6228
		x"40",	--6229
		x"17",	--6230
		x"42",	--6231
		x"36",	--6232
		x"37",	--6233
		x"b1",	--6234
		x"44",	--6235
		x"81",	--6236
		x"46",	--6237
		x"81",	--6238
		x"40",	--6239
		x"81",	--6240
		x"42",	--6241
		x"0d",	--6242
		x"08",	--6243
		x"b1",	--6244
		x"40",	--6245
		x"b1",	--6246
		x"42",	--6247
		x"b1",	--6248
		x"44",	--6249
		x"81",	--6250
		x"46",	--6251
		x"2d",	--6252
		x"0f",	--6253
		x"0f",	--6254
		x"0f",	--6255
		x"39",	--6256
		x"f0",	--6257
		x"09",	--6258
		x"0f",	--6259
		x"0f",	--6260
		x"8f",	--6261
		x"04",	--6262
		x"53",	--6263
		x"8f",	--6264
		x"06",	--6265
		x"e9",	--6266
		x"4f",	--6267
		x"0c",	--6268
		x"3d",	--6269
		x"80",	--6270
		x"0e",	--6271
		x"0f",	--6272
		x"b0",	--6273
		x"58",	--6274
		x"b0",	--6275
		x"02",	--6276
		x"b0",	--6277
		x"5c",	--6278
		x"04",	--6279
		x"05",	--6280
		x"1c",	--6281
		x"40",	--6282
		x"0c",	--6283
		x"0c",	--6284
		x"0b",	--6285
		x"0b",	--6286
		x"3b",	--6287
		x"f0",	--6288
		x"0c",	--6289
		x"3d",	--6290
		x"80",	--6291
		x"b0",	--6292
		x"58",	--6293
		x"0c",	--6294
		x"0d",	--6295
		x"0e",	--6296
		x"0f",	--6297
		x"b0",	--6298
		x"08",	--6299
		x"b0",	--6300
		x"02",	--6301
		x"8b",	--6302
		x"00",	--6303
		x"8b",	--6304
		x"02",	--6305
		x"91",	--6306
		x"40",	--6307
		x"81",	--6308
		x"42",	--6309
		x"b1",	--6310
		x"44",	--6311
		x"81",	--6312
		x"46",	--6313
		x"1c",	--6314
		x"40",	--6315
		x"0c",	--6316
		x"0c",	--6317
		x"07",	--6318
		x"07",	--6319
		x"37",	--6320
		x"f0",	--6321
		x"0e",	--6322
		x"0f",	--6323
		x"b0",	--6324
		x"02",	--6325
		x"87",	--6326
		x"00",	--6327
		x"87",	--6328
		x"02",	--6329
		x"10",	--6330
		x"1c",	--6331
		x"40",	--6332
		x"0c",	--6333
		x"0c",	--6334
		x"05",	--6335
		x"05",	--6336
		x"35",	--6337
		x"f0",	--6338
		x"0e",	--6339
		x"0f",	--6340
		x"b0",	--6341
		x"02",	--6342
		x"85",	--6343
		x"00",	--6344
		x"85",	--6345
		x"02",	--6346
		x"1d",	--6347
		x"44",	--6348
		x"0e",	--6349
		x"3f",	--6350
		x"80",	--6351
		x"b0",	--6352
		x"48",	--6353
		x"06",	--6354
		x"07",	--6355
		x"14",	--6356
		x"40",	--6357
		x"15",	--6358
		x"42",	--6359
		x"0b",	--6360
		x"05",	--6361
		x"28",	--6362
		x"1f",	--6363
		x"40",	--6364
		x"0f",	--6365
		x"0f",	--6366
		x"0a",	--6367
		x"0a",	--6368
		x"0a",	--6369
		x"3d",	--6370
		x"f0",	--6371
		x"0d",	--6372
		x"0f",	--6373
		x"0f",	--6374
		x"2e",	--6375
		x"1f",	--6376
		x"02",	--6377
		x"b0",	--6378
		x"5c",	--6379
		x"0c",	--6380
		x"0d",	--6381
		x"0e",	--6382
		x"0f",	--6383
		x"b0",	--6384
		x"58",	--6385
		x"8a",	--6386
		x"00",	--6387
		x"8a",	--6388
		x"02",	--6389
		x"0c",	--6390
		x"3d",	--6391
		x"80",	--6392
		x"0e",	--6393
		x"0f",	--6394
		x"b0",	--6395
		x"58",	--6396
		x"06",	--6397
		x"07",	--6398
		x"34",	--6399
		x"35",	--6400
		x"2b",	--6401
		x"d6",	--6402
		x"91",	--6403
		x"40",	--6404
		x"44",	--6405
		x"91",	--6406
		x"42",	--6407
		x"46",	--6408
		x"04",	--6409
		x"05",	--6410
		x"07",	--6411
		x"37",	--6412
		x"1f",	--6413
		x"40",	--6414
		x"0f",	--6415
		x"0f",	--6416
		x"0f",	--6417
		x"0f",	--6418
		x"0f",	--6419
		x"2c",	--6420
		x"1d",	--6421
		x"02",	--6422
		x"1e",	--6423
		x"12",	--6424
		x"1f",	--6425
		x"14",	--6426
		x"b0",	--6427
		x"58",	--6428
		x"0c",	--6429
		x"0d",	--6430
		x"0e",	--6431
		x"0f",	--6432
		x"b0",	--6433
		x"bc",	--6434
		x"08",	--6435
		x"09",	--6436
		x"1a",	--6437
		x"0b",	--6438
		x"26",	--6439
		x"81",	--6440
		x"4e",	--6441
		x"0a",	--6442
		x"03",	--6443
		x"81",	--6444
		x"4c",	--6445
		x"06",	--6446
		x"05",	--6447
		x"04",	--6448
		x"0b",	--6449
		x"da",	--6450
		x"04",	--6451
		x"d8",	--6452
		x"3f",	--6453
		x"50",	--6454
		x"0f",	--6455
		x"0f",	--6456
		x"8f",	--6457
		x"00",	--6458
		x"8f",	--6459
		x"02",	--6460
		x"b1",	--6461
		x"44",	--6462
		x"b1",	--6463
		x"46",	--6464
		x"27",	--6465
		x"14",	--6466
		x"05",	--6467
		x"81",	--6468
		x"46",	--6469
		x"06",	--6470
		x"06",	--6471
		x"08",	--6472
		x"09",	--6473
		x"0a",	--6474
		x"0b",	--6475
		x"db",	--6476
		x"b1",	--6477
		x"03",	--6478
		x"86",	--6479
		x"08",	--6480
		x"91",	--6481
		x"86",	--6482
		x"3b",	--6483
		x"81",	--6484
		x"86",	--6485
		x"09",	--6486
		x"30",	--6487
		x"02",	--6488
		x"b1",	--6489
		x"03",	--6490
		x"86",	--6491
		x"02",	--6492
		x"30",	--6493
		x"02",	--6494
		x"cf",	--6495
		x"16",	--6496
		x"40",	--6497
		x"17",	--6498
		x"42",	--6499
		x"05",	--6500
		x"0a",	--6501
		x"0b",	--6502
		x"07",	--6503
		x"16",	--6504
		x"1f",	--6505
		x"40",	--6506
		x"0f",	--6507
		x"0f",	--6508
		x"3e",	--6509
		x"50",	--6510
		x"0e",	--6511
		x"0f",	--6512
		x"0f",	--6513
		x"2c",	--6514
		x"1d",	--6515
		x"02",	--6516
		x"0e",	--6517
		x"0f",	--6518
		x"b0",	--6519
		x"bc",	--6520
		x"0a",	--6521
		x"0b",	--6522
		x"36",	--6523
		x"37",	--6524
		x"25",	--6525
		x"e8",	--6526
		x"81",	--6527
		x"50",	--6528
		x"03",	--6529
		x"81",	--6530
		x"52",	--6531
		x"02",	--6532
		x"3b",	--6533
		x"00",	--6534
		x"18",	--6535
		x"60",	--6536
		x"88",	--6537
		x"00",	--6538
		x"88",	--6539
		x"02",	--6540
		x"30",	--6541
		x"02",	--6542
		x"16",	--6543
		x"40",	--6544
		x"17",	--6545
		x"42",	--6546
		x"05",	--6547
		x"0a",	--6548
		x"0b",	--6549
		x"07",	--6550
		x"16",	--6551
		x"1f",	--6552
		x"40",	--6553
		x"0f",	--6554
		x"0f",	--6555
		x"39",	--6556
		x"50",	--6557
		x"09",	--6558
		x"0f",	--6559
		x"0f",	--6560
		x"2c",	--6561
		x"1d",	--6562
		x"02",	--6563
		x"0e",	--6564
		x"0f",	--6565
		x"b0",	--6566
		x"bc",	--6567
		x"0a",	--6568
		x"0b",	--6569
		x"36",	--6570
		x"37",	--6571
		x"25",	--6572
		x"e8",	--6573
		x"0c",	--6574
		x"0d",	--6575
		x"81",	--6576
		x"50",	--6577
		x"03",	--6578
		x"81",	--6579
		x"52",	--6580
		x"02",	--6581
		x"3b",	--6582
		x"00",	--6583
		x"18",	--6584
		x"60",	--6585
		x"88",	--6586
		x"00",	--6587
		x"88",	--6588
		x"02",	--6589
		x"1e",	--6590
		x"50",	--6591
		x"1f",	--6592
		x"52",	--6593
		x"b0",	--6594
		x"08",	--6595
		x"05",	--6596
		x"35",	--6597
		x"54",	--6598
		x"16",	--6599
		x"07",	--6600
		x"06",	--6601
		x"3c",	--6602
		x"3d",	--6603
		x"b0",	--6604
		x"bc",	--6605
		x"16",	--6606
		x"07",	--6607
		x"81",	--6608
		x"42",	--6609
		x"06",	--6610
		x"17",	--6611
		x"42",	--6612
		x"f4",	--6613
		x"81",	--6614
		x"40",	--6615
		x"f1",	--6616
		x"0a",	--6617
		x"0b",	--6618
		x"81",	--6619
		x"50",	--6620
		x"03",	--6621
		x"81",	--6622
		x"52",	--6623
		x"02",	--6624
		x"3b",	--6625
		x"00",	--6626
		x"19",	--6627
		x"60",	--6628
		x"89",	--6629
		x"04",	--6630
		x"89",	--6631
		x"06",	--6632
		x"30",	--6633
		x"02",	--6634
		x"1f",	--6635
		x"5c",	--6636
		x"0f",	--6637
		x"0f",	--6638
		x"3a",	--6639
		x"50",	--6640
		x"0a",	--6641
		x"0a",	--6642
		x"1a",	--6643
		x"48",	--6644
		x"81",	--6645
		x"44",	--6646
		x"16",	--6647
		x"04",	--6648
		x"17",	--6649
		x"06",	--6650
		x"1f",	--6651
		x"40",	--6652
		x"0f",	--6653
		x"0f",	--6654
		x"39",	--6655
		x"50",	--6656
		x"09",	--6657
		x"09",	--6658
		x"19",	--6659
		x"54",	--6660
		x"81",	--6661
		x"4c",	--6662
		x"28",	--6663
		x"19",	--6664
		x"02",	--6665
		x"0c",	--6666
		x"0d",	--6667
		x"0e",	--6668
		x"0f",	--6669
		x"b0",	--6670
		x"bc",	--6671
		x"0a",	--6672
		x"0b",	--6673
		x"0c",	--6674
		x"0d",	--6675
		x"0e",	--6676
		x"0f",	--6677
		x"b0",	--6678
		x"08",	--6679
		x"0c",	--6680
		x"0d",	--6681
		x"0e",	--6682
		x"0f",	--6683
		x"b0",	--6684
		x"bc",	--6685
		x"18",	--6686
		x"4c",	--6687
		x"88",	--6688
		x"00",	--6689
		x"88",	--6690
		x"02",	--6691
		x"19",	--6692
		x"44",	--6693
		x"89",	--6694
		x"04",	--6695
		x"89",	--6696
		x"06",	--6697
		x"34",	--6698
		x"35",	--6699
		x"a1",	--6700
		x"54",	--6701
		x"12",	--6702
		x"1c",	--6703
		x"40",	--6704
		x"1d",	--6705
		x"42",	--6706
		x"81",	--6707
		x"54",	--6708
		x"81",	--6709
		x"48",	--6710
		x"08",	--6711
		x"09",	--6712
		x"38",	--6713
		x"39",	--6714
		x"81",	--6715
		x"5c",	--6716
		x"81",	--6717
		x"5e",	--6718
		x"04",	--6719
		x"05",	--6720
		x"a1",	--6721
		x"48",	--6722
		x"05",	--6723
		x"04",	--6724
		x"15",	--6725
		x"a4",	--6726
		x"14",	--6727
		x"a2",	--6728
		x"1c",	--6729
		x"40",	--6730
		x"1d",	--6731
		x"42",	--6732
		x"81",	--6733
		x"54",	--6734
		x"81",	--6735
		x"48",	--6736
		x"09",	--6737
		x"0a",	--6738
		x"39",	--6739
		x"3a",	--6740
		x"81",	--6741
		x"5c",	--6742
		x"81",	--6743
		x"5e",	--6744
		x"04",	--6745
		x"05",	--6746
		x"43",	--6747
		x"1f",	--6748
		x"5c",	--6749
		x"0f",	--6750
		x"0f",	--6751
		x"3a",	--6752
		x"50",	--6753
		x"0a",	--6754
		x"0a",	--6755
		x"1a",	--6756
		x"48",	--6757
		x"81",	--6758
		x"44",	--6759
		x"16",	--6760
		x"04",	--6761
		x"17",	--6762
		x"06",	--6763
		x"1f",	--6764
		x"40",	--6765
		x"0f",	--6766
		x"0f",	--6767
		x"39",	--6768
		x"50",	--6769
		x"09",	--6770
		x"09",	--6771
		x"19",	--6772
		x"54",	--6773
		x"81",	--6774
		x"4c",	--6775
		x"28",	--6776
		x"19",	--6777
		x"02",	--6778
		x"0c",	--6779
		x"0d",	--6780
		x"0e",	--6781
		x"0f",	--6782
		x"b0",	--6783
		x"bc",	--6784
		x"0a",	--6785
		x"0b",	--6786
		x"0c",	--6787
		x"0d",	--6788
		x"0e",	--6789
		x"0f",	--6790
		x"b0",	--6791
		x"08",	--6792
		x"0c",	--6793
		x"0d",	--6794
		x"0e",	--6795
		x"0f",	--6796
		x"b0",	--6797
		x"bc",	--6798
		x"18",	--6799
		x"4c",	--6800
		x"88",	--6801
		x"00",	--6802
		x"88",	--6803
		x"02",	--6804
		x"19",	--6805
		x"44",	--6806
		x"89",	--6807
		x"04",	--6808
		x"89",	--6809
		x"06",	--6810
		x"34",	--6811
		x"35",	--6812
		x"a1",	--6813
		x"54",	--6814
		x"a1",	--6815
		x"48",	--6816
		x"05",	--6817
		x"04",	--6818
		x"15",	--6819
		x"b7",	--6820
		x"24",	--6821
		x"b5",	--6822
		x"16",	--6823
		x"40",	--6824
		x"17",	--6825
		x"42",	--6826
		x"05",	--6827
		x"0a",	--6828
		x"0b",	--6829
		x"15",	--6830
		x"1f",	--6831
		x"40",	--6832
		x"0f",	--6833
		x"0f",	--6834
		x"3d",	--6835
		x"50",	--6836
		x"0d",	--6837
		x"0f",	--6838
		x"0f",	--6839
		x"2c",	--6840
		x"1d",	--6841
		x"02",	--6842
		x"0e",	--6843
		x"0f",	--6844
		x"b0",	--6845
		x"bc",	--6846
		x"0a",	--6847
		x"0b",	--6848
		x"36",	--6849
		x"37",	--6850
		x"25",	--6851
		x"07",	--6852
		x"04",	--6853
		x"17",	--6854
		x"e7",	--6855
		x"26",	--6856
		x"e5",	--6857
		x"81",	--6858
		x"50",	--6859
		x"16",	--6860
		x"81",	--6861
		x"52",	--6862
		x"13",	--6863
		x"18",	--6864
		x"60",	--6865
		x"98",	--6866
		x"50",	--6867
		x"00",	--6868
		x"98",	--6869
		x"52",	--6870
		x"02",	--6871
		x"98",	--6872
		x"54",	--6873
		x"04",	--6874
		x"98",	--6875
		x"56",	--6876
		x"06",	--6877
		x"88",	--6878
		x"08",	--6879
		x"88",	--6880
		x"0a",	--6881
		x"1e",	--6882
		x"1d",	--6883
		x"50",	--6884
		x"1e",	--6885
		x"52",	--6886
		x"3e",	--6887
		x"00",	--6888
		x"18",	--6889
		x"60",	--6890
		x"88",	--6891
		x"00",	--6892
		x"88",	--6893
		x"02",	--6894
		x"1d",	--6895
		x"54",	--6896
		x"1e",	--6897
		x"56",	--6898
		x"3e",	--6899
		x"00",	--6900
		x"88",	--6901
		x"04",	--6902
		x"88",	--6903
		x"06",	--6904
		x"0d",	--6905
		x"0e",	--6906
		x"3e",	--6907
		x"00",	--6908
		x"88",	--6909
		x"08",	--6910
		x"88",	--6911
		x"0a",	--6912
		x"1f",	--6913
		x"58",	--6914
		x"3f",	--6915
		x"07",	--6916
		x"31",	--6917
		x"74",	--6918
		x"34",	--6919
		x"35",	--6920
		x"36",	--6921
		x"37",	--6922
		x"38",	--6923
		x"39",	--6924
		x"3a",	--6925
		x"3b",	--6926
		x"30",	--6927
		x"0b",	--6928
		x"0a",	--6929
		x"31",	--6930
		x"0c",	--6931
		x"0d",	--6932
		x"3c",	--6933
		x"3d",	--6934
		x"ff",	--6935
		x"3d",	--6936
		x"49",	--6937
		x"06",	--6938
		x"3d",	--6939
		x"4a",	--6940
		x"06",	--6941
		x"3c",	--6942
		x"d9",	--6943
		x"03",	--6944
		x"0c",	--6945
		x"0d",	--6946
		x"26",	--6947
		x"3d",	--6948
		x"80",	--6949
		x"05",	--6950
		x"0c",	--6951
		x"0d",	--6952
		x"b0",	--6953
		x"08",	--6954
		x"2f",	--6955
		x"0d",	--6956
		x"b0",	--6957
		x"ce",	--6958
		x"0a",	--6959
		x"0b",	--6960
		x"3a",	--6961
		x"03",	--6962
		x"0b",	--6963
		x"1c",	--6964
		x"04",	--6965
		x"1d",	--6966
		x"06",	--6967
		x"2e",	--6968
		x"1f",	--6969
		x"02",	--6970
		x"1a",	--6971
		x"02",	--6972
		x"0b",	--6973
		x"0e",	--6974
		x"2a",	--6975
		x"02",	--6976
		x"0b",	--6977
		x"0f",	--6978
		x"2e",	--6979
		x"1f",	--6980
		x"02",	--6981
		x"0a",	--6982
		x"0f",	--6983
		x"0b",	--6984
		x"0d",	--6985
		x"b0",	--6986
		x"ea",	--6987
		x"0e",	--6988
		x"13",	--6989
		x"b0",	--6990
		x"c4",	--6991
		x"21",	--6992
		x"02",	--6993
		x"b0",	--6994
		x"ea",	--6995
		x"3f",	--6996
		x"00",	--6997
		x"04",	--6998
		x"13",	--6999
		x"b0",	--7000
		x"c4",	--7001
		x"21",	--7002
		x"31",	--7003
		x"3a",	--7004
		x"3b",	--7005
		x"30",	--7006
		x"b0",	--7007
		x"20",	--7008
		x"30",	--7009
		x"0b",	--7010
		x"0a",	--7011
		x"09",	--7012
		x"08",	--7013
		x"07",	--7014
		x"06",	--7015
		x"05",	--7016
		x"04",	--7017
		x"31",	--7018
		x"08",	--7019
		x"09",	--7020
		x"81",	--7021
		x"00",	--7022
		x"81",	--7023
		x"02",	--7024
		x"0a",	--7025
		x"0b",	--7026
		x"3a",	--7027
		x"3b",	--7028
		x"ff",	--7029
		x"3b",	--7030
		x"00",	--7031
		x"04",	--7032
		x"b0",	--7033
		x"02",	--7034
		x"0e",	--7035
		x"9b",	--7036
		x"0c",	--7037
		x"0d",	--7038
		x"0e",	--7039
		x"0f",	--7040
		x"b0",	--7041
		x"58",	--7042
		x"0a",	--7043
		x"0b",	--7044
		x"0c",	--7045
		x"0d",	--7046
		x"b0",	--7047
		x"58",	--7048
		x"06",	--7049
		x"07",	--7050
		x"3c",	--7051
		x"d3",	--7052
		x"3d",	--7053
		x"2e",	--7054
		x"0e",	--7055
		x"0f",	--7056
		x"b0",	--7057
		x"58",	--7058
		x"3c",	--7059
		x"34",	--7060
		x"3d",	--7061
		x"d7",	--7062
		x"b0",	--7063
		x"08",	--7064
		x"0c",	--7065
		x"0d",	--7066
		x"0e",	--7067
		x"0f",	--7068
		x"b0",	--7069
		x"58",	--7070
		x"3c",	--7071
		x"1b",	--7072
		x"3d",	--7073
		x"38",	--7074
		x"b0",	--7075
		x"bc",	--7076
		x"0c",	--7077
		x"0d",	--7078
		x"0e",	--7079
		x"0f",	--7080
		x"b0",	--7081
		x"58",	--7082
		x"3c",	--7083
		x"01",	--7084
		x"3d",	--7085
		x"50",	--7086
		x"b0",	--7087
		x"08",	--7088
		x"0c",	--7089
		x"0d",	--7090
		x"0e",	--7091
		x"0f",	--7092
		x"b0",	--7093
		x"58",	--7094
		x"3c",	--7095
		x"89",	--7096
		x"3d",	--7097
		x"08",	--7098
		x"b0",	--7099
		x"bc",	--7100
		x"04",	--7101
		x"05",	--7102
		x"81",	--7103
		x"1a",	--7104
		x"19",	--7105
		x"0c",	--7106
		x"0d",	--7107
		x"0e",	--7108
		x"0f",	--7109
		x"b0",	--7110
		x"58",	--7111
		x"3c",	--7112
		x"ab",	--7113
		x"3d",	--7114
		x"2a",	--7115
		x"b0",	--7116
		x"08",	--7117
		x"0c",	--7118
		x"0d",	--7119
		x"0e",	--7120
		x"0f",	--7121
		x"b0",	--7122
		x"58",	--7123
		x"0c",	--7124
		x"0d",	--7125
		x"0e",	--7126
		x"0f",	--7127
		x"b0",	--7128
		x"bc",	--7129
		x"3b",	--7130
		x"0c",	--7131
		x"3d",	--7132
		x"00",	--7133
		x"2e",	--7134
		x"1f",	--7135
		x"02",	--7136
		x"b0",	--7137
		x"58",	--7138
		x"81",	--7139
		x"04",	--7140
		x"81",	--7141
		x"06",	--7142
		x"0c",	--7143
		x"0d",	--7144
		x"0e",	--7145
		x"0f",	--7146
		x"b0",	--7147
		x"58",	--7148
		x"0c",	--7149
		x"0d",	--7150
		x"1e",	--7151
		x"04",	--7152
		x"1f",	--7153
		x"06",	--7154
		x"b0",	--7155
		x"08",	--7156
		x"0c",	--7157
		x"0d",	--7158
		x"0e",	--7159
		x"0f",	--7160
		x"b0",	--7161
		x"58",	--7162
		x"2c",	--7163
		x"1d",	--7164
		x"02",	--7165
		x"b0",	--7166
		x"08",	--7167
		x"0a",	--7168
		x"0b",	--7169
		x"3c",	--7170
		x"ab",	--7171
		x"3d",	--7172
		x"2a",	--7173
		x"0e",	--7174
		x"0f",	--7175
		x"b0",	--7176
		x"58",	--7177
		x"0c",	--7178
		x"0d",	--7179
		x"0e",	--7180
		x"0f",	--7181
		x"b0",	--7182
		x"bc",	--7183
		x"0c",	--7184
		x"0d",	--7185
		x"0e",	--7186
		x"0f",	--7187
		x"b0",	--7188
		x"08",	--7189
		x"08",	--7190
		x"09",	--7191
		x"0e",	--7192
		x"0f",	--7193
		x"31",	--7194
		x"34",	--7195
		x"35",	--7196
		x"36",	--7197
		x"37",	--7198
		x"38",	--7199
		x"39",	--7200
		x"3a",	--7201
		x"3b",	--7202
		x"30",	--7203
		x"0b",	--7204
		x"0a",	--7205
		x"09",	--7206
		x"08",	--7207
		x"07",	--7208
		x"07",	--7209
		x"08",	--7210
		x"09",	--7211
		x"0c",	--7212
		x"0d",	--7213
		x"3c",	--7214
		x"3d",	--7215
		x"ff",	--7216
		x"0c",	--7217
		x"02",	--7218
		x"0d",	--7219
		x"a8",	--7220
		x"3d",	--7221
		x"80",	--7222
		x"05",	--7223
		x"0c",	--7224
		x"0d",	--7225
		x"b0",	--7226
		x"bc",	--7227
		x"a0",	--7228
		x"3d",	--7229
		x"80",	--7230
		x"0a",	--7231
		x"0c",	--7232
		x"0d",	--7233
		x"7e",	--7234
		x"07",	--7235
		x"12",	--7236
		x"0d",	--7237
		x"0c",	--7238
		x"7e",	--7239
		x"fb",	--7240
		x"1b",	--7241
		x"0c",	--7242
		x"3d",	--7243
		x"00",	--7244
		x"b0",	--7245
		x"58",	--7246
		x"08",	--7247
		x"09",	--7248
		x"0a",	--7249
		x"0b",	--7250
		x"0a",	--7251
		x"3b",	--7252
		x"80",	--7253
		x"0c",	--7254
		x"0d",	--7255
		x"8d",	--7256
		x"8d",	--7257
		x"8d",	--7258
		x"8d",	--7259
		x"7e",	--7260
		x"07",	--7261
		x"0d",	--7262
		x"0c",	--7263
		x"7e",	--7264
		x"fc",	--7265
		x"3c",	--7266
		x"e7",	--7267
		x"3d",	--7268
		x"0a",	--7269
		x"0e",	--7270
		x"8e",	--7271
		x"8e",	--7272
		x"8e",	--7273
		x"8e",	--7274
		x"0b",	--7275
		x"0c",	--7276
		x"0d",	--7277
		x"0d",	--7278
		x"15",	--7279
		x"03",	--7280
		x"3c",	--7281
		x"ff",	--7282
		x"11",	--7283
		x"3a",	--7284
		x"ca",	--7285
		x"3b",	--7286
		x"49",	--7287
		x"0f",	--7288
		x"04",	--7289
		x"3a",	--7290
		x"ca",	--7291
		x"3b",	--7292
		x"49",	--7293
		x"3c",	--7294
		x"ca",	--7295
		x"3d",	--7296
		x"49",	--7297
		x"0e",	--7298
		x"0f",	--7299
		x"56",	--7300
		x"0d",	--7301
		x"14",	--7302
		x"02",	--7303
		x"1c",	--7304
		x"11",	--7305
		x"0a",	--7306
		x"0b",	--7307
		x"0b",	--7308
		x"7f",	--7309
		x"07",	--7310
		x"0a",	--7311
		x"0b",	--7312
		x"7f",	--7313
		x"fc",	--7314
		x"38",	--7315
		x"39",	--7316
		x"7f",	--7317
		x"08",	--7318
		x"09",	--7319
		x"0e",	--7320
		x"0f",	--7321
		x"42",	--7322
		x"3d",	--7323
		x"05",	--7324
		x"0d",	--7325
		x"27",	--7326
		x"3c",	--7327
		x"ea",	--7328
		x"24",	--7329
		x"0d",	--7330
		x"3d",	--7331
		x"00",	--7332
		x"37",	--7333
		x"31",	--7334
		x"0f",	--7335
		x"3e",	--7336
		x"ca",	--7337
		x"3f",	--7338
		x"49",	--7339
		x"0d",	--7340
		x"04",	--7341
		x"3e",	--7342
		x"ca",	--7343
		x"3f",	--7344
		x"49",	--7345
		x"3c",	--7346
		x"ca",	--7347
		x"3d",	--7348
		x"49",	--7349
		x"24",	--7350
		x"3e",	--7351
		x"60",	--7352
		x"3f",	--7353
		x"a2",	--7354
		x"0d",	--7355
		x"04",	--7356
		x"3e",	--7357
		x"60",	--7358
		x"3f",	--7359
		x"a2",	--7360
		x"3c",	--7361
		x"60",	--7362
		x"3d",	--7363
		x"a2",	--7364
		x"15",	--7365
		x"0a",	--7366
		x"0b",	--7367
		x"0b",	--7368
		x"3b",	--7369
		x"19",	--7370
		x"7f",	--7371
		x"07",	--7372
		x"0a",	--7373
		x"0b",	--7374
		x"7f",	--7375
		x"fc",	--7376
		x"0e",	--7377
		x"0f",	--7378
		x"3e",	--7379
		x"3f",	--7380
		x"7f",	--7381
		x"0e",	--7382
		x"0f",	--7383
		x"0c",	--7384
		x"3d",	--7385
		x"00",	--7386
		x"b0",	--7387
		x"58",	--7388
		x"37",	--7389
		x"38",	--7390
		x"39",	--7391
		x"3a",	--7392
		x"3b",	--7393
		x"30",	--7394
		x"b0",	--7395
		x"48",	--7396
		x"30",	--7397
		x"0b",	--7398
		x"0a",	--7399
		x"09",	--7400
		x"08",	--7401
		x"07",	--7402
		x"06",	--7403
		x"05",	--7404
		x"04",	--7405
		x"21",	--7406
		x"06",	--7407
		x"07",	--7408
		x"08",	--7409
		x"09",	--7410
		x"38",	--7411
		x"39",	--7412
		x"ff",	--7413
		x"0c",	--7414
		x"0d",	--7415
		x"7a",	--7416
		x"07",	--7417
		x"12",	--7418
		x"0d",	--7419
		x"0c",	--7420
		x"7a",	--7421
		x"fb",	--7422
		x"3c",	--7423
		x"81",	--7424
		x"3d",	--7425
		x"0d",	--7426
		x"05",	--7427
		x"1d",	--7428
		x"57",	--7429
		x"3c",	--7430
		x"17",	--7431
		x"54",	--7432
		x"0a",	--7433
		x"0b",	--7434
		x"0d",	--7435
		x"09",	--7436
		x"81",	--7437
		x"00",	--7438
		x"38",	--7439
		x"39",	--7440
		x"7f",	--7441
		x"6d",	--7442
		x"7d",	--7443
		x"1f",	--7444
		x"1d",	--7445
		x"3c",	--7446
		x"ca",	--7447
		x"3d",	--7448
		x"49",	--7449
		x"b0",	--7450
		x"bc",	--7451
		x"0c",	--7452
		x"0d",	--7453
		x"b0",	--7454
		x"1c",	--7455
		x"0f",	--7456
		x"43",	--7457
		x"42",	--7458
		x"0b",	--7459
		x"03",	--7460
		x"0a",	--7461
		x"0b",	--7462
		x"3d",	--7463
		x"08",	--7464
		x"02",	--7465
		x"09",	--7466
		x"39",	--7467
		x"0a",	--7468
		x"3b",	--7469
		x"80",	--7470
		x"35",	--7471
		x"09",	--7472
		x"08",	--7473
		x"7d",	--7474
		x"4d",	--7475
		x"fb",	--7476
		x"04",	--7477
		x"05",	--7478
		x"04",	--7479
		x"05",	--7480
		x"04",	--7481
		x"02",	--7482
		x"05",	--7483
		x"2a",	--7484
		x"3c",	--7485
		x"ca",	--7486
		x"3d",	--7487
		x"49",	--7488
		x"b0",	--7489
		x"bc",	--7490
		x"0c",	--7491
		x"0d",	--7492
		x"b0",	--7493
		x"1c",	--7494
		x"0f",	--7495
		x"1c",	--7496
		x"1b",	--7497
		x"07",	--7498
		x"0e",	--7499
		x"0a",	--7500
		x"3b",	--7501
		x"80",	--7502
		x"6c",	--7503
		x"7c",	--7504
		x"1f",	--7505
		x"4c",	--7506
		x"04",	--7507
		x"0b",	--7508
		x"0a",	--7509
		x"7c",	--7510
		x"fa",	--7511
		x"0a",	--7512
		x"0b",	--7513
		x"0a",	--7514
		x"0b",	--7515
		x"08",	--7516
		x"39",	--7517
		x"80",	--7518
		x"07",	--7519
		x"0c",	--7520
		x"0d",	--7521
		x"b0",	--7522
		x"bc",	--7523
		x"02",	--7524
		x"0e",	--7525
		x"0f",	--7526
		x"21",	--7527
		x"34",	--7528
		x"35",	--7529
		x"36",	--7530
		x"37",	--7531
		x"38",	--7532
		x"39",	--7533
		x"3a",	--7534
		x"3b",	--7535
		x"30",	--7536
		x"b0",	--7537
		x"cc",	--7538
		x"30",	--7539
		x"0b",	--7540
		x"0a",	--7541
		x"0a",	--7542
		x"0b",	--7543
		x"0c",	--7544
		x"3d",	--7545
		x"00",	--7546
		x"b0",	--7547
		x"6c",	--7548
		x"0f",	--7549
		x"07",	--7550
		x"0e",	--7551
		x"0f",	--7552
		x"b0",	--7553
		x"02",	--7554
		x"3a",	--7555
		x"3b",	--7556
		x"30",	--7557
		x"0c",	--7558
		x"3d",	--7559
		x"00",	--7560
		x"0e",	--7561
		x"0f",	--7562
		x"b0",	--7563
		x"08",	--7564
		x"b0",	--7565
		x"02",	--7566
		x"0e",	--7567
		x"3f",	--7568
		x"00",	--7569
		x"3a",	--7570
		x"3b",	--7571
		x"30",	--7572
		x"0b",	--7573
		x"0a",	--7574
		x"09",	--7575
		x"08",	--7576
		x"07",	--7577
		x"06",	--7578
		x"05",	--7579
		x"04",	--7580
		x"31",	--7581
		x"fa",	--7582
		x"08",	--7583
		x"6b",	--7584
		x"6b",	--7585
		x"67",	--7586
		x"6c",	--7587
		x"6c",	--7588
		x"e9",	--7589
		x"6b",	--7590
		x"02",	--7591
		x"30",	--7592
		x"aa",	--7593
		x"6c",	--7594
		x"e3",	--7595
		x"6c",	--7596
		x"bb",	--7597
		x"6b",	--7598
		x"df",	--7599
		x"91",	--7600
		x"02",	--7601
		x"00",	--7602
		x"1b",	--7603
		x"02",	--7604
		x"14",	--7605
		x"04",	--7606
		x"15",	--7607
		x"06",	--7608
		x"16",	--7609
		x"04",	--7610
		x"17",	--7611
		x"06",	--7612
		x"2c",	--7613
		x"0c",	--7614
		x"09",	--7615
		x"0c",	--7616
		x"bf",	--7617
		x"39",	--7618
		x"20",	--7619
		x"50",	--7620
		x"1c",	--7621
		x"d7",	--7622
		x"81",	--7623
		x"02",	--7624
		x"81",	--7625
		x"04",	--7626
		x"4c",	--7627
		x"7c",	--7628
		x"1f",	--7629
		x"0b",	--7630
		x"0a",	--7631
		x"0b",	--7632
		x"12",	--7633
		x"0b",	--7634
		x"0a",	--7635
		x"7c",	--7636
		x"fb",	--7637
		x"81",	--7638
		x"02",	--7639
		x"81",	--7640
		x"04",	--7641
		x"1c",	--7642
		x"0d",	--7643
		x"79",	--7644
		x"1f",	--7645
		x"04",	--7646
		x"0c",	--7647
		x"0d",	--7648
		x"79",	--7649
		x"fc",	--7650
		x"3c",	--7651
		x"3d",	--7652
		x"0c",	--7653
		x"0d",	--7654
		x"1a",	--7655
		x"0b",	--7656
		x"0c",	--7657
		x"02",	--7658
		x"0d",	--7659
		x"e5",	--7660
		x"16",	--7661
		x"02",	--7662
		x"17",	--7663
		x"04",	--7664
		x"06",	--7665
		x"07",	--7666
		x"5f",	--7667
		x"01",	--7668
		x"5f",	--7669
		x"01",	--7670
		x"28",	--7671
		x"c8",	--7672
		x"01",	--7673
		x"a8",	--7674
		x"02",	--7675
		x"0e",	--7676
		x"0f",	--7677
		x"0e",	--7678
		x"0f",	--7679
		x"88",	--7680
		x"04",	--7681
		x"88",	--7682
		x"06",	--7683
		x"f8",	--7684
		x"03",	--7685
		x"00",	--7686
		x"0f",	--7687
		x"4d",	--7688
		x"0f",	--7689
		x"31",	--7690
		x"06",	--7691
		x"34",	--7692
		x"35",	--7693
		x"36",	--7694
		x"37",	--7695
		x"38",	--7696
		x"39",	--7697
		x"3a",	--7698
		x"3b",	--7699
		x"30",	--7700
		x"2b",	--7701
		x"67",	--7702
		x"81",	--7703
		x"00",	--7704
		x"04",	--7705
		x"05",	--7706
		x"5f",	--7707
		x"01",	--7708
		x"5f",	--7709
		x"01",	--7710
		x"d8",	--7711
		x"4f",	--7712
		x"68",	--7713
		x"0e",	--7714
		x"0f",	--7715
		x"0e",	--7716
		x"0f",	--7717
		x"0f",	--7718
		x"69",	--7719
		x"c8",	--7720
		x"01",	--7721
		x"a8",	--7722
		x"02",	--7723
		x"88",	--7724
		x"04",	--7725
		x"88",	--7726
		x"06",	--7727
		x"0c",	--7728
		x"0d",	--7729
		x"3c",	--7730
		x"3d",	--7731
		x"3d",	--7732
		x"ff",	--7733
		x"05",	--7734
		x"3d",	--7735
		x"00",	--7736
		x"17",	--7737
		x"3c",	--7738
		x"15",	--7739
		x"1b",	--7740
		x"02",	--7741
		x"3b",	--7742
		x"0e",	--7743
		x"0f",	--7744
		x"0a",	--7745
		x"3b",	--7746
		x"0c",	--7747
		x"0d",	--7748
		x"3c",	--7749
		x"3d",	--7750
		x"3d",	--7751
		x"ff",	--7752
		x"f5",	--7753
		x"3c",	--7754
		x"88",	--7755
		x"04",	--7756
		x"88",	--7757
		x"06",	--7758
		x"88",	--7759
		x"02",	--7760
		x"f8",	--7761
		x"03",	--7762
		x"00",	--7763
		x"0f",	--7764
		x"b3",	--7765
		x"0c",	--7766
		x"0d",	--7767
		x"1c",	--7768
		x"0d",	--7769
		x"12",	--7770
		x"0f",	--7771
		x"0e",	--7772
		x"0a",	--7773
		x"0b",	--7774
		x"0a",	--7775
		x"0b",	--7776
		x"88",	--7777
		x"04",	--7778
		x"88",	--7779
		x"06",	--7780
		x"98",	--7781
		x"02",	--7782
		x"0f",	--7783
		x"a1",	--7784
		x"6b",	--7785
		x"9f",	--7786
		x"ad",	--7787
		x"00",	--7788
		x"9d",	--7789
		x"02",	--7790
		x"02",	--7791
		x"9d",	--7792
		x"04",	--7793
		x"04",	--7794
		x"9d",	--7795
		x"06",	--7796
		x"06",	--7797
		x"5e",	--7798
		x"01",	--7799
		x"5e",	--7800
		x"01",	--7801
		x"cd",	--7802
		x"01",	--7803
		x"0f",	--7804
		x"8c",	--7805
		x"06",	--7806
		x"07",	--7807
		x"9a",	--7808
		x"39",	--7809
		x"19",	--7810
		x"39",	--7811
		x"20",	--7812
		x"8f",	--7813
		x"3e",	--7814
		x"3c",	--7815
		x"b6",	--7816
		x"c1",	--7817
		x"0e",	--7818
		x"0f",	--7819
		x"0e",	--7820
		x"0f",	--7821
		x"97",	--7822
		x"0f",	--7823
		x"79",	--7824
		x"d8",	--7825
		x"01",	--7826
		x"a8",	--7827
		x"02",	--7828
		x"3e",	--7829
		x"3f",	--7830
		x"1e",	--7831
		x"0f",	--7832
		x"88",	--7833
		x"04",	--7834
		x"88",	--7835
		x"06",	--7836
		x"92",	--7837
		x"0c",	--7838
		x"7b",	--7839
		x"81",	--7840
		x"00",	--7841
		x"81",	--7842
		x"02",	--7843
		x"81",	--7844
		x"04",	--7845
		x"4d",	--7846
		x"7d",	--7847
		x"1f",	--7848
		x"0c",	--7849
		x"4b",	--7850
		x"0c",	--7851
		x"0d",	--7852
		x"12",	--7853
		x"0d",	--7854
		x"0c",	--7855
		x"7b",	--7856
		x"fb",	--7857
		x"81",	--7858
		x"02",	--7859
		x"81",	--7860
		x"04",	--7861
		x"1c",	--7862
		x"0d",	--7863
		x"79",	--7864
		x"1f",	--7865
		x"04",	--7866
		x"0c",	--7867
		x"0d",	--7868
		x"79",	--7869
		x"fc",	--7870
		x"3c",	--7871
		x"3d",	--7872
		x"0c",	--7873
		x"0d",	--7874
		x"1a",	--7875
		x"0b",	--7876
		x"0c",	--7877
		x"04",	--7878
		x"0d",	--7879
		x"02",	--7880
		x"0a",	--7881
		x"0b",	--7882
		x"14",	--7883
		x"02",	--7884
		x"15",	--7885
		x"04",	--7886
		x"04",	--7887
		x"05",	--7888
		x"49",	--7889
		x"0a",	--7890
		x"0b",	--7891
		x"18",	--7892
		x"6c",	--7893
		x"33",	--7894
		x"df",	--7895
		x"01",	--7896
		x"01",	--7897
		x"2f",	--7898
		x"3f",	--7899
		x"3e",	--7900
		x"2c",	--7901
		x"31",	--7902
		x"e0",	--7903
		x"81",	--7904
		x"04",	--7905
		x"81",	--7906
		x"06",	--7907
		x"81",	--7908
		x"00",	--7909
		x"81",	--7910
		x"02",	--7911
		x"0e",	--7912
		x"3e",	--7913
		x"18",	--7914
		x"0f",	--7915
		x"2f",	--7916
		x"b0",	--7917
		x"c4",	--7918
		x"0e",	--7919
		x"3e",	--7920
		x"10",	--7921
		x"0f",	--7922
		x"b0",	--7923
		x"c4",	--7924
		x"0d",	--7925
		x"3d",	--7926
		x"0e",	--7927
		x"3e",	--7928
		x"10",	--7929
		x"0f",	--7930
		x"3f",	--7931
		x"18",	--7932
		x"b0",	--7933
		x"2a",	--7934
		x"b0",	--7935
		x"e6",	--7936
		x"31",	--7937
		x"20",	--7938
		x"30",	--7939
		x"31",	--7940
		x"e0",	--7941
		x"81",	--7942
		x"04",	--7943
		x"81",	--7944
		x"06",	--7945
		x"81",	--7946
		x"00",	--7947
		x"81",	--7948
		x"02",	--7949
		x"0e",	--7950
		x"3e",	--7951
		x"18",	--7952
		x"0f",	--7953
		x"2f",	--7954
		x"b0",	--7955
		x"c4",	--7956
		x"0e",	--7957
		x"3e",	--7958
		x"10",	--7959
		x"0f",	--7960
		x"b0",	--7961
		x"c4",	--7962
		x"d1",	--7963
		x"11",	--7964
		x"0d",	--7965
		x"3d",	--7966
		x"0e",	--7967
		x"3e",	--7968
		x"10",	--7969
		x"0f",	--7970
		x"3f",	--7971
		x"18",	--7972
		x"b0",	--7973
		x"2a",	--7974
		x"b0",	--7975
		x"e6",	--7976
		x"31",	--7977
		x"20",	--7978
		x"30",	--7979
		x"0b",	--7980
		x"0a",	--7981
		x"09",	--7982
		x"08",	--7983
		x"07",	--7984
		x"06",	--7985
		x"05",	--7986
		x"04",	--7987
		x"31",	--7988
		x"dc",	--7989
		x"81",	--7990
		x"04",	--7991
		x"81",	--7992
		x"06",	--7993
		x"81",	--7994
		x"00",	--7995
		x"81",	--7996
		x"02",	--7997
		x"0e",	--7998
		x"3e",	--7999
		x"18",	--8000
		x"0f",	--8001
		x"2f",	--8002
		x"b0",	--8003
		x"c4",	--8004
		x"0e",	--8005
		x"3e",	--8006
		x"10",	--8007
		x"0f",	--8008
		x"b0",	--8009
		x"c4",	--8010
		x"5f",	--8011
		x"18",	--8012
		x"6f",	--8013
		x"b6",	--8014
		x"5e",	--8015
		x"10",	--8016
		x"6e",	--8017
		x"d9",	--8018
		x"6f",	--8019
		x"ae",	--8020
		x"6e",	--8021
		x"e2",	--8022
		x"6f",	--8023
		x"ac",	--8024
		x"6e",	--8025
		x"d1",	--8026
		x"14",	--8027
		x"1c",	--8028
		x"15",	--8029
		x"1e",	--8030
		x"18",	--8031
		x"14",	--8032
		x"19",	--8033
		x"16",	--8034
		x"3c",	--8035
		x"20",	--8036
		x"0e",	--8037
		x"0f",	--8038
		x"06",	--8039
		x"07",	--8040
		x"81",	--8041
		x"20",	--8042
		x"81",	--8043
		x"22",	--8044
		x"0a",	--8045
		x"0b",	--8046
		x"81",	--8047
		x"20",	--8048
		x"08",	--8049
		x"08",	--8050
		x"09",	--8051
		x"12",	--8052
		x"05",	--8053
		x"04",	--8054
		x"b1",	--8055
		x"20",	--8056
		x"19",	--8057
		x"14",	--8058
		x"0d",	--8059
		x"0a",	--8060
		x"0b",	--8061
		x"0e",	--8062
		x"0f",	--8063
		x"1c",	--8064
		x"0d",	--8065
		x"0b",	--8066
		x"03",	--8067
		x"0b",	--8068
		x"0c",	--8069
		x"0d",	--8070
		x"0e",	--8071
		x"0f",	--8072
		x"06",	--8073
		x"07",	--8074
		x"09",	--8075
		x"e5",	--8076
		x"16",	--8077
		x"07",	--8078
		x"e2",	--8079
		x"0a",	--8080
		x"f5",	--8081
		x"f2",	--8082
		x"81",	--8083
		x"20",	--8084
		x"81",	--8085
		x"22",	--8086
		x"0c",	--8087
		x"1a",	--8088
		x"1a",	--8089
		x"1a",	--8090
		x"12",	--8091
		x"06",	--8092
		x"26",	--8093
		x"81",	--8094
		x"0a",	--8095
		x"5d",	--8096
		x"d1",	--8097
		x"11",	--8098
		x"19",	--8099
		x"83",	--8100
		x"c1",	--8101
		x"09",	--8102
		x"0c",	--8103
		x"3c",	--8104
		x"3f",	--8105
		x"00",	--8106
		x"18",	--8107
		x"1d",	--8108
		x"0a",	--8109
		x"3d",	--8110
		x"1a",	--8111
		x"20",	--8112
		x"1b",	--8113
		x"22",	--8114
		x"0c",	--8115
		x"0e",	--8116
		x"0f",	--8117
		x"0b",	--8118
		x"2a",	--8119
		x"0a",	--8120
		x"0b",	--8121
		x"3d",	--8122
		x"3f",	--8123
		x"00",	--8124
		x"f5",	--8125
		x"81",	--8126
		x"20",	--8127
		x"81",	--8128
		x"22",	--8129
		x"81",	--8130
		x"0a",	--8131
		x"0c",	--8132
		x"0d",	--8133
		x"3c",	--8134
		x"7f",	--8135
		x"0d",	--8136
		x"3c",	--8137
		x"40",	--8138
		x"44",	--8139
		x"81",	--8140
		x"0c",	--8141
		x"81",	--8142
		x"0e",	--8143
		x"f1",	--8144
		x"03",	--8145
		x"08",	--8146
		x"0f",	--8147
		x"3f",	--8148
		x"b0",	--8149
		x"e6",	--8150
		x"31",	--8151
		x"24",	--8152
		x"34",	--8153
		x"35",	--8154
		x"36",	--8155
		x"37",	--8156
		x"38",	--8157
		x"39",	--8158
		x"3a",	--8159
		x"3b",	--8160
		x"30",	--8161
		x"1e",	--8162
		x"0f",	--8163
		x"d3",	--8164
		x"3a",	--8165
		x"03",	--8166
		x"08",	--8167
		x"1e",	--8168
		x"10",	--8169
		x"1c",	--8170
		x"20",	--8171
		x"1d",	--8172
		x"22",	--8173
		x"12",	--8174
		x"0d",	--8175
		x"0c",	--8176
		x"06",	--8177
		x"07",	--8178
		x"06",	--8179
		x"37",	--8180
		x"00",	--8181
		x"81",	--8182
		x"20",	--8183
		x"81",	--8184
		x"22",	--8185
		x"12",	--8186
		x"0f",	--8187
		x"0e",	--8188
		x"1a",	--8189
		x"0f",	--8190
		x"e7",	--8191
		x"81",	--8192
		x"0a",	--8193
		x"a6",	--8194
		x"6e",	--8195
		x"36",	--8196
		x"5f",	--8197
		x"d1",	--8198
		x"11",	--8199
		x"19",	--8200
		x"20",	--8201
		x"c1",	--8202
		x"19",	--8203
		x"0f",	--8204
		x"3f",	--8205
		x"18",	--8206
		x"c5",	--8207
		x"0d",	--8208
		x"ba",	--8209
		x"0c",	--8210
		x"0d",	--8211
		x"3c",	--8212
		x"80",	--8213
		x"0d",	--8214
		x"0c",	--8215
		x"b3",	--8216
		x"0d",	--8217
		x"b1",	--8218
		x"81",	--8219
		x"20",	--8220
		x"03",	--8221
		x"81",	--8222
		x"22",	--8223
		x"ab",	--8224
		x"3e",	--8225
		x"40",	--8226
		x"0f",	--8227
		x"3e",	--8228
		x"80",	--8229
		x"3f",	--8230
		x"a4",	--8231
		x"4d",	--8232
		x"7b",	--8233
		x"4f",	--8234
		x"de",	--8235
		x"5f",	--8236
		x"d1",	--8237
		x"11",	--8238
		x"19",	--8239
		x"06",	--8240
		x"c1",	--8241
		x"11",	--8242
		x"0f",	--8243
		x"3f",	--8244
		x"10",	--8245
		x"9e",	--8246
		x"4f",	--8247
		x"f8",	--8248
		x"6f",	--8249
		x"f1",	--8250
		x"3f",	--8251
		x"3e",	--8252
		x"97",	--8253
		x"0b",	--8254
		x"0a",	--8255
		x"09",	--8256
		x"08",	--8257
		x"07",	--8258
		x"31",	--8259
		x"e8",	--8260
		x"81",	--8261
		x"04",	--8262
		x"81",	--8263
		x"06",	--8264
		x"81",	--8265
		x"00",	--8266
		x"81",	--8267
		x"02",	--8268
		x"0e",	--8269
		x"3e",	--8270
		x"10",	--8271
		x"0f",	--8272
		x"2f",	--8273
		x"b0",	--8274
		x"c4",	--8275
		x"0e",	--8276
		x"3e",	--8277
		x"0f",	--8278
		x"b0",	--8279
		x"c4",	--8280
		x"5f",	--8281
		x"10",	--8282
		x"6f",	--8283
		x"5d",	--8284
		x"5e",	--8285
		x"08",	--8286
		x"6e",	--8287
		x"82",	--8288
		x"d1",	--8289
		x"09",	--8290
		x"11",	--8291
		x"6f",	--8292
		x"58",	--8293
		x"6f",	--8294
		x"56",	--8295
		x"6e",	--8296
		x"6f",	--8297
		x"6e",	--8298
		x"4c",	--8299
		x"1d",	--8300
		x"12",	--8301
		x"1d",	--8302
		x"0a",	--8303
		x"81",	--8304
		x"12",	--8305
		x"1e",	--8306
		x"14",	--8307
		x"1f",	--8308
		x"16",	--8309
		x"18",	--8310
		x"0c",	--8311
		x"19",	--8312
		x"0e",	--8313
		x"0f",	--8314
		x"1e",	--8315
		x"0e",	--8316
		x"0f",	--8317
		x"3d",	--8318
		x"81",	--8319
		x"12",	--8320
		x"37",	--8321
		x"1f",	--8322
		x"0c",	--8323
		x"3d",	--8324
		x"00",	--8325
		x"0a",	--8326
		x"0b",	--8327
		x"0b",	--8328
		x"0a",	--8329
		x"0b",	--8330
		x"0e",	--8331
		x"0f",	--8332
		x"12",	--8333
		x"0d",	--8334
		x"0c",	--8335
		x"0e",	--8336
		x"0f",	--8337
		x"37",	--8338
		x"0b",	--8339
		x"0f",	--8340
		x"f7",	--8341
		x"f2",	--8342
		x"0e",	--8343
		x"f4",	--8344
		x"ef",	--8345
		x"09",	--8346
		x"e5",	--8347
		x"0e",	--8348
		x"e3",	--8349
		x"dd",	--8350
		x"0c",	--8351
		x"0d",	--8352
		x"3c",	--8353
		x"7f",	--8354
		x"0d",	--8355
		x"3c",	--8356
		x"40",	--8357
		x"1c",	--8358
		x"81",	--8359
		x"14",	--8360
		x"81",	--8361
		x"16",	--8362
		x"0f",	--8363
		x"3f",	--8364
		x"10",	--8365
		x"b0",	--8366
		x"e6",	--8367
		x"31",	--8368
		x"18",	--8369
		x"37",	--8370
		x"38",	--8371
		x"39",	--8372
		x"3a",	--8373
		x"3b",	--8374
		x"30",	--8375
		x"e1",	--8376
		x"10",	--8377
		x"0f",	--8378
		x"3f",	--8379
		x"10",	--8380
		x"f0",	--8381
		x"4f",	--8382
		x"fa",	--8383
		x"3f",	--8384
		x"3e",	--8385
		x"eb",	--8386
		x"0d",	--8387
		x"e2",	--8388
		x"0c",	--8389
		x"0d",	--8390
		x"3c",	--8391
		x"80",	--8392
		x"0d",	--8393
		x"0c",	--8394
		x"db",	--8395
		x"0d",	--8396
		x"d9",	--8397
		x"0e",	--8398
		x"02",	--8399
		x"0f",	--8400
		x"d5",	--8401
		x"3a",	--8402
		x"40",	--8403
		x"0b",	--8404
		x"3a",	--8405
		x"80",	--8406
		x"3b",	--8407
		x"ce",	--8408
		x"81",	--8409
		x"14",	--8410
		x"81",	--8411
		x"16",	--8412
		x"81",	--8413
		x"12",	--8414
		x"0f",	--8415
		x"3f",	--8416
		x"10",	--8417
		x"cb",	--8418
		x"0f",	--8419
		x"3f",	--8420
		x"c8",	--8421
		x"31",	--8422
		x"e8",	--8423
		x"81",	--8424
		x"04",	--8425
		x"81",	--8426
		x"06",	--8427
		x"81",	--8428
		x"00",	--8429
		x"81",	--8430
		x"02",	--8431
		x"0e",	--8432
		x"3e",	--8433
		x"10",	--8434
		x"0f",	--8435
		x"2f",	--8436
		x"b0",	--8437
		x"c4",	--8438
		x"0e",	--8439
		x"3e",	--8440
		x"0f",	--8441
		x"b0",	--8442
		x"c4",	--8443
		x"e1",	--8444
		x"10",	--8445
		x"0d",	--8446
		x"e1",	--8447
		x"08",	--8448
		x"0a",	--8449
		x"0e",	--8450
		x"3e",	--8451
		x"0f",	--8452
		x"3f",	--8453
		x"10",	--8454
		x"b0",	--8455
		x"e8",	--8456
		x"31",	--8457
		x"18",	--8458
		x"30",	--8459
		x"1f",	--8460
		x"fb",	--8461
		x"31",	--8462
		x"e8",	--8463
		x"81",	--8464
		x"04",	--8465
		x"81",	--8466
		x"06",	--8467
		x"81",	--8468
		x"00",	--8469
		x"81",	--8470
		x"02",	--8471
		x"0e",	--8472
		x"3e",	--8473
		x"10",	--8474
		x"0f",	--8475
		x"2f",	--8476
		x"b0",	--8477
		x"c4",	--8478
		x"0e",	--8479
		x"3e",	--8480
		x"0f",	--8481
		x"b0",	--8482
		x"c4",	--8483
		x"e1",	--8484
		x"10",	--8485
		x"0d",	--8486
		x"e1",	--8487
		x"08",	--8488
		x"0a",	--8489
		x"0e",	--8490
		x"3e",	--8491
		x"0f",	--8492
		x"3f",	--8493
		x"10",	--8494
		x"b0",	--8495
		x"e8",	--8496
		x"31",	--8497
		x"18",	--8498
		x"30",	--8499
		x"3f",	--8500
		x"fb",	--8501
		x"31",	--8502
		x"e8",	--8503
		x"81",	--8504
		x"04",	--8505
		x"81",	--8506
		x"06",	--8507
		x"81",	--8508
		x"00",	--8509
		x"81",	--8510
		x"02",	--8511
		x"0e",	--8512
		x"3e",	--8513
		x"10",	--8514
		x"0f",	--8515
		x"2f",	--8516
		x"b0",	--8517
		x"c4",	--8518
		x"0e",	--8519
		x"3e",	--8520
		x"0f",	--8521
		x"b0",	--8522
		x"c4",	--8523
		x"e1",	--8524
		x"10",	--8525
		x"0d",	--8526
		x"e1",	--8527
		x"08",	--8528
		x"0a",	--8529
		x"0e",	--8530
		x"3e",	--8531
		x"0f",	--8532
		x"3f",	--8533
		x"10",	--8534
		x"b0",	--8535
		x"e8",	--8536
		x"31",	--8537
		x"18",	--8538
		x"30",	--8539
		x"3f",	--8540
		x"fb",	--8541
		x"31",	--8542
		x"e8",	--8543
		x"81",	--8544
		x"04",	--8545
		x"81",	--8546
		x"06",	--8547
		x"81",	--8548
		x"00",	--8549
		x"81",	--8550
		x"02",	--8551
		x"0e",	--8552
		x"3e",	--8553
		x"10",	--8554
		x"0f",	--8555
		x"2f",	--8556
		x"b0",	--8557
		x"c4",	--8558
		x"0e",	--8559
		x"3e",	--8560
		x"0f",	--8561
		x"b0",	--8562
		x"c4",	--8563
		x"e1",	--8564
		x"10",	--8565
		x"0d",	--8566
		x"e1",	--8567
		x"08",	--8568
		x"0a",	--8569
		x"0e",	--8570
		x"3e",	--8571
		x"0f",	--8572
		x"3f",	--8573
		x"10",	--8574
		x"b0",	--8575
		x"e8",	--8576
		x"31",	--8577
		x"18",	--8578
		x"30",	--8579
		x"1f",	--8580
		x"fb",	--8581
		x"31",	--8582
		x"e8",	--8583
		x"81",	--8584
		x"04",	--8585
		x"81",	--8586
		x"06",	--8587
		x"81",	--8588
		x"00",	--8589
		x"81",	--8590
		x"02",	--8591
		x"0e",	--8592
		x"3e",	--8593
		x"10",	--8594
		x"0f",	--8595
		x"2f",	--8596
		x"b0",	--8597
		x"c4",	--8598
		x"0e",	--8599
		x"3e",	--8600
		x"0f",	--8601
		x"b0",	--8602
		x"c4",	--8603
		x"e1",	--8604
		x"10",	--8605
		x"0d",	--8606
		x"e1",	--8607
		x"08",	--8608
		x"0a",	--8609
		x"0e",	--8610
		x"3e",	--8611
		x"0f",	--8612
		x"3f",	--8613
		x"10",	--8614
		x"b0",	--8615
		x"e8",	--8616
		x"31",	--8617
		x"18",	--8618
		x"30",	--8619
		x"1f",	--8620
		x"fb",	--8621
		x"0b",	--8622
		x"0a",	--8623
		x"31",	--8624
		x"f1",	--8625
		x"03",	--8626
		x"00",	--8627
		x"0d",	--8628
		x"0d",	--8629
		x"0d",	--8630
		x"0d",	--8631
		x"4c",	--8632
		x"c1",	--8633
		x"01",	--8634
		x"0e",	--8635
		x"0b",	--8636
		x"0f",	--8637
		x"09",	--8638
		x"e1",	--8639
		x"00",	--8640
		x"0f",	--8641
		x"b0",	--8642
		x"e6",	--8643
		x"31",	--8644
		x"3a",	--8645
		x"3b",	--8646
		x"30",	--8647
		x"b1",	--8648
		x"1e",	--8649
		x"02",	--8650
		x"4c",	--8651
		x"1b",	--8652
		x"0a",	--8653
		x"0b",	--8654
		x"81",	--8655
		x"04",	--8656
		x"81",	--8657
		x"06",	--8658
		x"0e",	--8659
		x"0f",	--8660
		x"b0",	--8661
		x"74",	--8662
		x"3f",	--8663
		x"1f",	--8664
		x"e7",	--8665
		x"81",	--8666
		x"04",	--8667
		x"81",	--8668
		x"06",	--8669
		x"4e",	--8670
		x"7e",	--8671
		x"1f",	--8672
		x"0f",	--8673
		x"3e",	--8674
		x"1e",	--8675
		x"0e",	--8676
		x"81",	--8677
		x"02",	--8678
		x"d9",	--8679
		x"0e",	--8680
		x"10",	--8681
		x"0a",	--8682
		x"0b",	--8683
		x"3a",	--8684
		x"3b",	--8685
		x"1a",	--8686
		x"0b",	--8687
		x"de",	--8688
		x"91",	--8689
		x"04",	--8690
		x"04",	--8691
		x"91",	--8692
		x"06",	--8693
		x"06",	--8694
		x"7e",	--8695
		x"f8",	--8696
		x"e8",	--8697
		x"3f",	--8698
		x"00",	--8699
		x"ed",	--8700
		x"0e",	--8701
		x"3f",	--8702
		x"00",	--8703
		x"c3",	--8704
		x"31",	--8705
		x"f4",	--8706
		x"81",	--8707
		x"00",	--8708
		x"81",	--8709
		x"02",	--8710
		x"0e",	--8711
		x"2e",	--8712
		x"0f",	--8713
		x"b0",	--8714
		x"c4",	--8715
		x"5f",	--8716
		x"04",	--8717
		x"6f",	--8718
		x"28",	--8719
		x"27",	--8720
		x"6f",	--8721
		x"07",	--8722
		x"1d",	--8723
		x"06",	--8724
		x"0d",	--8725
		x"21",	--8726
		x"3d",	--8727
		x"1f",	--8728
		x"09",	--8729
		x"c1",	--8730
		x"05",	--8731
		x"26",	--8732
		x"3e",	--8733
		x"3f",	--8734
		x"ff",	--8735
		x"31",	--8736
		x"0c",	--8737
		x"30",	--8738
		x"1e",	--8739
		x"08",	--8740
		x"1f",	--8741
		x"0a",	--8742
		x"3c",	--8743
		x"1e",	--8744
		x"4c",	--8745
		x"4d",	--8746
		x"7d",	--8747
		x"1f",	--8748
		x"0f",	--8749
		x"c1",	--8750
		x"05",	--8751
		x"ef",	--8752
		x"3e",	--8753
		x"3f",	--8754
		x"1e",	--8755
		x"0f",	--8756
		x"31",	--8757
		x"0c",	--8758
		x"30",	--8759
		x"0e",	--8760
		x"0f",	--8761
		x"31",	--8762
		x"0c",	--8763
		x"30",	--8764
		x"12",	--8765
		x"0f",	--8766
		x"0e",	--8767
		x"7d",	--8768
		x"fb",	--8769
		x"eb",	--8770
		x"0e",	--8771
		x"3f",	--8772
		x"00",	--8773
		x"31",	--8774
		x"0c",	--8775
		x"30",	--8776
		x"0b",	--8777
		x"0a",	--8778
		x"09",	--8779
		x"08",	--8780
		x"31",	--8781
		x"0a",	--8782
		x"0b",	--8783
		x"c1",	--8784
		x"01",	--8785
		x"0e",	--8786
		x"0d",	--8787
		x"0b",	--8788
		x"0b",	--8789
		x"e1",	--8790
		x"00",	--8791
		x"0f",	--8792
		x"b0",	--8793
		x"e6",	--8794
		x"31",	--8795
		x"38",	--8796
		x"39",	--8797
		x"3a",	--8798
		x"3b",	--8799
		x"30",	--8800
		x"f1",	--8801
		x"03",	--8802
		x"00",	--8803
		x"b1",	--8804
		x"1e",	--8805
		x"02",	--8806
		x"81",	--8807
		x"04",	--8808
		x"81",	--8809
		x"06",	--8810
		x"0e",	--8811
		x"0f",	--8812
		x"b0",	--8813
		x"74",	--8814
		x"3f",	--8815
		x"0f",	--8816
		x"18",	--8817
		x"e5",	--8818
		x"81",	--8819
		x"04",	--8820
		x"81",	--8821
		x"06",	--8822
		x"4e",	--8823
		x"7e",	--8824
		x"1f",	--8825
		x"06",	--8826
		x"3e",	--8827
		x"1e",	--8828
		x"0e",	--8829
		x"81",	--8830
		x"02",	--8831
		x"d7",	--8832
		x"91",	--8833
		x"04",	--8834
		x"04",	--8835
		x"91",	--8836
		x"06",	--8837
		x"06",	--8838
		x"7e",	--8839
		x"f8",	--8840
		x"f1",	--8841
		x"0e",	--8842
		x"3e",	--8843
		x"1e",	--8844
		x"1c",	--8845
		x"0d",	--8846
		x"48",	--8847
		x"78",	--8848
		x"1f",	--8849
		x"04",	--8850
		x"0c",	--8851
		x"0d",	--8852
		x"78",	--8853
		x"fc",	--8854
		x"3c",	--8855
		x"3d",	--8856
		x"0c",	--8857
		x"0d",	--8858
		x"18",	--8859
		x"09",	--8860
		x"0c",	--8861
		x"04",	--8862
		x"0d",	--8863
		x"02",	--8864
		x"08",	--8865
		x"09",	--8866
		x"7e",	--8867
		x"1f",	--8868
		x"0e",	--8869
		x"0d",	--8870
		x"0e",	--8871
		x"0d",	--8872
		x"0e",	--8873
		x"81",	--8874
		x"04",	--8875
		x"81",	--8876
		x"06",	--8877
		x"3e",	--8878
		x"1e",	--8879
		x"0e",	--8880
		x"81",	--8881
		x"02",	--8882
		x"a4",	--8883
		x"12",	--8884
		x"0b",	--8885
		x"0a",	--8886
		x"7e",	--8887
		x"fb",	--8888
		x"ec",	--8889
		x"0b",	--8890
		x"0a",	--8891
		x"09",	--8892
		x"1f",	--8893
		x"17",	--8894
		x"3e",	--8895
		x"00",	--8896
		x"2c",	--8897
		x"3a",	--8898
		x"18",	--8899
		x"0b",	--8900
		x"39",	--8901
		x"0c",	--8902
		x"0d",	--8903
		x"4f",	--8904
		x"4f",	--8905
		x"17",	--8906
		x"3c",	--8907
		x"46",	--8908
		x"6e",	--8909
		x"0f",	--8910
		x"0a",	--8911
		x"0b",	--8912
		x"0f",	--8913
		x"39",	--8914
		x"3a",	--8915
		x"3b",	--8916
		x"30",	--8917
		x"3f",	--8918
		x"00",	--8919
		x"0f",	--8920
		x"3a",	--8921
		x"0b",	--8922
		x"39",	--8923
		x"18",	--8924
		x"0c",	--8925
		x"0d",	--8926
		x"4f",	--8927
		x"4f",	--8928
		x"e9",	--8929
		x"12",	--8930
		x"0d",	--8931
		x"0c",	--8932
		x"7f",	--8933
		x"fb",	--8934
		x"e3",	--8935
		x"3a",	--8936
		x"10",	--8937
		x"0b",	--8938
		x"39",	--8939
		x"10",	--8940
		x"ef",	--8941
		x"3a",	--8942
		x"20",	--8943
		x"0b",	--8944
		x"09",	--8945
		x"ea",	--8946
		x"0b",	--8947
		x"0a",	--8948
		x"09",	--8949
		x"08",	--8950
		x"07",	--8951
		x"0d",	--8952
		x"1e",	--8953
		x"04",	--8954
		x"1f",	--8955
		x"06",	--8956
		x"5a",	--8957
		x"01",	--8958
		x"6c",	--8959
		x"6c",	--8960
		x"70",	--8961
		x"6c",	--8962
		x"6a",	--8963
		x"6c",	--8964
		x"36",	--8965
		x"0e",	--8966
		x"32",	--8967
		x"1b",	--8968
		x"02",	--8969
		x"3b",	--8970
		x"82",	--8971
		x"6d",	--8972
		x"3b",	--8973
		x"80",	--8974
		x"5e",	--8975
		x"0c",	--8976
		x"0d",	--8977
		x"3c",	--8978
		x"7f",	--8979
		x"0d",	--8980
		x"3c",	--8981
		x"40",	--8982
		x"40",	--8983
		x"3e",	--8984
		x"3f",	--8985
		x"0f",	--8986
		x"0f",	--8987
		x"4a",	--8988
		x"0d",	--8989
		x"3d",	--8990
		x"7f",	--8991
		x"12",	--8992
		x"0f",	--8993
		x"0e",	--8994
		x"12",	--8995
		x"0f",	--8996
		x"0e",	--8997
		x"12",	--8998
		x"0f",	--8999
		x"0e",	--9000
		x"12",	--9001
		x"0f",	--9002
		x"0e",	--9003
		x"12",	--9004
		x"0f",	--9005
		x"0e",	--9006
		x"12",	--9007
		x"0f",	--9008
		x"0e",	--9009
		x"12",	--9010
		x"0f",	--9011
		x"0e",	--9012
		x"3e",	--9013
		x"3f",	--9014
		x"7f",	--9015
		x"4d",	--9016
		x"05",	--9017
		x"0f",	--9018
		x"cc",	--9019
		x"4d",	--9020
		x"0e",	--9021
		x"0f",	--9022
		x"4d",	--9023
		x"0d",	--9024
		x"0d",	--9025
		x"0d",	--9026
		x"0d",	--9027
		x"0d",	--9028
		x"0d",	--9029
		x"0d",	--9030
		x"0c",	--9031
		x"3c",	--9032
		x"7f",	--9033
		x"0c",	--9034
		x"4f",	--9035
		x"0f",	--9036
		x"0f",	--9037
		x"0f",	--9038
		x"0d",	--9039
		x"0d",	--9040
		x"0f",	--9041
		x"37",	--9042
		x"38",	--9043
		x"39",	--9044
		x"3a",	--9045
		x"3b",	--9046
		x"30",	--9047
		x"0d",	--9048
		x"be",	--9049
		x"0c",	--9050
		x"0d",	--9051
		x"3c",	--9052
		x"80",	--9053
		x"0d",	--9054
		x"0c",	--9055
		x"02",	--9056
		x"0d",	--9057
		x"b8",	--9058
		x"3e",	--9059
		x"40",	--9060
		x"0f",	--9061
		x"b4",	--9062
		x"12",	--9063
		x"0f",	--9064
		x"0e",	--9065
		x"0d",	--9066
		x"3d",	--9067
		x"80",	--9068
		x"b2",	--9069
		x"7d",	--9070
		x"0e",	--9071
		x"0f",	--9072
		x"cd",	--9073
		x"0e",	--9074
		x"3f",	--9075
		x"10",	--9076
		x"3e",	--9077
		x"3f",	--9078
		x"7f",	--9079
		x"7d",	--9080
		x"c5",	--9081
		x"37",	--9082
		x"82",	--9083
		x"07",	--9084
		x"37",	--9085
		x"1a",	--9086
		x"4f",	--9087
		x"0c",	--9088
		x"0d",	--9089
		x"4b",	--9090
		x"7b",	--9091
		x"1f",	--9092
		x"05",	--9093
		x"12",	--9094
		x"0d",	--9095
		x"0c",	--9096
		x"7b",	--9097
		x"fb",	--9098
		x"18",	--9099
		x"09",	--9100
		x"77",	--9101
		x"1f",	--9102
		x"04",	--9103
		x"08",	--9104
		x"09",	--9105
		x"77",	--9106
		x"fc",	--9107
		x"38",	--9108
		x"39",	--9109
		x"08",	--9110
		x"09",	--9111
		x"1e",	--9112
		x"0f",	--9113
		x"08",	--9114
		x"04",	--9115
		x"09",	--9116
		x"02",	--9117
		x"0e",	--9118
		x"0f",	--9119
		x"08",	--9120
		x"09",	--9121
		x"08",	--9122
		x"09",	--9123
		x"0e",	--9124
		x"0f",	--9125
		x"3e",	--9126
		x"7f",	--9127
		x"0f",	--9128
		x"3e",	--9129
		x"40",	--9130
		x"26",	--9131
		x"38",	--9132
		x"3f",	--9133
		x"09",	--9134
		x"0e",	--9135
		x"0f",	--9136
		x"12",	--9137
		x"0f",	--9138
		x"0e",	--9139
		x"12",	--9140
		x"0f",	--9141
		x"0e",	--9142
		x"12",	--9143
		x"0f",	--9144
		x"0e",	--9145
		x"12",	--9146
		x"0f",	--9147
		x"0e",	--9148
		x"12",	--9149
		x"0f",	--9150
		x"0e",	--9151
		x"12",	--9152
		x"0f",	--9153
		x"0e",	--9154
		x"12",	--9155
		x"0f",	--9156
		x"0e",	--9157
		x"3e",	--9158
		x"3f",	--9159
		x"7f",	--9160
		x"5d",	--9161
		x"39",	--9162
		x"00",	--9163
		x"72",	--9164
		x"4d",	--9165
		x"70",	--9166
		x"08",	--9167
		x"09",	--9168
		x"da",	--9169
		x"0f",	--9170
		x"d8",	--9171
		x"0e",	--9172
		x"0f",	--9173
		x"3e",	--9174
		x"80",	--9175
		x"0f",	--9176
		x"0e",	--9177
		x"04",	--9178
		x"38",	--9179
		x"40",	--9180
		x"09",	--9181
		x"d0",	--9182
		x"0f",	--9183
		x"ce",	--9184
		x"f9",	--9185
		x"0b",	--9186
		x"0a",	--9187
		x"2a",	--9188
		x"5b",	--9189
		x"02",	--9190
		x"3b",	--9191
		x"7f",	--9192
		x"1d",	--9193
		x"02",	--9194
		x"12",	--9195
		x"0d",	--9196
		x"12",	--9197
		x"0d",	--9198
		x"12",	--9199
		x"0d",	--9200
		x"12",	--9201
		x"0d",	--9202
		x"12",	--9203
		x"0d",	--9204
		x"12",	--9205
		x"0d",	--9206
		x"12",	--9207
		x"0d",	--9208
		x"4d",	--9209
		x"5f",	--9210
		x"03",	--9211
		x"3f",	--9212
		x"80",	--9213
		x"0f",	--9214
		x"0f",	--9215
		x"ce",	--9216
		x"01",	--9217
		x"0d",	--9218
		x"2d",	--9219
		x"0a",	--9220
		x"51",	--9221
		x"be",	--9222
		x"82",	--9223
		x"02",	--9224
		x"0c",	--9225
		x"0d",	--9226
		x"0c",	--9227
		x"0d",	--9228
		x"0c",	--9229
		x"0d",	--9230
		x"0c",	--9231
		x"0d",	--9232
		x"0c",	--9233
		x"0d",	--9234
		x"0c",	--9235
		x"0d",	--9236
		x"0c",	--9237
		x"0d",	--9238
		x"0c",	--9239
		x"0d",	--9240
		x"fe",	--9241
		x"03",	--9242
		x"00",	--9243
		x"3d",	--9244
		x"00",	--9245
		x"0b",	--9246
		x"3f",	--9247
		x"81",	--9248
		x"0c",	--9249
		x"0d",	--9250
		x"0a",	--9251
		x"3f",	--9252
		x"3d",	--9253
		x"00",	--9254
		x"f9",	--9255
		x"8e",	--9256
		x"02",	--9257
		x"8e",	--9258
		x"04",	--9259
		x"8e",	--9260
		x"06",	--9261
		x"3a",	--9262
		x"3b",	--9263
		x"30",	--9264
		x"3d",	--9265
		x"ff",	--9266
		x"2a",	--9267
		x"3d",	--9268
		x"81",	--9269
		x"8e",	--9270
		x"02",	--9271
		x"fe",	--9272
		x"03",	--9273
		x"00",	--9274
		x"0c",	--9275
		x"0d",	--9276
		x"0c",	--9277
		x"0d",	--9278
		x"0c",	--9279
		x"0d",	--9280
		x"0c",	--9281
		x"0d",	--9282
		x"0c",	--9283
		x"0d",	--9284
		x"0c",	--9285
		x"0d",	--9286
		x"0c",	--9287
		x"0d",	--9288
		x"0c",	--9289
		x"0d",	--9290
		x"0a",	--9291
		x"0b",	--9292
		x"0a",	--9293
		x"3b",	--9294
		x"00",	--9295
		x"8e",	--9296
		x"04",	--9297
		x"8e",	--9298
		x"06",	--9299
		x"3a",	--9300
		x"3b",	--9301
		x"30",	--9302
		x"0b",	--9303
		x"ad",	--9304
		x"ee",	--9305
		x"00",	--9306
		x"3a",	--9307
		x"3b",	--9308
		x"30",	--9309
		x"0a",	--9310
		x"0c",	--9311
		x"0c",	--9312
		x"0d",	--9313
		x"0c",	--9314
		x"3d",	--9315
		x"10",	--9316
		x"0c",	--9317
		x"02",	--9318
		x"0d",	--9319
		x"08",	--9320
		x"de",	--9321
		x"00",	--9322
		x"e4",	--9323
		x"0b",	--9324
		x"f2",	--9325
		x"ee",	--9326
		x"00",	--9327
		x"e3",	--9328
		x"ce",	--9329
		x"00",	--9330
		x"dc",	--9331
		x"0b",	--9332
		x"6d",	--9333
		x"6d",	--9334
		x"12",	--9335
		x"6c",	--9336
		x"6c",	--9337
		x"0f",	--9338
		x"6d",	--9339
		x"41",	--9340
		x"6c",	--9341
		x"11",	--9342
		x"6d",	--9343
		x"0d",	--9344
		x"6c",	--9345
		x"14",	--9346
		x"5d",	--9347
		x"01",	--9348
		x"5d",	--9349
		x"01",	--9350
		x"14",	--9351
		x"4d",	--9352
		x"09",	--9353
		x"1e",	--9354
		x"0f",	--9355
		x"3b",	--9356
		x"30",	--9357
		x"6c",	--9358
		x"28",	--9359
		x"ce",	--9360
		x"01",	--9361
		x"f7",	--9362
		x"3e",	--9363
		x"0f",	--9364
		x"3b",	--9365
		x"30",	--9366
		x"cf",	--9367
		x"01",	--9368
		x"f0",	--9369
		x"3e",	--9370
		x"f8",	--9371
		x"1b",	--9372
		x"02",	--9373
		x"1c",	--9374
		x"02",	--9375
		x"0c",	--9376
		x"e6",	--9377
		x"0b",	--9378
		x"16",	--9379
		x"1b",	--9380
		x"04",	--9381
		x"1f",	--9382
		x"06",	--9383
		x"1c",	--9384
		x"04",	--9385
		x"1e",	--9386
		x"06",	--9387
		x"0e",	--9388
		x"da",	--9389
		x"0f",	--9390
		x"02",	--9391
		x"0c",	--9392
		x"d6",	--9393
		x"0f",	--9394
		x"06",	--9395
		x"0e",	--9396
		x"02",	--9397
		x"0b",	--9398
		x"02",	--9399
		x"0e",	--9400
		x"d1",	--9401
		x"4d",	--9402
		x"ce",	--9403
		x"3e",	--9404
		x"d6",	--9405
		x"6c",	--9406
		x"d7",	--9407
		x"5e",	--9408
		x"01",	--9409
		x"5f",	--9410
		x"01",	--9411
		x"0e",	--9412
		x"c5",	--9413
		x"1e",	--9414
		x"4a",	--9415
		x"1e",	--9416
		x"0b",	--9417
		x"1d",	--9418
		x"48",	--9419
		x"cd",	--9420
		x"00",	--9421
		x"1d",	--9422
		x"82",	--9423
		x"48",	--9424
		x"3e",	--9425
		x"82",	--9426
		x"4a",	--9427
		x"30",	--9428
		x"3f",	--9429
		x"30",	--9430
		x"0b",	--9431
		x"0a",	--9432
		x"21",	--9433
		x"81",	--9434
		x"00",	--9435
		x"1a",	--9436
		x"48",	--9437
		x"1b",	--9438
		x"4a",	--9439
		x"0d",	--9440
		x"0e",	--9441
		x"3f",	--9442
		x"8c",	--9443
		x"b0",	--9444
		x"e0",	--9445
		x"0f",	--9446
		x"05",	--9447
		x"0e",	--9448
		x"0e",	--9449
		x"ce",	--9450
		x"ff",	--9451
		x"04",	--9452
		x"1e",	--9453
		x"48",	--9454
		x"ce",	--9455
		x"00",	--9456
		x"21",	--9457
		x"3a",	--9458
		x"3b",	--9459
		x"30",	--9460
		x"92",	--9461
		x"02",	--9462
		x"48",	--9463
		x"b2",	--9464
		x"ff",	--9465
		x"4a",	--9466
		x"0e",	--9467
		x"3e",	--9468
		x"06",	--9469
		x"1f",	--9470
		x"04",	--9471
		x"b0",	--9472
		x"ae",	--9473
		x"30",	--9474
		x"92",	--9475
		x"02",	--9476
		x"48",	--9477
		x"92",	--9478
		x"04",	--9479
		x"4a",	--9480
		x"0e",	--9481
		x"3e",	--9482
		x"1f",	--9483
		x"06",	--9484
		x"b0",	--9485
		x"ae",	--9486
		x"30",	--9487
		x"0c",	--9488
		x"82",	--9489
		x"48",	--9490
		x"b2",	--9491
		x"ff",	--9492
		x"4a",	--9493
		x"0e",	--9494
		x"0f",	--9495
		x"b0",	--9496
		x"ae",	--9497
		x"30",	--9498
		x"82",	--9499
		x"48",	--9500
		x"82",	--9501
		x"4a",	--9502
		x"0e",	--9503
		x"0f",	--9504
		x"b0",	--9505
		x"ae",	--9506
		x"30",	--9507
		x"0b",	--9508
		x"0a",	--9509
		x"09",	--9510
		x"08",	--9511
		x"07",	--9512
		x"06",	--9513
		x"05",	--9514
		x"04",	--9515
		x"31",	--9516
		x"08",	--9517
		x"81",	--9518
		x"04",	--9519
		x"09",	--9520
		x"1f",	--9521
		x"1a",	--9522
		x"1d",	--9523
		x"1c",	--9524
		x"4c",	--9525
		x"04",	--9526
		x"84",	--9527
		x"45",	--9528
		x"4e",	--9529
		x"7e",	--9530
		x"40",	--9531
		x"11",	--9532
		x"f1",	--9533
		x"30",	--9534
		x"00",	--9535
		x"0e",	--9536
		x"8e",	--9537
		x"5e",	--9538
		x"03",	--9539
		x"7e",	--9540
		x"58",	--9541
		x"02",	--9542
		x"7e",	--9543
		x"78",	--9544
		x"c1",	--9545
		x"01",	--9546
		x"0c",	--9547
		x"2c",	--9548
		x"0f",	--9549
		x"7e",	--9550
		x"20",	--9551
		x"04",	--9552
		x"f1",	--9553
		x"30",	--9554
		x"00",	--9555
		x"04",	--9556
		x"4c",	--9557
		x"05",	--9558
		x"c1",	--9559
		x"00",	--9560
		x"0c",	--9561
		x"1c",	--9562
		x"01",	--9563
		x"0c",	--9564
		x"0a",	--9565
		x"8c",	--9566
		x"8c",	--9567
		x"8c",	--9568
		x"8c",	--9569
		x"0b",	--9570
		x"06",	--9571
		x"0c",	--9572
		x"8c",	--9573
		x"8c",	--9574
		x"8c",	--9575
		x"8c",	--9576
		x"07",	--9577
		x"0a",	--9578
		x"0b",	--9579
		x"0e",	--9580
		x"8e",	--9581
		x"c1",	--9582
		x"02",	--9583
		x"6e",	--9584
		x"02",	--9585
		x"07",	--9586
		x"01",	--9587
		x"37",	--9588
		x"4f",	--9589
		x"7f",	--9590
		x"10",	--9591
		x"3c",	--9592
		x"1d",	--9593
		x"04",	--9594
		x"3d",	--9595
		x"1d",	--9596
		x"cd",	--9597
		x"00",	--9598
		x"fc",	--9599
		x"1d",	--9600
		x"04",	--9601
		x"09",	--9602
		x"02",	--9603
		x"09",	--9604
		x"01",	--9605
		x"09",	--9606
		x"e1",	--9607
		x"02",	--9608
		x"05",	--9609
		x"09",	--9610
		x"02",	--9611
		x"09",	--9612
		x"01",	--9613
		x"09",	--9614
		x"05",	--9615
		x"07",	--9616
		x"01",	--9617
		x"05",	--9618
		x"4f",	--9619
		x"0d",	--9620
		x"f1",	--9621
		x"20",	--9622
		x"06",	--9623
		x"06",	--9624
		x"0b",	--9625
		x"0e",	--9626
		x"0f",	--9627
		x"0f",	--9628
		x"6f",	--9629
		x"8f",	--9630
		x"16",	--9631
		x"88",	--9632
		x"01",	--9633
		x"06",	--9634
		x"06",	--9635
		x"f6",	--9636
		x"0b",	--9637
		x"f1",	--9638
		x"30",	--9639
		x"06",	--9640
		x"05",	--9641
		x"05",	--9642
		x"5f",	--9643
		x"06",	--9644
		x"8f",	--9645
		x"88",	--9646
		x"1b",	--9647
		x"0f",	--9648
		x"0f",	--9649
		x"0f",	--9650
		x"f7",	--9651
		x"0a",	--9652
		x"06",	--9653
		x"0b",	--9654
		x"07",	--9655
		x"1b",	--9656
		x"0f",	--9657
		x"0f",	--9658
		x"6f",	--9659
		x"8f",	--9660
		x"16",	--9661
		x"88",	--9662
		x"06",	--9663
		x"f7",	--9664
		x"e1",	--9665
		x"02",	--9666
		x"02",	--9667
		x"4a",	--9668
		x"08",	--9669
		x"1a",	--9670
		x"04",	--9671
		x"0a",	--9672
		x"0d",	--9673
		x"3f",	--9674
		x"30",	--9675
		x"88",	--9676
		x"7a",	--9677
		x"4a",	--9678
		x"fa",	--9679
		x"44",	--9680
		x"0b",	--9681
		x"f3",	--9682
		x"37",	--9683
		x"8f",	--9684
		x"88",	--9685
		x"1b",	--9686
		x"0f",	--9687
		x"0f",	--9688
		x"6f",	--9689
		x"4f",	--9690
		x"07",	--9691
		x"07",	--9692
		x"f5",	--9693
		x"04",	--9694
		x"3f",	--9695
		x"20",	--9696
		x"88",	--9697
		x"1b",	--9698
		x"0b",	--9699
		x"fa",	--9700
		x"0f",	--9701
		x"31",	--9702
		x"34",	--9703
		x"35",	--9704
		x"36",	--9705
		x"37",	--9706
		x"38",	--9707
		x"39",	--9708
		x"3a",	--9709
		x"3b",	--9710
		x"30",	--9711
		x"0b",	--9712
		x"0a",	--9713
		x"09",	--9714
		x"08",	--9715
		x"07",	--9716
		x"06",	--9717
		x"05",	--9718
		x"04",	--9719
		x"31",	--9720
		x"b6",	--9721
		x"81",	--9722
		x"3a",	--9723
		x"06",	--9724
		x"05",	--9725
		x"81",	--9726
		x"3e",	--9727
		x"c1",	--9728
		x"2f",	--9729
		x"c1",	--9730
		x"2b",	--9731
		x"c1",	--9732
		x"2e",	--9733
		x"c1",	--9734
		x"2a",	--9735
		x"81",	--9736
		x"30",	--9737
		x"81",	--9738
		x"26",	--9739
		x"07",	--9740
		x"81",	--9741
		x"2c",	--9742
		x"0e",	--9743
		x"3e",	--9744
		x"1c",	--9745
		x"81",	--9746
		x"1c",	--9747
		x"30",	--9748
		x"5a",	--9749
		x"0f",	--9750
		x"1f",	--9751
		x"81",	--9752
		x"40",	--9753
		x"07",	--9754
		x"1e",	--9755
		x"7e",	--9756
		x"25",	--9757
		x"13",	--9758
		x"81",	--9759
		x"00",	--9760
		x"81",	--9761
		x"02",	--9762
		x"81",	--9763
		x"3e",	--9764
		x"c1",	--9765
		x"2f",	--9766
		x"c1",	--9767
		x"2b",	--9768
		x"c1",	--9769
		x"2e",	--9770
		x"c1",	--9771
		x"2a",	--9772
		x"81",	--9773
		x"30",	--9774
		x"30",	--9775
		x"50",	--9776
		x"05",	--9777
		x"8e",	--9778
		x"0f",	--9779
		x"91",	--9780
		x"3c",	--9781
		x"91",	--9782
		x"2c",	--9783
		x"30",	--9784
		x"36",	--9785
		x"7e",	--9786
		x"63",	--9787
		x"c5",	--9788
		x"7e",	--9789
		x"64",	--9790
		x"27",	--9791
		x"7e",	--9792
		x"30",	--9793
		x"94",	--9794
		x"7e",	--9795
		x"31",	--9796
		x"1a",	--9797
		x"7e",	--9798
		x"2a",	--9799
		x"77",	--9800
		x"7e",	--9801
		x"2b",	--9802
		x"0a",	--9803
		x"7e",	--9804
		x"23",	--9805
		x"42",	--9806
		x"7e",	--9807
		x"25",	--9808
		x"e0",	--9809
		x"7e",	--9810
		x"20",	--9811
		x"32",	--9812
		x"56",	--9813
		x"7e",	--9814
		x"2d",	--9815
		x"49",	--9816
		x"7e",	--9817
		x"2e",	--9818
		x"5b",	--9819
		x"7e",	--9820
		x"2b",	--9821
		x"28",	--9822
		x"47",	--9823
		x"7e",	--9824
		x"3a",	--9825
		x"8c",	--9826
		x"7e",	--9827
		x"58",	--9828
		x"21",	--9829
		x"e9",	--9830
		x"7e",	--9831
		x"6f",	--9832
		x"24",	--9833
		x"7e",	--9834
		x"70",	--9835
		x"0a",	--9836
		x"7e",	--9837
		x"69",	--9838
		x"e3",	--9839
		x"7e",	--9840
		x"6c",	--9841
		x"22",	--9842
		x"7e",	--9843
		x"64",	--9844
		x"11",	--9845
		x"dc",	--9846
		x"7e",	--9847
		x"73",	--9848
		x"98",	--9849
		x"7e",	--9850
		x"74",	--9851
		x"04",	--9852
		x"7e",	--9853
		x"70",	--9854
		x"07",	--9855
		x"b8",	--9856
		x"7e",	--9857
		x"75",	--9858
		x"d1",	--9859
		x"7e",	--9860
		x"78",	--9861
		x"d2",	--9862
		x"19",	--9863
		x"3e",	--9864
		x"18",	--9865
		x"2c",	--9866
		x"08",	--9867
		x"30",	--9868
		x"24",	--9869
		x"b1",	--9870
		x"28",	--9871
		x"cb",	--9872
		x"f1",	--9873
		x"00",	--9874
		x"30",	--9875
		x"54",	--9876
		x"69",	--9877
		x"59",	--9878
		x"6e",	--9879
		x"04",	--9880
		x"7e",	--9881
		x"fe",	--9882
		x"6e",	--9883
		x"01",	--9884
		x"5e",	--9885
		x"c1",	--9886
		x"00",	--9887
		x"30",	--9888
		x"54",	--9889
		x"f1",	--9890
		x"10",	--9891
		x"00",	--9892
		x"30",	--9893
		x"54",	--9894
		x"f1",	--9895
		x"2b",	--9896
		x"02",	--9897
		x"30",	--9898
		x"54",	--9899
		x"f1",	--9900
		x"2b",	--9901
		x"02",	--9902
		x"02",	--9903
		x"30",	--9904
		x"54",	--9905
		x"f1",	--9906
		x"20",	--9907
		x"02",	--9908
		x"30",	--9909
		x"54",	--9910
		x"c1",	--9911
		x"2a",	--9912
		x"02",	--9913
		x"30",	--9914
		x"3a",	--9915
		x"d1",	--9916
		x"2e",	--9917
		x"30",	--9918
		x"54",	--9919
		x"0e",	--9920
		x"2e",	--9921
		x"2a",	--9922
		x"0a",	--9923
		x"03",	--9924
		x"81",	--9925
		x"26",	--9926
		x"0d",	--9927
		x"c1",	--9928
		x"2e",	--9929
		x"02",	--9930
		x"30",	--9931
		x"4a",	--9932
		x"f1",	--9933
		x"10",	--9934
		x"00",	--9935
		x"3a",	--9936
		x"81",	--9937
		x"26",	--9938
		x"91",	--9939
		x"26",	--9940
		x"05",	--9941
		x"27",	--9942
		x"81",	--9943
		x"26",	--9944
		x"15",	--9945
		x"c1",	--9946
		x"2e",	--9947
		x"12",	--9948
		x"69",	--9949
		x"79",	--9950
		x"10",	--9951
		x"5e",	--9952
		x"01",	--9953
		x"4e",	--9954
		x"4e",	--9955
		x"0e",	--9956
		x"0e",	--9957
		x"4e",	--9958
		x"6a",	--9959
		x"7a",	--9960
		x"7f",	--9961
		x"4a",	--9962
		x"c1",	--9963
		x"00",	--9964
		x"30",	--9965
		x"54",	--9966
		x"1a",	--9967
		x"26",	--9968
		x"0a",	--9969
		x"0c",	--9970
		x"0c",	--9971
		x"0c",	--9972
		x"0a",	--9973
		x"81",	--9974
		x"26",	--9975
		x"b1",	--9976
		x"d0",	--9977
		x"26",	--9978
		x"8e",	--9979
		x"81",	--9980
		x"26",	--9981
		x"d1",	--9982
		x"2a",	--9983
		x"30",	--9984
		x"54",	--9985
		x"07",	--9986
		x"27",	--9987
		x"6e",	--9988
		x"c1",	--9989
		x"2e",	--9990
		x"03",	--9991
		x"c1",	--9992
		x"2a",	--9993
		x"26",	--9994
		x"c1",	--9995
		x"04",	--9996
		x"c1",	--9997
		x"05",	--9998
		x"0e",	--9999
		x"2e",	--10000
		x"03",	--10001
		x"07",	--10002
		x"27",	--10003
		x"2e",	--10004
		x"c1",	--10005
		x"2e",	--10006
		x"07",	--10007
		x"e1",	--10008
		x"01",	--10009
		x"1f",	--10010
		x"26",	--10011
		x"c1",	--10012
		x"03",	--10013
		x"06",	--10014
		x"c1",	--10015
		x"2a",	--10016
		x"03",	--10017
		x"91",	--10018
		x"26",	--10019
		x"30",	--10020
		x"0e",	--10021
		x"02",	--10022
		x"3e",	--10023
		x"46",	--10024
		x"11",	--10025
		x"04",	--10026
		x"11",	--10027
		x"04",	--10028
		x"1d",	--10029
		x"34",	--10030
		x"1f",	--10031
		x"3e",	--10032
		x"b0",	--10033
		x"48",	--10034
		x"21",	--10035
		x"81",	--10036
		x"2c",	--10037
		x"05",	--10038
		x"30",	--10039
		x"36",	--10040
		x"07",	--10041
		x"27",	--10042
		x"29",	--10043
		x"81",	--10044
		x"1e",	--10045
		x"5e",	--10046
		x"09",	--10047
		x"01",	--10048
		x"4e",	--10049
		x"4e",	--10050
		x"4e",	--10051
		x"4e",	--10052
		x"6a",	--10053
		x"7a",	--10054
		x"f7",	--10055
		x"4a",	--10056
		x"c1",	--10057
		x"00",	--10058
		x"05",	--10059
		x"b1",	--10060
		x"10",	--10061
		x"28",	--10062
		x"53",	--10063
		x"d1",	--10064
		x"01",	--10065
		x"06",	--10066
		x"e1",	--10067
		x"00",	--10068
		x"b1",	--10069
		x"0a",	--10070
		x"28",	--10071
		x"03",	--10072
		x"b1",	--10073
		x"10",	--10074
		x"28",	--10075
		x"6b",	--10076
		x"6b",	--10077
		x"24",	--10078
		x"0c",	--10079
		x"3c",	--10080
		x"28",	--10081
		x"17",	--10082
		x"02",	--10083
		x"16",	--10084
		x"04",	--10085
		x"1b",	--10086
		x"06",	--10087
		x"81",	--10088
		x"1e",	--10089
		x"81",	--10090
		x"20",	--10091
		x"81",	--10092
		x"22",	--10093
		x"81",	--10094
		x"24",	--10095
		x"d1",	--10096
		x"2b",	--10097
		x"08",	--10098
		x"06",	--10099
		x"07",	--10100
		x"04",	--10101
		x"06",	--10102
		x"02",	--10103
		x"0b",	--10104
		x"02",	--10105
		x"c1",	--10106
		x"2b",	--10107
		x"0b",	--10108
		x"0b",	--10109
		x"0b",	--10110
		x"c1",	--10111
		x"2f",	--10112
		x"05",	--10113
		x"20",	--10114
		x"5b",	--10115
		x"07",	--10116
		x"0d",	--10117
		x"27",	--10118
		x"28",	--10119
		x"1b",	--10120
		x"02",	--10121
		x"81",	--10122
		x"1e",	--10123
		x"81",	--10124
		x"20",	--10125
		x"d1",	--10126
		x"2b",	--10127
		x"08",	--10128
		x"09",	--10129
		x"06",	--10130
		x"27",	--10131
		x"2b",	--10132
		x"81",	--10133
		x"1e",	--10134
		x"d1",	--10135
		x"2b",	--10136
		x"0b",	--10137
		x"02",	--10138
		x"c1",	--10139
		x"2b",	--10140
		x"0b",	--10141
		x"0b",	--10142
		x"0b",	--10143
		x"c1",	--10144
		x"2f",	--10145
		x"05",	--10146
		x"f1",	--10147
		x"00",	--10148
		x"12",	--10149
		x"c1",	--10150
		x"2b",	--10151
		x"0f",	--10152
		x"68",	--10153
		x"b1",	--10154
		x"10",	--10155
		x"28",	--10156
		x"03",	--10157
		x"78",	--10158
		x"40",	--10159
		x"05",	--10160
		x"b1",	--10161
		x"28",	--10162
		x"04",	--10163
		x"78",	--10164
		x"20",	--10165
		x"c1",	--10166
		x"00",	--10167
		x"68",	--10168
		x"68",	--10169
		x"30",	--10170
		x"c1",	--10171
		x"2f",	--10172
		x"2d",	--10173
		x"f1",	--10174
		x"2d",	--10175
		x"02",	--10176
		x"68",	--10177
		x"11",	--10178
		x"b1",	--10179
		x"1e",	--10180
		x"b1",	--10181
		x"20",	--10182
		x"b1",	--10183
		x"22",	--10184
		x"b1",	--10185
		x"24",	--10186
		x"91",	--10187
		x"1e",	--10188
		x"81",	--10189
		x"20",	--10190
		x"81",	--10191
		x"22",	--10192
		x"81",	--10193
		x"24",	--10194
		x"17",	--10195
		x"58",	--10196
		x"0f",	--10197
		x"1a",	--10198
		x"1e",	--10199
		x"1b",	--10200
		x"20",	--10201
		x"3a",	--10202
		x"3b",	--10203
		x"0e",	--10204
		x"0f",	--10205
		x"1e",	--10206
		x"0f",	--10207
		x"81",	--10208
		x"1e",	--10209
		x"81",	--10210
		x"20",	--10211
		x"06",	--10212
		x"1a",	--10213
		x"1e",	--10214
		x"3a",	--10215
		x"1a",	--10216
		x"81",	--10217
		x"1e",	--10218
		x"c1",	--10219
		x"1b",	--10220
		x"68",	--10221
		x"6a",	--10222
		x"16",	--10223
		x"1e",	--10224
		x"91",	--10225
		x"20",	--10226
		x"3c",	--10227
		x"18",	--10228
		x"22",	--10229
		x"14",	--10230
		x"24",	--10231
		x"07",	--10232
		x"37",	--10233
		x"1a",	--10234
		x"09",	--10235
		x"91",	--10236
		x"28",	--10237
		x"32",	--10238
		x"1b",	--10239
		x"28",	--10240
		x"8b",	--10241
		x"8b",	--10242
		x"8b",	--10243
		x"8b",	--10244
		x"81",	--10245
		x"34",	--10246
		x"81",	--10247
		x"36",	--10248
		x"81",	--10249
		x"38",	--10250
		x"11",	--10251
		x"3a",	--10252
		x"11",	--10253
		x"3a",	--10254
		x"11",	--10255
		x"3a",	--10256
		x"11",	--10257
		x"3a",	--10258
		x"0c",	--10259
		x"1d",	--10260
		x"44",	--10261
		x"0e",	--10262
		x"0f",	--10263
		x"b0",	--10264
		x"ea",	--10265
		x"31",	--10266
		x"0b",	--10267
		x"3c",	--10268
		x"0a",	--10269
		x"05",	--10270
		x"7b",	--10271
		x"30",	--10272
		x"c7",	--10273
		x"00",	--10274
		x"0c",	--10275
		x"4b",	--10276
		x"d1",	--10277
		x"01",	--10278
		x"03",	--10279
		x"7a",	--10280
		x"37",	--10281
		x"02",	--10282
		x"7a",	--10283
		x"57",	--10284
		x"4a",	--10285
		x"c7",	--10286
		x"00",	--10287
		x"06",	--10288
		x"36",	--10289
		x"11",	--10290
		x"3a",	--10291
		x"11",	--10292
		x"3a",	--10293
		x"11",	--10294
		x"3a",	--10295
		x"11",	--10296
		x"3a",	--10297
		x"0c",	--10298
		x"1d",	--10299
		x"44",	--10300
		x"0e",	--10301
		x"0f",	--10302
		x"b0",	--10303
		x"c4",	--10304
		x"31",	--10305
		x"09",	--10306
		x"81",	--10307
		x"3c",	--10308
		x"08",	--10309
		x"04",	--10310
		x"37",	--10311
		x"0c",	--10312
		x"b2",	--10313
		x"0d",	--10314
		x"b0",	--10315
		x"0e",	--10316
		x"ae",	--10317
		x"0f",	--10318
		x"ac",	--10319
		x"81",	--10320
		x"1e",	--10321
		x"81",	--10322
		x"20",	--10323
		x"81",	--10324
		x"22",	--10325
		x"81",	--10326
		x"24",	--10327
		x"6c",	--10328
		x"58",	--10329
		x"3e",	--10330
		x"14",	--10331
		x"1e",	--10332
		x"17",	--10333
		x"20",	--10334
		x"08",	--10335
		x"38",	--10336
		x"1a",	--10337
		x"19",	--10338
		x"28",	--10339
		x"89",	--10340
		x"89",	--10341
		x"89",	--10342
		x"89",	--10343
		x"1c",	--10344
		x"28",	--10345
		x"0d",	--10346
		x"0e",	--10347
		x"0f",	--10348
		x"b0",	--10349
		x"ee",	--10350
		x"0b",	--10351
		x"3e",	--10352
		x"0a",	--10353
		x"05",	--10354
		x"7b",	--10355
		x"30",	--10356
		x"c8",	--10357
		x"00",	--10358
		x"0c",	--10359
		x"4b",	--10360
		x"d1",	--10361
		x"01",	--10362
		x"03",	--10363
		x"7a",	--10364
		x"37",	--10365
		x"02",	--10366
		x"7a",	--10367
		x"57",	--10368
		x"4a",	--10369
		x"c8",	--10370
		x"00",	--10371
		x"06",	--10372
		x"36",	--10373
		x"1c",	--10374
		x"28",	--10375
		x"0d",	--10376
		x"0e",	--10377
		x"0f",	--10378
		x"b0",	--10379
		x"b8",	--10380
		x"04",	--10381
		x"07",	--10382
		x"38",	--10383
		x"0e",	--10384
		x"d0",	--10385
		x"0f",	--10386
		x"ce",	--10387
		x"81",	--10388
		x"1e",	--10389
		x"81",	--10390
		x"20",	--10391
		x"2c",	--10392
		x"17",	--10393
		x"1e",	--10394
		x"08",	--10395
		x"38",	--10396
		x"1a",	--10397
		x"1e",	--10398
		x"28",	--10399
		x"0f",	--10400
		x"b0",	--10401
		x"5e",	--10402
		x"0d",	--10403
		x"3f",	--10404
		x"0a",	--10405
		x"05",	--10406
		x"7d",	--10407
		x"30",	--10408
		x"c8",	--10409
		x"00",	--10410
		x"0c",	--10411
		x"4d",	--10412
		x"d1",	--10413
		x"01",	--10414
		x"03",	--10415
		x"7c",	--10416
		x"37",	--10417
		x"02",	--10418
		x"7c",	--10419
		x"57",	--10420
		x"4c",	--10421
		x"c8",	--10422
		x"00",	--10423
		x"06",	--10424
		x"36",	--10425
		x"1e",	--10426
		x"28",	--10427
		x"0f",	--10428
		x"b0",	--10429
		x"44",	--10430
		x"07",	--10431
		x"38",	--10432
		x"0f",	--10433
		x"db",	--10434
		x"81",	--10435
		x"1e",	--10436
		x"b1",	--10437
		x"0a",	--10438
		x"28",	--10439
		x"02",	--10440
		x"c1",	--10441
		x"02",	--10442
		x"c1",	--10443
		x"2e",	--10444
		x"2a",	--10445
		x"0f",	--10446
		x"3f",	--10447
		x"1c",	--10448
		x"81",	--10449
		x"42",	--10450
		x"1a",	--10451
		x"1c",	--10452
		x"8a",	--10453
		x"8a",	--10454
		x"8a",	--10455
		x"8a",	--10456
		x"81",	--10457
		x"44",	--10458
		x"81",	--10459
		x"46",	--10460
		x"0a",	--10461
		x"8a",	--10462
		x"8a",	--10463
		x"8a",	--10464
		x"8a",	--10465
		x"81",	--10466
		x"48",	--10467
		x"1c",	--10468
		x"42",	--10469
		x"1d",	--10470
		x"44",	--10471
		x"1c",	--10472
		x"46",	--10473
		x"1d",	--10474
		x"48",	--10475
		x"2c",	--10476
		x"1c",	--10477
		x"26",	--10478
		x"0e",	--10479
		x"e1",	--10480
		x"01",	--10481
		x"5e",	--10482
		x"26",	--10483
		x"4e",	--10484
		x"c1",	--10485
		x"03",	--10486
		x"06",	--10487
		x"c1",	--10488
		x"2a",	--10489
		x"03",	--10490
		x"91",	--10491
		x"26",	--10492
		x"30",	--10493
		x"11",	--10494
		x"04",	--10495
		x"11",	--10496
		x"04",	--10497
		x"1d",	--10498
		x"34",	--10499
		x"0e",	--10500
		x"1e",	--10501
		x"1f",	--10502
		x"3e",	--10503
		x"b0",	--10504
		x"48",	--10505
		x"21",	--10506
		x"81",	--10507
		x"2c",	--10508
		x"0d",	--10509
		x"7f",	--10510
		x"8f",	--10511
		x"91",	--10512
		x"3c",	--10513
		x"0e",	--10514
		x"0e",	--10515
		x"19",	--10516
		x"40",	--10517
		x"f7",	--10518
		x"81",	--10519
		x"3e",	--10520
		x"81",	--10521
		x"2c",	--10522
		x"07",	--10523
		x"0e",	--10524
		x"91",	--10525
		x"26",	--10526
		x"30",	--10527
		x"d1",	--10528
		x"2e",	--10529
		x"c1",	--10530
		x"2a",	--10531
		x"03",	--10532
		x"05",	--10533
		x"d1",	--10534
		x"2a",	--10535
		x"81",	--10536
		x"26",	--10537
		x"17",	--10538
		x"16",	--10539
		x"40",	--10540
		x"6e",	--10541
		x"4e",	--10542
		x"02",	--10543
		x"30",	--10544
		x"2c",	--10545
		x"1f",	--10546
		x"2c",	--10547
		x"31",	--10548
		x"4a",	--10549
		x"34",	--10550
		x"35",	--10551
		x"36",	--10552
		x"37",	--10553
		x"38",	--10554
		x"39",	--10555
		x"3a",	--10556
		x"3b",	--10557
		x"30",	--10558
		x"0d",	--10559
		x"0f",	--10560
		x"04",	--10561
		x"3d",	--10562
		x"03",	--10563
		x"3f",	--10564
		x"1f",	--10565
		x"0e",	--10566
		x"03",	--10567
		x"5d",	--10568
		x"3e",	--10569
		x"1e",	--10570
		x"0d",	--10571
		x"b0",	--10572
		x"44",	--10573
		x"3d",	--10574
		x"6d",	--10575
		x"02",	--10576
		x"3e",	--10577
		x"1e",	--10578
		x"5d",	--10579
		x"02",	--10580
		x"3f",	--10581
		x"1f",	--10582
		x"30",	--10583
		x"b0",	--10584
		x"7e",	--10585
		x"0f",	--10586
		x"30",	--10587
		x"0b",	--10588
		x"0a",	--10589
		x"09",	--10590
		x"79",	--10591
		x"20",	--10592
		x"0a",	--10593
		x"0b",	--10594
		x"0c",	--10595
		x"0d",	--10596
		x"0e",	--10597
		x"0f",	--10598
		x"0c",	--10599
		x"0d",	--10600
		x"0d",	--10601
		x"06",	--10602
		x"02",	--10603
		x"0c",	--10604
		x"03",	--10605
		x"0c",	--10606
		x"0d",	--10607
		x"1e",	--10608
		x"19",	--10609
		x"f2",	--10610
		x"39",	--10611
		x"3a",	--10612
		x"3b",	--10613
		x"30",	--10614
		x"b0",	--10615
		x"b8",	--10616
		x"0e",	--10617
		x"0f",	--10618
		x"30",	--10619
		x"0b",	--10620
		x"0b",	--10621
		x"0f",	--10622
		x"06",	--10623
		x"3b",	--10624
		x"03",	--10625
		x"3e",	--10626
		x"3f",	--10627
		x"1e",	--10628
		x"0f",	--10629
		x"0d",	--10630
		x"05",	--10631
		x"5b",	--10632
		x"3c",	--10633
		x"3d",	--10634
		x"1c",	--10635
		x"0d",	--10636
		x"b0",	--10637
		x"b8",	--10638
		x"6b",	--10639
		x"04",	--10640
		x"3c",	--10641
		x"3d",	--10642
		x"1c",	--10643
		x"0d",	--10644
		x"5b",	--10645
		x"04",	--10646
		x"3e",	--10647
		x"3f",	--10648
		x"1e",	--10649
		x"0f",	--10650
		x"3b",	--10651
		x"30",	--10652
		x"b0",	--10653
		x"f8",	--10654
		x"0e",	--10655
		x"0f",	--10656
		x"30",	--10657
		x"7c",	--10658
		x"10",	--10659
		x"0d",	--10660
		x"0e",	--10661
		x"0f",	--10662
		x"0e",	--10663
		x"0e",	--10664
		x"02",	--10665
		x"0e",	--10666
		x"1f",	--10667
		x"1c",	--10668
		x"f8",	--10669
		x"30",	--10670
		x"b0",	--10671
		x"44",	--10672
		x"0f",	--10673
		x"30",	--10674
		x"07",	--10675
		x"06",	--10676
		x"05",	--10677
		x"04",	--10678
		x"30",	--10679
		x"40",	--10680
		x"04",	--10681
		x"05",	--10682
		x"06",	--10683
		x"07",	--10684
		x"08",	--10685
		x"09",	--10686
		x"0a",	--10687
		x"0b",	--10688
		x"0c",	--10689
		x"0d",	--10690
		x"0e",	--10691
		x"0f",	--10692
		x"08",	--10693
		x"09",	--10694
		x"0a",	--10695
		x"0b",	--10696
		x"0b",	--10697
		x"0e",	--10698
		x"08",	--10699
		x"0a",	--10700
		x"0b",	--10701
		x"05",	--10702
		x"09",	--10703
		x"08",	--10704
		x"02",	--10705
		x"08",	--10706
		x"05",	--10707
		x"08",	--10708
		x"09",	--10709
		x"0a",	--10710
		x"0b",	--10711
		x"1c",	--10712
		x"91",	--10713
		x"00",	--10714
		x"e5",	--10715
		x"21",	--10716
		x"34",	--10717
		x"35",	--10718
		x"36",	--10719
		x"37",	--10720
		x"30",	--10721
		x"0b",	--10722
		x"0a",	--10723
		x"09",	--10724
		x"08",	--10725
		x"18",	--10726
		x"0a",	--10727
		x"19",	--10728
		x"0c",	--10729
		x"1a",	--10730
		x"0e",	--10731
		x"1b",	--10732
		x"10",	--10733
		x"b0",	--10734
		x"66",	--10735
		x"38",	--10736
		x"39",	--10737
		x"3a",	--10738
		x"3b",	--10739
		x"30",	--10740
		x"0b",	--10741
		x"0a",	--10742
		x"09",	--10743
		x"08",	--10744
		x"18",	--10745
		x"0a",	--10746
		x"19",	--10747
		x"0c",	--10748
		x"1a",	--10749
		x"0e",	--10750
		x"1b",	--10751
		x"10",	--10752
		x"b0",	--10753
		x"66",	--10754
		x"0c",	--10755
		x"0d",	--10756
		x"0e",	--10757
		x"0f",	--10758
		x"38",	--10759
		x"39",	--10760
		x"3a",	--10761
		x"3b",	--10762
		x"30",	--10763
		x"0b",	--10764
		x"0a",	--10765
		x"09",	--10766
		x"08",	--10767
		x"07",	--10768
		x"18",	--10769
		x"0c",	--10770
		x"19",	--10771
		x"0e",	--10772
		x"1a",	--10773
		x"10",	--10774
		x"1b",	--10775
		x"12",	--10776
		x"b0",	--10777
		x"66",	--10778
		x"17",	--10779
		x"14",	--10780
		x"87",	--10781
		x"00",	--10782
		x"87",	--10783
		x"02",	--10784
		x"87",	--10785
		x"04",	--10786
		x"87",	--10787
		x"06",	--10788
		x"37",	--10789
		x"38",	--10790
		x"39",	--10791
		x"3a",	--10792
		x"3b",	--10793
		x"30",	--10794
		x"00",	--10795
		x"32",	--10796
		x"f0",	--10797
		x"fd",	--10798
		x"7a",	--10799
		x"00",	--10800
		x"64",	--10801
		x"25",	--10802
		x"20",	--10803
		x"64",	--10804
		x"25",	--10805
		x"0d",	--10806
		x"00",	--10807
		x"20",	--10808
		x"25",	--10809
		x"20",	--10810
		x"0d",	--10811
		x"00",	--10812
		x"c2",	--10813
		x"ea",	--10814
		x"f0",	--10815
		x"f8",	--10816
		x"00",	--10817
		x"08",	--10818
		x"da",	--10819
		x"e2",	--10820
		x"0d",	--10821
		x"3d",	--10822
		x"3d",	--10823
		x"3d",	--10824
		x"20",	--10825
		x"61",	--10826
		x"63",	--10827
		x"6c",	--10828
		x"4d",	--10829
		x"55",	--10830
		x"3d",	--10831
		x"3d",	--10832
		x"3d",	--10833
		x"0d",	--10834
		x"00",	--10835
		x"6e",	--10836
		x"65",	--10837
		x"61",	--10838
		x"74",	--10839
		x"76",	--10840
		x"20",	--10841
		x"6f",	--10842
		x"65",	--10843
		x"77",	--10844
		x"69",	--10845
		x"65",	--10846
		x"72",	--10847
		x"61",	--10848
		x"00",	--10849
		x"75",	--10850
		x"7a",	--10851
		x"72",	--10852
		x"70",	--10853
		x"6d",	--10854
		x"65",	--10855
		x"63",	--10856
		x"64",	--10857
		x"72",	--10858
		x"73",	--10859
		x"65",	--10860
		x"64",	--10861
		x"63",	--10862
		x"6e",	--10863
		x"72",	--10864
		x"6c",	--10865
		x"65",	--10866
		x"00",	--10867
		x"64",	--10868
		x"6d",	--10869
		x"74",	--10870
		x"79",	--10871
		x"73",	--10872
		x"65",	--10873
		x"64",	--10874
		x"63",	--10875
		x"6e",	--10876
		x"69",	--10877
		x"75",	--10878
		x"61",	--10879
		x"69",	--10880
		x"6e",	--10881
		x"6f",	--10882
		x"73",	--10883
		x"61",	--10884
		x"6c",	--10885
		x"20",	--10886
		x"76",	--10887
		x"69",	--10888
		x"61",	--10889
		x"63",	--10890
		x"00",	--10891
		x"6f",	--10892
		x"6d",	--10893
		x"62",	--10894
		x"6f",	--10895
		x"6c",	--10896
		x"61",	--10897
		x"65",	--10898
		x"00",	--10899
		x"0a",	--10900
		x"08",	--10901
		x"08",	--10902
		x"25",	--10903
		x"00",	--10904
		x"50",	--10905
		x"0a",	--10906
		x"44",	--10907
		x"57",	--10908
		x"0d",	--10909
		x"00",	--10910
		x"49",	--10911
		x"48",	--10912
		x"0d",	--10913
		x"00",	--10914
		x"45",	--10915
		x"54",	--10916
		x"0a",	--10917
		x"53",	--10918
		x"6f",	--10919
		x"0d",	--10920
		x"00",	--10921
		x"6f",	--10922
		x"72",	--10923
		x"63",	--10924
		x"20",	--10925
		x"73",	--10926
		x"67",	--10927
		x"3a",	--10928
		x"0a",	--10929
		x"09",	--10930
		x"63",	--10931
		x"5b",	--10932
		x"5d",	--10933
		x"4c",	--10934
		x"46",	--10935
		x"20",	--10936
		x"49",	--10937
		x"48",	--10938
		x"20",	--10939
		x"54",	--10940
		x"4d",	--10941
		x"4f",	--10942
		x"54",	--10943
		x"0d",	--10944
		x"00",	--10945
		x"64",	--10946
		x"25",	--10947
		x"0d",	--10948
		x"00",	--10949
		x"6f",	--10950
		x"20",	--10951
		x"6d",	--10952
		x"6c",	--10953
		x"6d",	--10954
		x"6e",	--10955
		x"65",	--10956
		x"20",	--10957
		x"65",	--10958
		x"0d",	--10959
		x"00",	--10960
		x"61",	--10961
		x"74",	--10962
		x"6e",	--10963
		x"20",	--10964
		x"6f",	--10965
		x"20",	--10966
		x"20",	--10967
		x"65",	--10968
		x"20",	--10969
		x"62",	--10970
		x"6e",	--10971
		x"66",	--10972
		x"6c",	--10973
		x"0d",	--10974
		x"00",	--10975
		x"65",	--10976
		x"73",	--10977
		x"6f",	--10978
		x"6c",	--10979
		x"20",	--10980
		x"6f",	--10981
		x"20",	--10982
		x"65",	--10983
		x"20",	--10984
		x"68",	--10985
		x"74",	--10986
		x"0a",	--10987
		x"25",	--10988
		x"20",	--10989
		x"73",	--10990
		x"6e",	--10991
		x"74",	--10992
		x"61",	--10993
		x"6e",	--10994
		x"6d",	--10995
		x"65",	--10996
		x"0d",	--10997
		x"00",	--10998
		x"74",	--10999
		x"70",	--11000
		x"0a",	--11001
		x"65",	--11002
		x"72",	--11003
		x"72",	--11004
		x"20",	--11005
		x"69",	--11006
		x"73",	--11007
		x"6e",	--11008
		x"20",	--11009
		x"72",	--11010
		x"75",	--11011
		x"65",	--11012
		x"74",	--11013
		x"0a",	--11014
		x"63",	--11015
		x"72",	--11016
		x"65",	--11017
		x"74",	--11018
		x"75",	--11019
		x"61",	--11020
		x"65",	--11021
		x"0d",	--11022
		x"00",	--11023
		x"25",	--11024
		x"20",	--11025
		x"45",	--11026
		x"54",	--11027
		x"52",	--11028
		x"47",	--11029
		x"54",	--11030
		x"3c",	--11031
		x"49",	--11032
		x"45",	--11033
		x"55",	--11034
		x"3e",	--11035
		x"0a",	--11036
		x"25",	--11037
		x"20",	--11038
		x"64",	--11039
		x"0a",	--11040
		x"25",	--11041
		x"64",	--11042
		x"25",	--11043
		x"64",	--11044
		x"25",	--11045
		x"0d",	--11046
		x"00",	--11047
		x"64",	--11048
		x"25",	--11049
		x"0d",	--11050
		x"00",	--11051
		x"25",	--11052
		x"20",	--11053
		x"0d",	--11054
		x"00",	--11055
		x"6f",	--11056
		x"62",	--11057
		x"68",	--11058
		x"6e",	--11059
		x"20",	--11060
		x"65",	--11061
		x"0a",	--11062
		x"59",	--11063
		x"20",	--11064
		x"6e",	--11065
		x"66",	--11066
		x"6f",	--11067
		x"74",	--11068
		x"0a",	--11069
		x"59",	--11070
		x"20",	--11071
		x"6e",	--11072
		x"74",	--11073
		x"65",	--11074
		x"72",	--11075
		x"67",	--11076
		x"74",	--11077
		x"0a",	--11078
		x"59",	--11079
		x"20",	--11080
		x"6e",	--11081
		x"74",	--11082
		x"65",	--11083
		x"6c",	--11084
		x"66",	--11085
		x"0d",	--11086
		x"00",	--11087
		x"64",	--11088
		x"0a",	--11089
		x"73",	--11090
		x"6f",	--11091
		x"0d",	--11092
		x"00",	--11093
		x"72",	--11094
		x"6e",	--11095
		x"3a",	--11096
		x"6f",	--11097
		x"61",	--11098
		x"69",	--11099
		x"6e",	--11100
		x"0a",	--11101
		x"6c",	--11102
		x"66",	--11103
		x"3a",	--11104
		x"6f",	--11105
		x"61",	--11106
		x"69",	--11107
		x"6e",	--11108
		x"0a",	--11109
		x"72",	--11110
		x"67",	--11111
		x"74",	--11112
		x"72",	--11113
		x"74",	--11114
		x"74",	--11115
		x"6f",	--11116
		x"0d",	--11117
		x"00",	--11118
		x"6f",	--11119
		x"6d",	--11120
		x"6e",	--11121
		x"20",	--11122
		x"63",	--11123
		x"69",	--11124
		x"61",	--11125
		x"65",	--11126
		x"0d",	--11127
		x"00",	--11128
		x"6f",	--11129
		x"6d",	--11130
		x"6e",	--11131
		x"20",	--11132
		x"65",	--11133
		x"63",	--11134
		x"69",	--11135
		x"61",	--11136
		x"65",	--11137
		x"0d",	--11138
		x"00",	--11139
		x"f4",	--11140
		x"f4",	--11141
		x"f4",	--11142
		x"f4",	--11143
		x"00",	--11144
		x"77",	--11145
		x"69",	--11146
		x"65",	--11147
		x"0d",	--11148
		x"65",	--11149
		x"72",	--11150
		x"72",	--11151
		x"20",	--11152
		x"69",	--11153
		x"73",	--11154
		x"6e",	--11155
		x"20",	--11156
		x"72",	--11157
		x"75",	--11158
		x"65",	--11159
		x"74",	--11160
		x"0a",	--11161
		x"63",	--11162
		x"72",	--11163
		x"65",	--11164
		x"74",	--11165
		x"75",	--11166
		x"61",	--11167
		x"65",	--11168
		x"0d",	--11169
		x"00",	--11170
		x"25",	--11171
		x"20",	--11172
		x"45",	--11173
		x"49",	--11174
		x"54",	--11175
		x"52",	--11176
		x"56",	--11177
		x"4c",	--11178
		x"45",	--11179
		x"0a",	--11180
		x"72",	--11181
		x"25",	--11182
		x"20",	--11183
		x"3d",	--11184
		x"64",	--11185
		x"0a",	--11186
		x"09",	--11187
		x"73",	--11188
		x"52",	--11189
		x"47",	--11190
		x"53",	--11191
		x"45",	--11192
		x"0d",	--11193
		x"00",	--11194
		x"65",	--11195
		x"64",	--11196
		x"0d",	--11197
		x"25",	--11198
		x"20",	--11199
		x"73",	--11200
		x"0a",	--11201
		x"25",	--11202
		x"3a",	--11203
		x"6e",	--11204
		x"20",	--11205
		x"75",	--11206
		x"68",	--11207
		x"63",	--11208
		x"6d",	--11209
		x"61",	--11210
		x"64",	--11211
		x"0a",	--11212
		x"28",	--11213
		x"56",	--11214
		x"56",	--11215
		x"56",	--11216
		x"56",	--11217
		x"56",	--11218
		x"56",	--11219
		x"56",	--11220
		x"56",	--11221
		x"56",	--11222
		x"56",	--11223
		x"56",	--11224
		x"56",	--11225
		x"56",	--11226
		x"56",	--11227
		x"56",	--11228
		x"56",	--11229
		x"56",	--11230
		x"56",	--11231
		x"56",	--11232
		x"56",	--11233
		x"56",	--11234
		x"56",	--11235
		x"56",	--11236
		x"56",	--11237
		x"56",	--11238
		x"56",	--11239
		x"56",	--11240
		x"56",	--11241
		x"1a",	--11242
		x"56",	--11243
		x"56",	--11244
		x"56",	--11245
		x"56",	--11246
		x"56",	--11247
		x"56",	--11248
		x"56",	--11249
		x"56",	--11250
		x"56",	--11251
		x"56",	--11252
		x"56",	--11253
		x"56",	--11254
		x"56",	--11255
		x"56",	--11256
		x"56",	--11257
		x"56",	--11258
		x"56",	--11259
		x"56",	--11260
		x"56",	--11261
		x"56",	--11262
		x"56",	--11263
		x"56",	--11264
		x"56",	--11265
		x"56",	--11266
		x"56",	--11267
		x"56",	--11268
		x"56",	--11269
		x"56",	--11270
		x"56",	--11271
		x"56",	--11272
		x"56",	--11273
		x"0c",	--11274
		x"fe",	--11275
		x"f0",	--11276
		x"56",	--11277
		x"56",	--11278
		x"56",	--11279
		x"56",	--11280
		x"56",	--11281
		x"56",	--11282
		x"56",	--11283
		x"d8",	--11284
		x"56",	--11285
		x"c6",	--11286
		x"56",	--11287
		x"56",	--11288
		x"56",	--11289
		x"56",	--11290
		x"aa",	--11291
		x"56",	--11292
		x"56",	--11293
		x"56",	--11294
		x"9c",	--11295
		x"8a",	--11296
		x"30",	--11297
		x"32",	--11298
		x"34",	--11299
		x"36",	--11300
		x"38",	--11301
		x"61",	--11302
		x"63",	--11303
		x"65",	--11304
		x"00",	--11305
		x"38",	--11306
		x"ed",	--11307
		x"da",	--11308
		x"49",	--11309
		x"5e",	--11310
		x"7b",	--11311
		x"da",	--11312
		x"c9",	--11313
		x"69",	--11314
		x"ac",	--11315
		x"68",	--11316
		x"22",	--11317
		x"b4",	--11318
		x"14",	--11319
		x"68",	--11320
		x"a2",	--11321
		x"00",	--11322
		x"c9",	--11323
		x"00",	--11324
		x"49",	--11325
		x"00",	--11326
		x"96",	--11327
		x"00",	--11328
		x"c9",	--11329
		x"00",	--11330
		x"fb",	--11331
		x"00",	--11332
		x"16",	--11333
		x"00",	--11334
		x"2f",	--11335
		x"00",	--11336
		x"49",	--11337
		x"00",	--11338
		x"62",	--11339
		x"00",	--11340
		x"7b",	--11341
		x"00",	--11342
		x"8a",	--11343
		x"00",	--11344
		x"96",	--11345
		x"00",	--11346
		x"a3",	--11347
		x"00",	--11348
		x"af",	--11349
		x"00",	--11350
		x"bc",	--11351
		x"00",	--11352
		x"c9",	--11353
		x"00",	--11354
		x"d5",	--11355
		x"00",	--11356
		x"e2",	--11357
		x"00",	--11358
		x"ee",	--11359
		x"00",	--11360
		x"fb",	--11361
		x"00",	--11362
		x"03",	--11363
		x"00",	--11364
		x"0a",	--11365
		x"00",	--11366
		x"10",	--11367
		x"00",	--11368
		x"16",	--11369
		x"00",	--11370
		x"1d",	--11371
		x"00",	--11372
		x"23",	--11373
		x"00",	--11374
		x"29",	--11375
		x"00",	--11376
		x"2f",	--11377
		x"00",	--11378
		x"36",	--11379
		x"00",	--11380
		x"3c",	--11381
		x"00",	--11382
		x"42",	--11383
		x"00",	--11384
		x"49",	--11385
		x"a2",	--11386
		x"00",	--11387
		x"f9",	--11388
		x"00",	--11389
		x"83",	--11390
		x"00",	--11391
		x"6e",	--11392
		x"00",	--11393
		x"4e",	--11394
		x"00",	--11395
		x"44",	--11396
		x"00",	--11397
		x"15",	--11398
		x"00",	--11399
		x"29",	--11400
		x"00",	--11401
		x"fc",	--11402
		x"00",	--11403
		x"27",	--11404
		x"00",	--11405
		x"57",	--11406
		x"00",	--11407
		x"d1",	--11408
		x"00",	--11409
		x"f5",	--11410
		x"00",	--11411
		x"34",	--11412
		x"00",	--11413
		x"dd",	--11414
		x"00",	--11415
		x"c0",	--11416
		x"00",	--11417
		x"db",	--11418
		x"00",	--11419
		x"62",	--11420
		x"00",	--11421
		x"95",	--11422
		x"00",	--11423
		x"99",	--11424
		x"00",	--11425
		x"3c",	--11426
		x"00",	--11427
		x"43",	--11428
		x"00",	--11429
		x"90",	--11430
		x"00",	--11431
		x"41",	--11432
		x"00",	--11433
		x"fe",	--11434
		x"00",	--11435
		x"51",	--11436
		x"00",	--11437
		x"63",	--11438
		x"00",	--11439
		x"ab",	--11440
		x"00",	--11441
		x"de",	--11442
		x"00",	--11443
		x"bb",	--11444
		x"00",	--11445
		x"c5",	--11446
		x"00",	--11447
		x"61",	--11448
		x"00",	--11449
		x"b7",	--11450
		x"00",	--11451
		x"24",	--11452
		x"00",	--11453
		x"6e",	--11454
		x"00",	--11455
		x"3a",	--11456
		x"00",	--11457
		x"42",	--11458
		x"00",	--11459
		x"4d",	--11460
		x"00",	--11461
		x"d2",	--11462
		x"00",	--11463
		x"e0",	--11464
		x"00",	--11465
		x"06",	--11466
		x"00",	--11467
		x"49",	--11468
		x"00",	--11469
		x"2e",	--11470
		x"00",	--11471
		x"ea",	--11472
		x"00",	--11473
		x"09",	--11474
		x"00",	--11475
		x"d1",	--11476
		x"00",	--11477
		x"92",	--11478
		x"00",	--11479
		x"1c",	--11480
		x"00",	--11481
		x"fe",	--11482
		x"00",	--11483
		x"1d",	--11484
		x"00",	--11485
		x"eb",	--11486
		x"00",	--11487
		x"1c",	--11488
		x"00",	--11489
		x"b1",	--11490
		x"00",	--11491
		x"29",	--11492
		x"00",	--11493
		x"a7",	--11494
		x"00",	--11495
		x"3e",	--11496
		x"00",	--11497
		x"e8",	--11498
		x"00",	--11499
		x"82",	--11500
		x"00",	--11501
		x"35",	--11502
		x"00",	--11503
		x"f5",	--11504
		x"00",	--11505
		x"2e",	--11506
		x"00",	--11507
		x"bb",	--11508
		x"00",	--11509
		x"44",	--11510
		x"00",	--11511
		x"84",	--11512
		x"00",	--11513
		x"e9",	--11514
		x"00",	--11515
		x"9c",	--11516
		x"00",	--11517
		x"70",	--11518
		x"00",	--11519
		x"26",	--11520
		x"00",	--11521
		x"b4",	--11522
		x"00",	--11523
		x"5f",	--11524
		x"00",	--11525
		x"7e",	--11526
		x"00",	--11527
		x"41",	--11528
		x"00",	--11529
		x"39",	--11530
		x"00",	--11531
		x"91",	--11532
		x"00",	--11533
		x"d6",	--11534
		x"00",	--11535
		x"39",	--11536
		x"00",	--11537
		x"83",	--11538
		x"00",	--11539
		x"53",	--11540
		x"00",	--11541
		x"39",	--11542
		x"00",	--11543
		x"f4",	--11544
		x"00",	--11545
		x"9c",	--11546
		x"00",	--11547
		x"84",	--11548
		x"00",	--11549
		x"5f",	--11550
		x"00",	--11551
		x"8b",	--11552
		x"00",	--11553
		x"bd",	--11554
		x"00",	--11555
		x"f9",	--11556
		x"00",	--11557
		x"28",	--11558
		x"00",	--11559
		x"3b",	--11560
		x"00",	--11561
		x"1f",	--11562
		x"00",	--11563
		x"f8",	--11564
		x"00",	--11565
		x"97",	--11566
		x"00",	--11567
		x"ff",	--11568
		x"00",	--11569
		x"de",	--11570
		x"00",	--11571
		x"05",	--11572
		x"00",	--11573
		x"98",	--11574
		x"00",	--11575
		x"0f",	--11576
		x"00",	--11577
		x"ef",	--11578
		x"00",	--11579
		x"2f",	--11580
		x"00",	--11581
		x"11",	--11582
		x"00",	--11583
		x"8b",	--11584
		x"00",	--11585
		x"5a",	--11586
		x"00",	--11587
		x"0a",	--11588
		x"00",	--11589
		x"6d",	--11590
		x"00",	--11591
		x"1f",	--11592
		x"00",	--11593
		x"6d",	--11594
		x"00",	--11595
		x"36",	--11596
		x"00",	--11597
		x"7e",	--11598
		x"00",	--11599
		x"cf",	--11600
		x"00",	--11601
		x"27",	--11602
		x"00",	--11603
		x"cb",	--11604
		x"00",	--11605
		x"09",	--11606
		x"00",	--11607
		x"b7",	--11608
		x"00",	--11609
		x"4f",	--11610
		x"00",	--11611
		x"46",	--11612
		x"00",	--11613
		x"3f",	--11614
		x"00",	--11615
		x"66",	--11616
		x"00",	--11617
		x"9e",	--11618
		x"00",	--11619
		x"5f",	--11620
		x"00",	--11621
		x"ea",	--11622
		x"00",	--11623
		x"2d",	--11624
		x"00",	--11625
		x"75",	--11626
		x"00",	--11627
		x"27",	--11628
		x"00",	--11629
		x"ba",	--11630
		x"00",	--11631
		x"c7",	--11632
		x"00",	--11633
		x"eb",	--11634
		x"00",	--11635
		x"e5",	--11636
		x"00",	--11637
		x"f1",	--11638
		x"00",	--11639
		x"7b",	--11640
		x"00",	--11641
		x"3d",	--11642
		x"00",	--11643
		x"07",	--11644
		x"00",	--11645
		x"39",	--11646
		x"00",	--11647
		x"f7",	--11648
		x"00",	--11649
		x"8a",	--11650
		x"00",	--11651
		x"52",	--11652
		x"00",	--11653
		x"92",	--11654
		x"00",	--11655
		x"ea",	--11656
		x"00",	--11657
		x"6b",	--11658
		x"00",	--11659
		x"fb",	--11660
		x"00",	--11661
		x"5f",	--11662
		x"00",	--11663
		x"b1",	--11664
		x"00",	--11665
		x"1f",	--11666
		x"00",	--11667
		x"8d",	--11668
		x"00",	--11669
		x"5d",	--11670
		x"00",	--11671
		x"08",	--11672
		x"00",	--11673
		x"56",	--11674
		x"00",	--11675
		x"03",	--11676
		x"00",	--11677
		x"30",	--11678
		x"00",	--11679
		x"46",	--11680
		x"00",	--11681
		x"fc",	--11682
		x"00",	--11683
		x"7b",	--11684
		x"00",	--11685
		x"6b",	--11686
		x"00",	--11687
		x"ab",	--11688
		x"00",	--11689
		x"f0",	--11690
		x"00",	--11691
		x"cf",	--11692
		x"00",	--11693
		x"bc",	--11694
		x"00",	--11695
		x"20",	--11696
		x"00",	--11697
		x"9a",	--11698
		x"00",	--11699
		x"f4",	--11700
		x"00",	--11701
		x"36",	--11702
		x"00",	--11703
		x"1d",	--11704
		x"00",	--11705
		x"a9",	--11706
		x"00",	--11707
		x"e3",	--11708
		x"00",	--11709
		x"91",	--11710
		x"00",	--11711
		x"61",	--11712
		x"00",	--11713
		x"5e",	--11714
		x"00",	--11715
		x"e6",	--11716
		x"00",	--11717
		x"1b",	--11718
		x"00",	--11719
		x"08",	--11720
		x"00",	--11721
		x"65",	--11722
		x"00",	--11723
		x"99",	--11724
		x"00",	--11725
		x"85",	--11726
		x"00",	--11727
		x"5f",	--11728
		x"00",	--11729
		x"14",	--11730
		x"00",	--11731
		x"a0",	--11732
		x"00",	--11733
		x"68",	--11734
		x"00",	--11735
		x"40",	--11736
		x"00",	--11737
		x"8d",	--11738
		x"00",	--11739
		x"ff",	--11740
		x"00",	--11741
		x"d8",	--11742
		x"00",	--11743
		x"80",	--11744
		x"00",	--11745
		x"4d",	--11746
		x"00",	--11747
		x"73",	--11748
		x"00",	--11749
		x"27",	--11750
		x"00",	--11751
		x"31",	--11752
		x"00",	--11753
		x"06",	--11754
		x"00",	--11755
		x"06",	--11756
		x"00",	--11757
		x"15",	--11758
		x"00",	--11759
		x"56",	--11760
		x"00",	--11761
		x"ca",	--11762
		x"00",	--11763
		x"73",	--11764
		x"00",	--11765
		x"a8",	--11766
		x"00",	--11767
		x"c9",	--11768
		x"00",	--11769
		x"60",	--11770
		x"00",	--11771
		x"e2",	--11772
		x"00",	--11773
		x"7b",	--11774
		x"00",	--11775
		x"c0",	--11776
		x"00",	--11777
		x"8c",	--11778
		x"00",	--11779
		x"6b",	--11780
		x"00",	--11781
		x"04",	--11782
		x"07",	--11783
		x"09",	--11784
		x"00",	--11785
		x"c9",	--11786
		x"00",	--11787
		x"f0",	--11788
		x"00",	--11789
		x"da",	--11790
		x"00",	--11791
		x"a2",	--11792
		x"00",	--11793
		x"84",	--11794
		x"00",	--11795
		x"50",	--11796
		x"00",	--11797
		x"c2",	--11798
		x"00",	--11799
		x"d0",	--11800
		x"00",	--11801
		x"c4",	--11802
		x"00",	--11803
		x"c6",	--11804
		x"00",	--11805
		x"44",	--11806
		x"00",	--11807
		x"00",	--11808
		x"00",	--11809
		x"00",	--11810
		x"00",	--11811
		x"02",	--11812
		x"03",	--11813
		x"03",	--11814
		x"04",	--11815
		x"04",	--11816
		x"04",	--11817
		x"04",	--11818
		x"05",	--11819
		x"05",	--11820
		x"05",	--11821
		x"05",	--11822
		x"05",	--11823
		x"05",	--11824
		x"05",	--11825
		x"05",	--11826
		x"06",	--11827
		x"06",	--11828
		x"06",	--11829
		x"06",	--11830
		x"06",	--11831
		x"06",	--11832
		x"06",	--11833
		x"06",	--11834
		x"06",	--11835
		x"06",	--11836
		x"06",	--11837
		x"06",	--11838
		x"06",	--11839
		x"06",	--11840
		x"06",	--11841
		x"06",	--11842
		x"07",	--11843
		x"07",	--11844
		x"07",	--11845
		x"07",	--11846
		x"07",	--11847
		x"07",	--11848
		x"07",	--11849
		x"07",	--11850
		x"07",	--11851
		x"07",	--11852
		x"07",	--11853
		x"07",	--11854
		x"07",	--11855
		x"07",	--11856
		x"07",	--11857
		x"07",	--11858
		x"07",	--11859
		x"07",	--11860
		x"07",	--11861
		x"07",	--11862
		x"07",	--11863
		x"07",	--11864
		x"07",	--11865
		x"07",	--11866
		x"07",	--11867
		x"07",	--11868
		x"07",	--11869
		x"07",	--11870
		x"07",	--11871
		x"07",	--11872
		x"07",	--11873
		x"07",	--11874
		x"08",	--11875
		x"08",	--11876
		x"08",	--11877
		x"08",	--11878
		x"08",	--11879
		x"08",	--11880
		x"08",	--11881
		x"08",	--11882
		x"08",	--11883
		x"08",	--11884
		x"08",	--11885
		x"08",	--11886
		x"08",	--11887
		x"08",	--11888
		x"08",	--11889
		x"08",	--11890
		x"08",	--11891
		x"08",	--11892
		x"08",	--11893
		x"08",	--11894
		x"08",	--11895
		x"08",	--11896
		x"08",	--11897
		x"08",	--11898
		x"08",	--11899
		x"08",	--11900
		x"08",	--11901
		x"08",	--11902
		x"08",	--11903
		x"08",	--11904
		x"08",	--11905
		x"08",	--11906
		x"08",	--11907
		x"08",	--11908
		x"08",	--11909
		x"08",	--11910
		x"08",	--11911
		x"08",	--11912
		x"08",	--11913
		x"08",	--11914
		x"08",	--11915
		x"08",	--11916
		x"08",	--11917
		x"08",	--11918
		x"08",	--11919
		x"08",	--11920
		x"08",	--11921
		x"08",	--11922
		x"08",	--11923
		x"08",	--11924
		x"08",	--11925
		x"08",	--11926
		x"08",	--11927
		x"08",	--11928
		x"08",	--11929
		x"08",	--11930
		x"08",	--11931
		x"08",	--11932
		x"08",	--11933
		x"08",	--11934
		x"08",	--11935
		x"08",	--11936
		x"08",	--11937
		x"08",	--11938
		x"28",	--11939
		x"75",	--11940
		x"6c",	--11941
		x"00",	--11942
		x"ff",	--11943
		x"ff",	--11944
		x"ff",	--11945
		x"ff",	--11946
		x"68",	--11947
		x"6c",	--11948
		x"00",	--11949
		x"ff",	--11950
		x"ff",	--11951
		x"ff",	--11952
		x"ff",	--11953
		x"ff",	--11954
		x"ff",	--11955
		x"ff",	--11956
		x"ff",	--11957
		x"ff",	--11958
		x"ff",	--11959
		x"ff",	--11960
		x"ff",	--11961
		x"ff",	--11962
		x"ff",	--11963
		x"ff",	--11964
		x"ff",	--11965
		x"ff",	--11966
		x"ff",	--11967
		x"ff",	--11968
		x"ff",	--11969
		x"ff",	--11970
		x"ff",	--11971
		x"ff",	--11972
		x"ff",	--11973
		x"ff",	--11974
		x"ff",	--11975
		x"ff",	--11976
		x"ff",	--11977
		x"ff",	--11978
		x"ff",	--11979
		x"ff",	--11980
		x"ff",	--11981
		x"ff",	--11982
		x"ff",	--11983
		x"ff",	--11984
		x"ff",	--11985
		x"ff",	--11986
		x"ff",	--11987
		x"ff",	--11988
		x"ff",	--11989
		x"ff",	--11990
		x"ff",	--11991
		x"ff",	--11992
		x"ff",	--11993
		x"ff",	--11994
		x"ff",	--11995
		x"ff",	--11996
		x"ff",	--11997
		x"ff",	--11998
		x"ff",	--11999
		x"ff",	--12000
		x"ff",	--12001
		x"ff",	--12002
		x"ff",	--12003
		x"ff",	--12004
		x"ff",	--12005
		x"ff",	--12006
		x"ff",	--12007
		x"ff",	--12008
		x"ff",	--12009
		x"ff",	--12010
		x"ff",	--12011
		x"ff",	--12012
		x"ff",	--12013
		x"ff",	--12014
		x"ff",	--12015
		x"ff",	--12016
		x"ff",	--12017
		x"ff",	--12018
		x"ff",	--12019
		x"ff",	--12020
		x"ff",	--12021
		x"ff",	--12022
		x"ff",	--12023
		x"ff",	--12024
		x"ff",	--12025
		x"ff",	--12026
		x"ff",	--12027
		x"ff",	--12028
		x"ff",	--12029
		x"ff",	--12030
		x"ff",	--12031
		x"ff",	--12032
		x"ff",	--12033
		x"ff",	--12034
		x"ff",	--12035
		x"ff",	--12036
		x"ff",	--12037
		x"ff",	--12038
		x"ff",	--12039
		x"ff",	--12040
		x"ff",	--12041
		x"ff",	--12042
		x"ff",	--12043
		x"ff",	--12044
		x"ff",	--12045
		x"ff",	--12046
		x"ff",	--12047
		x"ff",	--12048
		x"ff",	--12049
		x"ff",	--12050
		x"ff",	--12051
		x"ff",	--12052
		x"ff",	--12053
		x"ff",	--12054
		x"ff",	--12055
		x"ff",	--12056
		x"ff",	--12057
		x"ff",	--12058
		x"ff",	--12059
		x"ff",	--12060
		x"ff",	--12061
		x"ff",	--12062
		x"ff",	--12063
		x"ff",	--12064
		x"ff",	--12065
		x"ff",	--12066
		x"ff",	--12067
		x"ff",	--12068
		x"ff",	--12069
		x"ff",	--12070
		x"ff",	--12071
		x"ff",	--12072
		x"ff",	--12073
		x"ff",	--12074
		x"ff",	--12075
		x"ff",	--12076
		x"ff",	--12077
		x"ff",	--12078
		x"ff",	--12079
		x"ff",	--12080
		x"ff",	--12081
		x"ff",	--12082
		x"ff",	--12083
		x"ff",	--12084
		x"ff",	--12085
		x"ff",	--12086
		x"ff",	--12087
		x"ff",	--12088
		x"ff",	--12089
		x"ff",	--12090
		x"ff",	--12091
		x"ff",	--12092
		x"ff",	--12093
		x"ff",	--12094
		x"ff",	--12095
		x"ff",	--12096
		x"ff",	--12097
		x"ff",	--12098
		x"ff",	--12099
		x"ff",	--12100
		x"ff",	--12101
		x"ff",	--12102
		x"ff",	--12103
		x"ff",	--12104
		x"ff",	--12105
		x"ff",	--12106
		x"ff",	--12107
		x"ff",	--12108
		x"ff",	--12109
		x"ff",	--12110
		x"ff",	--12111
		x"ff",	--12112
		x"ff",	--12113
		x"ff",	--12114
		x"ff",	--12115
		x"ff",	--12116
		x"ff",	--12117
		x"ff",	--12118
		x"ff",	--12119
		x"ff",	--12120
		x"ff",	--12121
		x"ff",	--12122
		x"ff",	--12123
		x"ff",	--12124
		x"ff",	--12125
		x"ff",	--12126
		x"ff",	--12127
		x"ff",	--12128
		x"ff",	--12129
		x"ff",	--12130
		x"ff",	--12131
		x"ff",	--12132
		x"ff",	--12133
		x"ff",	--12134
		x"ff",	--12135
		x"ff",	--12136
		x"ff",	--12137
		x"ff",	--12138
		x"ff",	--12139
		x"ff",	--12140
		x"ff",	--12141
		x"ff",	--12142
		x"ff",	--12143
		x"ff",	--12144
		x"ff",	--12145
		x"ff",	--12146
		x"ff",	--12147
		x"ff",	--12148
		x"ff",	--12149
		x"ff",	--12150
		x"ff",	--12151
		x"ff",	--12152
		x"ff",	--12153
		x"ff",	--12154
		x"ff",	--12155
		x"ff",	--12156
		x"ff",	--12157
		x"ff",	--12158
		x"ff",	--12159
		x"ff",	--12160
		x"ff",	--12161
		x"ff",	--12162
		x"ff",	--12163
		x"ff",	--12164
		x"ff",	--12165
		x"ff",	--12166
		x"ff",	--12167
		x"ff",	--12168
		x"ff",	--12169
		x"ff",	--12170
		x"ff",	--12171
		x"ff",	--12172
		x"ff",	--12173
		x"ff",	--12174
		x"ff",	--12175
		x"ff",	--12176
		x"ff",	--12177
		x"ff",	--12178
		x"ff",	--12179
		x"ff",	--12180
		x"ff",	--12181
		x"ff",	--12182
		x"ff",	--12183
		x"ff",	--12184
		x"ff",	--12185
		x"ff",	--12186
		x"ff",	--12187
		x"ff",	--12188
		x"ff",	--12189
		x"ff",	--12190
		x"ff",	--12191
		x"ff",	--12192
		x"ff",	--12193
		x"ff",	--12194
		x"ff",	--12195
		x"ff",	--12196
		x"ff",	--12197
		x"ff",	--12198
		x"ff",	--12199
		x"ff",	--12200
		x"ff",	--12201
		x"ff",	--12202
		x"ff",	--12203
		x"ff",	--12204
		x"ff",	--12205
		x"ff",	--12206
		x"ff",	--12207
		x"ff",	--12208
		x"ff",	--12209
		x"ff",	--12210
		x"ff",	--12211
		x"ff",	--12212
		x"ff",	--12213
		x"ff",	--12214
		x"ff",	--12215
		x"ff",	--12216
		x"ff",	--12217
		x"ff",	--12218
		x"ff",	--12219
		x"ff",	--12220
		x"ff",	--12221
		x"ff",	--12222
		x"ff",	--12223
		x"ff",	--12224
		x"ff",	--12225
		x"ff",	--12226
		x"ff",	--12227
		x"ff",	--12228
		x"ff",	--12229
		x"ff",	--12230
		x"ff",	--12231
		x"ff",	--12232
		x"ff",	--12233
		x"ff",	--12234
		x"ff",	--12235
		x"ff",	--12236
		x"ff",	--12237
		x"ff",	--12238
		x"ff",	--12239
		x"ff",	--12240
		x"ff",	--12241
		x"ff",	--12242
		x"ff",	--12243
		x"ff",	--12244
		x"ff",	--12245
		x"ff",	--12246
		x"ff",	--12247
		x"ff",	--12248
		x"ff",	--12249
		x"ff",	--12250
		x"ff",	--12251
		x"ff",	--12252
		x"ff",	--12253
		x"ff",	--12254
		x"ff",	--12255
		x"ff",	--12256
		x"ff",	--12257
		x"ff",	--12258
		x"ff",	--12259
		x"ff",	--12260
		x"ff",	--12261
		x"ff",	--12262
		x"ff",	--12263
		x"ff",	--12264
		x"ff",	--12265
		x"ff",	--12266
		x"ff",	--12267
		x"ff",	--12268
		x"ff",	--12269
		x"ff",	--12270
		x"ff",	--12271
		x"ff",	--12272
		x"ff",	--12273
		x"ff",	--12274
		x"ff",	--12275
		x"ff",	--12276
		x"ff",	--12277
		x"ff",	--12278
		x"ff",	--12279
		x"ff",	--12280
		x"ff",	--12281
		x"ff",	--12282
		x"ff",	--12283
		x"ff",	--12284
		x"ff",	--12285
		x"ff",	--12286
		x"ff",	--12287
		x"ff",	--12288
		x"ff",	--12289
		x"ff",	--12290
		x"ff",	--12291
		x"ff",	--12292
		x"ff",	--12293
		x"ff",	--12294
		x"ff",	--12295
		x"ff",	--12296
		x"ff",	--12297
		x"ff",	--12298
		x"ff",	--12299
		x"ff",	--12300
		x"ff",	--12301
		x"ff",	--12302
		x"ff",	--12303
		x"ff",	--12304
		x"ff",	--12305
		x"ff",	--12306
		x"ff",	--12307
		x"ff",	--12308
		x"ff",	--12309
		x"ff",	--12310
		x"ff",	--12311
		x"ff",	--12312
		x"ff",	--12313
		x"ff",	--12314
		x"ff",	--12315
		x"ff",	--12316
		x"ff",	--12317
		x"ff",	--12318
		x"ff",	--12319
		x"ff",	--12320
		x"ff",	--12321
		x"ff",	--12322
		x"ff",	--12323
		x"ff",	--12324
		x"ff",	--12325
		x"ff",	--12326
		x"ff",	--12327
		x"ff",	--12328
		x"ff",	--12329
		x"ff",	--12330
		x"ff",	--12331
		x"ff",	--12332
		x"ff",	--12333
		x"ff",	--12334
		x"ff",	--12335
		x"ff",	--12336
		x"ff",	--12337
		x"ff",	--12338
		x"ff",	--12339
		x"ff",	--12340
		x"ff",	--12341
		x"ff",	--12342
		x"ff",	--12343
		x"ff",	--12344
		x"ff",	--12345
		x"ff",	--12346
		x"ff",	--12347
		x"ff",	--12348
		x"ff",	--12349
		x"ff",	--12350
		x"ff",	--12351
		x"ff",	--12352
		x"ff",	--12353
		x"ff",	--12354
		x"ff",	--12355
		x"ff",	--12356
		x"ff",	--12357
		x"ff",	--12358
		x"ff",	--12359
		x"ff",	--12360
		x"ff",	--12361
		x"ff",	--12362
		x"ff",	--12363
		x"ff",	--12364
		x"ff",	--12365
		x"ff",	--12366
		x"ff",	--12367
		x"ff",	--12368
		x"ff",	--12369
		x"ff",	--12370
		x"ff",	--12371
		x"ff",	--12372
		x"ff",	--12373
		x"ff",	--12374
		x"ff",	--12375
		x"ff",	--12376
		x"ff",	--12377
		x"ff",	--12378
		x"ff",	--12379
		x"ff",	--12380
		x"ff",	--12381
		x"ff",	--12382
		x"ff",	--12383
		x"ff",	--12384
		x"ff",	--12385
		x"ff",	--12386
		x"ff",	--12387
		x"ff",	--12388
		x"ff",	--12389
		x"ff",	--12390
		x"ff",	--12391
		x"ff",	--12392
		x"ff",	--12393
		x"ff",	--12394
		x"ff",	--12395
		x"ff",	--12396
		x"ff",	--12397
		x"ff",	--12398
		x"ff",	--12399
		x"ff",	--12400
		x"ff",	--12401
		x"ff",	--12402
		x"ff",	--12403
		x"ff",	--12404
		x"ff",	--12405
		x"ff",	--12406
		x"ff",	--12407
		x"ff",	--12408
		x"ff",	--12409
		x"ff",	--12410
		x"ff",	--12411
		x"ff",	--12412
		x"ff",	--12413
		x"ff",	--12414
		x"ff",	--12415
		x"ff",	--12416
		x"ff",	--12417
		x"ff",	--12418
		x"ff",	--12419
		x"ff",	--12420
		x"ff",	--12421
		x"ff",	--12422
		x"ff",	--12423
		x"ff",	--12424
		x"ff",	--12425
		x"ff",	--12426
		x"ff",	--12427
		x"ff",	--12428
		x"ff",	--12429
		x"ff",	--12430
		x"ff",	--12431
		x"ff",	--12432
		x"ff",	--12433
		x"ff",	--12434
		x"ff",	--12435
		x"ff",	--12436
		x"ff",	--12437
		x"ff",	--12438
		x"ff",	--12439
		x"ff",	--12440
		x"ff",	--12441
		x"ff",	--12442
		x"ff",	--12443
		x"ff",	--12444
		x"ff",	--12445
		x"ff",	--12446
		x"ff",	--12447
		x"ff",	--12448
		x"ff",	--12449
		x"ff",	--12450
		x"ff",	--12451
		x"ff",	--12452
		x"ff",	--12453
		x"ff",	--12454
		x"ff",	--12455
		x"ff",	--12456
		x"ff",	--12457
		x"ff",	--12458
		x"ff",	--12459
		x"ff",	--12460
		x"ff",	--12461
		x"ff",	--12462
		x"ff",	--12463
		x"ff",	--12464
		x"ff",	--12465
		x"ff",	--12466
		x"ff",	--12467
		x"ff",	--12468
		x"ff",	--12469
		x"ff",	--12470
		x"ff",	--12471
		x"ff",	--12472
		x"ff",	--12473
		x"ff",	--12474
		x"ff",	--12475
		x"ff",	--12476
		x"ff",	--12477
		x"ff",	--12478
		x"ff",	--12479
		x"ff",	--12480
		x"ff",	--12481
		x"ff",	--12482
		x"ff",	--12483
		x"ff",	--12484
		x"ff",	--12485
		x"ff",	--12486
		x"ff",	--12487
		x"ff",	--12488
		x"ff",	--12489
		x"ff",	--12490
		x"ff",	--12491
		x"ff",	--12492
		x"ff",	--12493
		x"ff",	--12494
		x"ff",	--12495
		x"ff",	--12496
		x"ff",	--12497
		x"ff",	--12498
		x"ff",	--12499
		x"ff",	--12500
		x"ff",	--12501
		x"ff",	--12502
		x"ff",	--12503
		x"ff",	--12504
		x"ff",	--12505
		x"ff",	--12506
		x"ff",	--12507
		x"ff",	--12508
		x"ff",	--12509
		x"ff",	--12510
		x"ff",	--12511
		x"ff",	--12512
		x"ff",	--12513
		x"ff",	--12514
		x"ff",	--12515
		x"ff",	--12516
		x"ff",	--12517
		x"ff",	--12518
		x"ff",	--12519
		x"ff",	--12520
		x"ff",	--12521
		x"ff",	--12522
		x"ff",	--12523
		x"ff",	--12524
		x"ff",	--12525
		x"ff",	--12526
		x"ff",	--12527
		x"ff",	--12528
		x"ff",	--12529
		x"ff",	--12530
		x"ff",	--12531
		x"ff",	--12532
		x"ff",	--12533
		x"ff",	--12534
		x"ff",	--12535
		x"ff",	--12536
		x"ff",	--12537
		x"ff",	--12538
		x"ff",	--12539
		x"ff",	--12540
		x"ff",	--12541
		x"ff",	--12542
		x"ff",	--12543
		x"ff",	--12544
		x"ff",	--12545
		x"ff",	--12546
		x"ff",	--12547
		x"ff",	--12548
		x"ff",	--12549
		x"ff",	--12550
		x"ff",	--12551
		x"ff",	--12552
		x"ff",	--12553
		x"ff",	--12554
		x"ff",	--12555
		x"ff",	--12556
		x"ff",	--12557
		x"ff",	--12558
		x"ff",	--12559
		x"ff",	--12560
		x"ff",	--12561
		x"ff",	--12562
		x"ff",	--12563
		x"ff",	--12564
		x"ff",	--12565
		x"ff",	--12566
		x"ff",	--12567
		x"ff",	--12568
		x"ff",	--12569
		x"ff",	--12570
		x"ff",	--12571
		x"ff",	--12572
		x"ff",	--12573
		x"ff",	--12574
		x"ff",	--12575
		x"ff",	--12576
		x"ff",	--12577
		x"ff",	--12578
		x"ff",	--12579
		x"ff",	--12580
		x"ff",	--12581
		x"ff",	--12582
		x"ff",	--12583
		x"ff",	--12584
		x"ff",	--12585
		x"ff",	--12586
		x"ff",	--12587
		x"ff",	--12588
		x"ff",	--12589
		x"ff",	--12590
		x"ff",	--12591
		x"ff",	--12592
		x"ff",	--12593
		x"ff",	--12594
		x"ff",	--12595
		x"ff",	--12596
		x"ff",	--12597
		x"ff",	--12598
		x"ff",	--12599
		x"ff",	--12600
		x"ff",	--12601
		x"ff",	--12602
		x"ff",	--12603
		x"ff",	--12604
		x"ff",	--12605
		x"ff",	--12606
		x"ff",	--12607
		x"ff",	--12608
		x"ff",	--12609
		x"ff",	--12610
		x"ff",	--12611
		x"ff",	--12612
		x"ff",	--12613
		x"ff",	--12614
		x"ff",	--12615
		x"ff",	--12616
		x"ff",	--12617
		x"ff",	--12618
		x"ff",	--12619
		x"ff",	--12620
		x"ff",	--12621
		x"ff",	--12622
		x"ff",	--12623
		x"ff",	--12624
		x"ff",	--12625
		x"ff",	--12626
		x"ff",	--12627
		x"ff",	--12628
		x"ff",	--12629
		x"ff",	--12630
		x"ff",	--12631
		x"ff",	--12632
		x"ff",	--12633
		x"ff",	--12634
		x"ff",	--12635
		x"ff",	--12636
		x"ff",	--12637
		x"ff",	--12638
		x"ff",	--12639
		x"ff",	--12640
		x"ff",	--12641
		x"ff",	--12642
		x"ff",	--12643
		x"ff",	--12644
		x"ff",	--12645
		x"ff",	--12646
		x"ff",	--12647
		x"ff",	--12648
		x"ff",	--12649
		x"ff",	--12650
		x"ff",	--12651
		x"ff",	--12652
		x"ff",	--12653
		x"ff",	--12654
		x"ff",	--12655
		x"ff",	--12656
		x"ff",	--12657
		x"ff",	--12658
		x"ff",	--12659
		x"ff",	--12660
		x"ff",	--12661
		x"ff",	--12662
		x"ff",	--12663
		x"ff",	--12664
		x"ff",	--12665
		x"ff",	--12666
		x"ff",	--12667
		x"ff",	--12668
		x"ff",	--12669
		x"ff",	--12670
		x"ff",	--12671
		x"ff",	--12672
		x"ff",	--12673
		x"ff",	--12674
		x"ff",	--12675
		x"ff",	--12676
		x"ff",	--12677
		x"ff",	--12678
		x"ff",	--12679
		x"ff",	--12680
		x"ff",	--12681
		x"ff",	--12682
		x"ff",	--12683
		x"ff",	--12684
		x"ff",	--12685
		x"ff",	--12686
		x"ff",	--12687
		x"ff",	--12688
		x"ff",	--12689
		x"ff",	--12690
		x"ff",	--12691
		x"ff",	--12692
		x"ff",	--12693
		x"ff",	--12694
		x"ff",	--12695
		x"ff",	--12696
		x"ff",	--12697
		x"ff",	--12698
		x"ff",	--12699
		x"ff",	--12700
		x"ff",	--12701
		x"ff",	--12702
		x"ff",	--12703
		x"ff",	--12704
		x"ff",	--12705
		x"ff",	--12706
		x"ff",	--12707
		x"ff",	--12708
		x"ff",	--12709
		x"ff",	--12710
		x"ff",	--12711
		x"ff",	--12712
		x"ff",	--12713
		x"ff",	--12714
		x"ff",	--12715
		x"ff",	--12716
		x"ff",	--12717
		x"ff",	--12718
		x"ff",	--12719
		x"ff",	--12720
		x"ff",	--12721
		x"ff",	--12722
		x"ff",	--12723
		x"ff",	--12724
		x"ff",	--12725
		x"ff",	--12726
		x"ff",	--12727
		x"ff",	--12728
		x"ff",	--12729
		x"ff",	--12730
		x"ff",	--12731
		x"ff",	--12732
		x"ff",	--12733
		x"ff",	--12734
		x"ff",	--12735
		x"ff",	--12736
		x"ff",	--12737
		x"ff",	--12738
		x"ff",	--12739
		x"ff",	--12740
		x"ff",	--12741
		x"ff",	--12742
		x"ff",	--12743
		x"ff",	--12744
		x"ff",	--12745
		x"ff",	--12746
		x"ff",	--12747
		x"ff",	--12748
		x"ff",	--12749
		x"ff",	--12750
		x"ff",	--12751
		x"ff",	--12752
		x"ff",	--12753
		x"ff",	--12754
		x"ff",	--12755
		x"ff",	--12756
		x"ff",	--12757
		x"ff",	--12758
		x"ff",	--12759
		x"ff",	--12760
		x"ff",	--12761
		x"ff",	--12762
		x"ff",	--12763
		x"ff",	--12764
		x"ff",	--12765
		x"ff",	--12766
		x"ff",	--12767
		x"ff",	--12768
		x"ff",	--12769
		x"ff",	--12770
		x"ff",	--12771
		x"ff",	--12772
		x"ff",	--12773
		x"ff",	--12774
		x"ff",	--12775
		x"ff",	--12776
		x"ff",	--12777
		x"ff",	--12778
		x"ff",	--12779
		x"ff",	--12780
		x"ff",	--12781
		x"ff",	--12782
		x"ff",	--12783
		x"ff",	--12784
		x"ff",	--12785
		x"ff",	--12786
		x"ff",	--12787
		x"ff",	--12788
		x"ff",	--12789
		x"ff",	--12790
		x"ff",	--12791
		x"ff",	--12792
		x"ff",	--12793
		x"ff",	--12794
		x"ff",	--12795
		x"ff",	--12796
		x"ff",	--12797
		x"ff",	--12798
		x"ff",	--12799
		x"ff",	--12800
		x"ff",	--12801
		x"ff",	--12802
		x"ff",	--12803
		x"ff",	--12804
		x"ff",	--12805
		x"ff",	--12806
		x"ff",	--12807
		x"ff",	--12808
		x"ff",	--12809
		x"ff",	--12810
		x"ff",	--12811
		x"ff",	--12812
		x"ff",	--12813
		x"ff",	--12814
		x"ff",	--12815
		x"ff",	--12816
		x"ff",	--12817
		x"ff",	--12818
		x"ff",	--12819
		x"ff",	--12820
		x"ff",	--12821
		x"ff",	--12822
		x"ff",	--12823
		x"ff",	--12824
		x"ff",	--12825
		x"ff",	--12826
		x"ff",	--12827
		x"ff",	--12828
		x"ff",	--12829
		x"ff",	--12830
		x"ff",	--12831
		x"ff",	--12832
		x"ff",	--12833
		x"ff",	--12834
		x"ff",	--12835
		x"ff",	--12836
		x"ff",	--12837
		x"ff",	--12838
		x"ff",	--12839
		x"ff",	--12840
		x"ff",	--12841
		x"ff",	--12842
		x"ff",	--12843
		x"ff",	--12844
		x"ff",	--12845
		x"ff",	--12846
		x"ff",	--12847
		x"ff",	--12848
		x"ff",	--12849
		x"ff",	--12850
		x"ff",	--12851
		x"ff",	--12852
		x"ff",	--12853
		x"ff",	--12854
		x"ff",	--12855
		x"ff",	--12856
		x"ff",	--12857
		x"ff",	--12858
		x"ff",	--12859
		x"ff",	--12860
		x"ff",	--12861
		x"ff",	--12862
		x"ff",	--12863
		x"ff",	--12864
		x"ff",	--12865
		x"ff",	--12866
		x"ff",	--12867
		x"ff",	--12868
		x"ff",	--12869
		x"ff",	--12870
		x"ff",	--12871
		x"ff",	--12872
		x"ff",	--12873
		x"ff",	--12874
		x"ff",	--12875
		x"ff",	--12876
		x"ff",	--12877
		x"ff",	--12878
		x"ff",	--12879
		x"ff",	--12880
		x"ff",	--12881
		x"ff",	--12882
		x"ff",	--12883
		x"ff",	--12884
		x"ff",	--12885
		x"ff",	--12886
		x"ff",	--12887
		x"ff",	--12888
		x"ff",	--12889
		x"ff",	--12890
		x"ff",	--12891
		x"ff",	--12892
		x"ff",	--12893
		x"ff",	--12894
		x"ff",	--12895
		x"ff",	--12896
		x"ff",	--12897
		x"ff",	--12898
		x"ff",	--12899
		x"ff",	--12900
		x"ff",	--12901
		x"ff",	--12902
		x"ff",	--12903
		x"ff",	--12904
		x"ff",	--12905
		x"ff",	--12906
		x"ff",	--12907
		x"ff",	--12908
		x"ff",	--12909
		x"ff",	--12910
		x"ff",	--12911
		x"ff",	--12912
		x"ff",	--12913
		x"ff",	--12914
		x"ff",	--12915
		x"ff",	--12916
		x"ff",	--12917
		x"ff",	--12918
		x"ff",	--12919
		x"ff",	--12920
		x"ff",	--12921
		x"ff",	--12922
		x"ff",	--12923
		x"ff",	--12924
		x"ff",	--12925
		x"ff",	--12926
		x"ff",	--12927
		x"ff",	--12928
		x"ff",	--12929
		x"ff",	--12930
		x"ff",	--12931
		x"ff",	--12932
		x"ff",	--12933
		x"ff",	--12934
		x"ff",	--12935
		x"ff",	--12936
		x"ff",	--12937
		x"ff",	--12938
		x"ff",	--12939
		x"ff",	--12940
		x"ff",	--12941
		x"ff",	--12942
		x"ff",	--12943
		x"ff",	--12944
		x"ff",	--12945
		x"ff",	--12946
		x"ff",	--12947
		x"ff",	--12948
		x"ff",	--12949
		x"ff",	--12950
		x"ff",	--12951
		x"ff",	--12952
		x"ff",	--12953
		x"ff",	--12954
		x"ff",	--12955
		x"ff",	--12956
		x"ff",	--12957
		x"ff",	--12958
		x"ff",	--12959
		x"ff",	--12960
		x"ff",	--12961
		x"ff",	--12962
		x"ff",	--12963
		x"ff",	--12964
		x"ff",	--12965
		x"ff",	--12966
		x"ff",	--12967
		x"ff",	--12968
		x"ff",	--12969
		x"ff",	--12970
		x"ff",	--12971
		x"ff",	--12972
		x"ff",	--12973
		x"ff",	--12974
		x"ff",	--12975
		x"ff",	--12976
		x"ff",	--12977
		x"ff",	--12978
		x"ff",	--12979
		x"ff",	--12980
		x"ff",	--12981
		x"ff",	--12982
		x"ff",	--12983
		x"ff",	--12984
		x"ff",	--12985
		x"ff",	--12986
		x"ff",	--12987
		x"ff",	--12988
		x"ff",	--12989
		x"ff",	--12990
		x"ff",	--12991
		x"ff",	--12992
		x"ff",	--12993
		x"ff",	--12994
		x"ff",	--12995
		x"ff",	--12996
		x"ff",	--12997
		x"ff",	--12998
		x"ff",	--12999
		x"ff",	--13000
		x"ff",	--13001
		x"ff",	--13002
		x"ff",	--13003
		x"ff",	--13004
		x"ff",	--13005
		x"ff",	--13006
		x"ff",	--13007
		x"ff",	--13008
		x"ff",	--13009
		x"ff",	--13010
		x"ff",	--13011
		x"ff",	--13012
		x"ff",	--13013
		x"ff",	--13014
		x"ff",	--13015
		x"ff",	--13016
		x"ff",	--13017
		x"ff",	--13018
		x"ff",	--13019
		x"ff",	--13020
		x"ff",	--13021
		x"ff",	--13022
		x"ff",	--13023
		x"ff",	--13024
		x"ff",	--13025
		x"ff",	--13026
		x"ff",	--13027
		x"ff",	--13028
		x"ff",	--13029
		x"ff",	--13030
		x"ff",	--13031
		x"ff",	--13032
		x"ff",	--13033
		x"ff",	--13034
		x"ff",	--13035
		x"ff",	--13036
		x"ff",	--13037
		x"ff",	--13038
		x"ff",	--13039
		x"ff",	--13040
		x"ff",	--13041
		x"ff",	--13042
		x"ff",	--13043
		x"ff",	--13044
		x"ff",	--13045
		x"ff",	--13046
		x"ff",	--13047
		x"ff",	--13048
		x"ff",	--13049
		x"ff",	--13050
		x"ff",	--13051
		x"ff",	--13052
		x"ff",	--13053
		x"ff",	--13054
		x"ff",	--13055
		x"ff",	--13056
		x"ff",	--13057
		x"ff",	--13058
		x"ff",	--13059
		x"ff",	--13060
		x"ff",	--13061
		x"ff",	--13062
		x"ff",	--13063
		x"ff",	--13064
		x"ff",	--13065
		x"ff",	--13066
		x"ff",	--13067
		x"ff",	--13068
		x"ff",	--13069
		x"ff",	--13070
		x"ff",	--13071
		x"ff",	--13072
		x"ff",	--13073
		x"ff",	--13074
		x"ff",	--13075
		x"ff",	--13076
		x"ff",	--13077
		x"ff",	--13078
		x"ff",	--13079
		x"ff",	--13080
		x"ff",	--13081
		x"ff",	--13082
		x"ff",	--13083
		x"ff",	--13084
		x"ff",	--13085
		x"ff",	--13086
		x"ff",	--13087
		x"ff",	--13088
		x"ff",	--13089
		x"ff",	--13090
		x"ff",	--13091
		x"ff",	--13092
		x"ff",	--13093
		x"ff",	--13094
		x"ff",	--13095
		x"ff",	--13096
		x"ff",	--13097
		x"ff",	--13098
		x"ff",	--13099
		x"ff",	--13100
		x"ff",	--13101
		x"ff",	--13102
		x"ff",	--13103
		x"ff",	--13104
		x"ff",	--13105
		x"ff",	--13106
		x"ff",	--13107
		x"ff",	--13108
		x"ff",	--13109
		x"ff",	--13110
		x"ff",	--13111
		x"ff",	--13112
		x"ff",	--13113
		x"ff",	--13114
		x"ff",	--13115
		x"ff",	--13116
		x"ff",	--13117
		x"ff",	--13118
		x"ff",	--13119
		x"ff",	--13120
		x"ff",	--13121
		x"ff",	--13122
		x"ff",	--13123
		x"ff",	--13124
		x"ff",	--13125
		x"ff",	--13126
		x"ff",	--13127
		x"ff",	--13128
		x"ff",	--13129
		x"ff",	--13130
		x"ff",	--13131
		x"ff",	--13132
		x"ff",	--13133
		x"ff",	--13134
		x"ff",	--13135
		x"ff",	--13136
		x"ff",	--13137
		x"ff",	--13138
		x"ff",	--13139
		x"ff",	--13140
		x"ff",	--13141
		x"ff",	--13142
		x"ff",	--13143
		x"ff",	--13144
		x"ff",	--13145
		x"ff",	--13146
		x"ff",	--13147
		x"ff",	--13148
		x"ff",	--13149
		x"ff",	--13150
		x"ff",	--13151
		x"ff",	--13152
		x"ff",	--13153
		x"ff",	--13154
		x"ff",	--13155
		x"ff",	--13156
		x"ff",	--13157
		x"ff",	--13158
		x"ff",	--13159
		x"ff",	--13160
		x"ff",	--13161
		x"ff",	--13162
		x"ff",	--13163
		x"ff",	--13164
		x"ff",	--13165
		x"ff",	--13166
		x"ff",	--13167
		x"ff",	--13168
		x"ff",	--13169
		x"ff",	--13170
		x"ff",	--13171
		x"ff",	--13172
		x"ff",	--13173
		x"ff",	--13174
		x"ff",	--13175
		x"ff",	--13176
		x"ff",	--13177
		x"ff",	--13178
		x"ff",	--13179
		x"ff",	--13180
		x"ff",	--13181
		x"ff",	--13182
		x"ff",	--13183
		x"ff",	--13184
		x"ff",	--13185
		x"ff",	--13186
		x"ff",	--13187
		x"ff",	--13188
		x"ff",	--13189
		x"ff",	--13190
		x"ff",	--13191
		x"ff",	--13192
		x"ff",	--13193
		x"ff",	--13194
		x"ff",	--13195
		x"ff",	--13196
		x"ff",	--13197
		x"ff",	--13198
		x"ff",	--13199
		x"ff",	--13200
		x"ff",	--13201
		x"ff",	--13202
		x"ff",	--13203
		x"ff",	--13204
		x"ff",	--13205
		x"ff",	--13206
		x"ff",	--13207
		x"ff",	--13208
		x"ff",	--13209
		x"ff",	--13210
		x"ff",	--13211
		x"ff",	--13212
		x"ff",	--13213
		x"ff",	--13214
		x"ff",	--13215
		x"ff",	--13216
		x"ff",	--13217
		x"ff",	--13218
		x"ff",	--13219
		x"ff",	--13220
		x"ff",	--13221
		x"ff",	--13222
		x"ff",	--13223
		x"ff",	--13224
		x"ff",	--13225
		x"ff",	--13226
		x"ff",	--13227
		x"ff",	--13228
		x"ff",	--13229
		x"ff",	--13230
		x"ff",	--13231
		x"ff",	--13232
		x"ff",	--13233
		x"ff",	--13234
		x"ff",	--13235
		x"ff",	--13236
		x"ff",	--13237
		x"ff",	--13238
		x"ff",	--13239
		x"ff",	--13240
		x"ff",	--13241
		x"ff",	--13242
		x"ff",	--13243
		x"ff",	--13244
		x"ff",	--13245
		x"ff",	--13246
		x"ff",	--13247
		x"ff",	--13248
		x"ff",	--13249
		x"ff",	--13250
		x"ff",	--13251
		x"ff",	--13252
		x"ff",	--13253
		x"ff",	--13254
		x"ff",	--13255
		x"ff",	--13256
		x"ff",	--13257
		x"ff",	--13258
		x"ff",	--13259
		x"ff",	--13260
		x"ff",	--13261
		x"ff",	--13262
		x"ff",	--13263
		x"ff",	--13264
		x"ff",	--13265
		x"ff",	--13266
		x"ff",	--13267
		x"ff",	--13268
		x"ff",	--13269
		x"ff",	--13270
		x"ff",	--13271
		x"ff",	--13272
		x"ff",	--13273
		x"ff",	--13274
		x"ff",	--13275
		x"ff",	--13276
		x"ff",	--13277
		x"ff",	--13278
		x"ff",	--13279
		x"ff",	--13280
		x"ff",	--13281
		x"ff",	--13282
		x"ff",	--13283
		x"ff",	--13284
		x"ff",	--13285
		x"ff",	--13286
		x"ff",	--13287
		x"ff",	--13288
		x"ff",	--13289
		x"ff",	--13290
		x"ff",	--13291
		x"ff",	--13292
		x"ff",	--13293
		x"ff",	--13294
		x"ff",	--13295
		x"ff",	--13296
		x"ff",	--13297
		x"ff",	--13298
		x"ff",	--13299
		x"ff",	--13300
		x"ff",	--13301
		x"ff",	--13302
		x"ff",	--13303
		x"ff",	--13304
		x"ff",	--13305
		x"ff",	--13306
		x"ff",	--13307
		x"ff",	--13308
		x"ff",	--13309
		x"ff",	--13310
		x"ff",	--13311
		x"ff",	--13312
		x"ff",	--13313
		x"ff",	--13314
		x"ff",	--13315
		x"ff",	--13316
		x"ff",	--13317
		x"ff",	--13318
		x"ff",	--13319
		x"ff",	--13320
		x"ff",	--13321
		x"ff",	--13322
		x"ff",	--13323
		x"ff",	--13324
		x"ff",	--13325
		x"ff",	--13326
		x"ff",	--13327
		x"ff",	--13328
		x"ff",	--13329
		x"ff",	--13330
		x"ff",	--13331
		x"ff",	--13332
		x"ff",	--13333
		x"ff",	--13334
		x"ff",	--13335
		x"ff",	--13336
		x"ff",	--13337
		x"ff",	--13338
		x"ff",	--13339
		x"ff",	--13340
		x"ff",	--13341
		x"ff",	--13342
		x"ff",	--13343
		x"ff",	--13344
		x"ff",	--13345
		x"ff",	--13346
		x"ff",	--13347
		x"ff",	--13348
		x"ff",	--13349
		x"ff",	--13350
		x"ff",	--13351
		x"ff",	--13352
		x"ff",	--13353
		x"ff",	--13354
		x"ff",	--13355
		x"ff",	--13356
		x"ff",	--13357
		x"ff",	--13358
		x"ff",	--13359
		x"ff",	--13360
		x"ff",	--13361
		x"ff",	--13362
		x"ff",	--13363
		x"ff",	--13364
		x"ff",	--13365
		x"ff",	--13366
		x"ff",	--13367
		x"ff",	--13368
		x"ff",	--13369
		x"ff",	--13370
		x"ff",	--13371
		x"ff",	--13372
		x"ff",	--13373
		x"ff",	--13374
		x"ff",	--13375
		x"ff",	--13376
		x"ff",	--13377
		x"ff",	--13378
		x"ff",	--13379
		x"ff",	--13380
		x"ff",	--13381
		x"ff",	--13382
		x"ff",	--13383
		x"ff",	--13384
		x"ff",	--13385
		x"ff",	--13386
		x"ff",	--13387
		x"ff",	--13388
		x"ff",	--13389
		x"ff",	--13390
		x"ff",	--13391
		x"ff",	--13392
		x"ff",	--13393
		x"ff",	--13394
		x"ff",	--13395
		x"ff",	--13396
		x"ff",	--13397
		x"ff",	--13398
		x"ff",	--13399
		x"ff",	--13400
		x"ff",	--13401
		x"ff",	--13402
		x"ff",	--13403
		x"ff",	--13404
		x"ff",	--13405
		x"ff",	--13406
		x"ff",	--13407
		x"ff",	--13408
		x"ff",	--13409
		x"ff",	--13410
		x"ff",	--13411
		x"ff",	--13412
		x"ff",	--13413
		x"ff",	--13414
		x"ff",	--13415
		x"ff",	--13416
		x"ff",	--13417
		x"ff",	--13418
		x"ff",	--13419
		x"ff",	--13420
		x"ff",	--13421
		x"ff",	--13422
		x"ff",	--13423
		x"ff",	--13424
		x"ff",	--13425
		x"ff",	--13426
		x"ff",	--13427
		x"ff",	--13428
		x"ff",	--13429
		x"ff",	--13430
		x"ff",	--13431
		x"ff",	--13432
		x"ff",	--13433
		x"ff",	--13434
		x"ff",	--13435
		x"ff",	--13436
		x"ff",	--13437
		x"ff",	--13438
		x"ff",	--13439
		x"ff",	--13440
		x"ff",	--13441
		x"ff",	--13442
		x"ff",	--13443
		x"ff",	--13444
		x"ff",	--13445
		x"ff",	--13446
		x"ff",	--13447
		x"ff",	--13448
		x"ff",	--13449
		x"ff",	--13450
		x"ff",	--13451
		x"ff",	--13452
		x"ff",	--13453
		x"ff",	--13454
		x"ff",	--13455
		x"ff",	--13456
		x"ff",	--13457
		x"ff",	--13458
		x"ff",	--13459
		x"ff",	--13460
		x"ff",	--13461
		x"ff",	--13462
		x"ff",	--13463
		x"ff",	--13464
		x"ff",	--13465
		x"ff",	--13466
		x"ff",	--13467
		x"ff",	--13468
		x"ff",	--13469
		x"ff",	--13470
		x"ff",	--13471
		x"ff",	--13472
		x"ff",	--13473
		x"ff",	--13474
		x"ff",	--13475
		x"ff",	--13476
		x"ff",	--13477
		x"ff",	--13478
		x"ff",	--13479
		x"ff",	--13480
		x"ff",	--13481
		x"ff",	--13482
		x"ff",	--13483
		x"ff",	--13484
		x"ff",	--13485
		x"ff",	--13486
		x"ff",	--13487
		x"ff",	--13488
		x"ff",	--13489
		x"ff",	--13490
		x"ff",	--13491
		x"ff",	--13492
		x"ff",	--13493
		x"ff",	--13494
		x"ff",	--13495
		x"ff",	--13496
		x"ff",	--13497
		x"ff",	--13498
		x"ff",	--13499
		x"ff",	--13500
		x"ff",	--13501
		x"ff",	--13502
		x"ff",	--13503
		x"ff",	--13504
		x"ff",	--13505
		x"ff",	--13506
		x"ff",	--13507
		x"ff",	--13508
		x"ff",	--13509
		x"ff",	--13510
		x"ff",	--13511
		x"ff",	--13512
		x"ff",	--13513
		x"ff",	--13514
		x"ff",	--13515
		x"ff",	--13516
		x"ff",	--13517
		x"ff",	--13518
		x"ff",	--13519
		x"ff",	--13520
		x"ff",	--13521
		x"ff",	--13522
		x"ff",	--13523
		x"ff",	--13524
		x"ff",	--13525
		x"ff",	--13526
		x"ff",	--13527
		x"ff",	--13528
		x"ff",	--13529
		x"ff",	--13530
		x"ff",	--13531
		x"ff",	--13532
		x"ff",	--13533
		x"ff",	--13534
		x"ff",	--13535
		x"ff",	--13536
		x"ff",	--13537
		x"ff",	--13538
		x"ff",	--13539
		x"ff",	--13540
		x"ff",	--13541
		x"ff",	--13542
		x"ff",	--13543
		x"ff",	--13544
		x"ff",	--13545
		x"ff",	--13546
		x"ff",	--13547
		x"ff",	--13548
		x"ff",	--13549
		x"ff",	--13550
		x"ff",	--13551
		x"ff",	--13552
		x"ff",	--13553
		x"ff",	--13554
		x"ff",	--13555
		x"ff",	--13556
		x"ff",	--13557
		x"ff",	--13558
		x"ff",	--13559
		x"ff",	--13560
		x"ff",	--13561
		x"ff",	--13562
		x"ff",	--13563
		x"ff",	--13564
		x"ff",	--13565
		x"ff",	--13566
		x"ff",	--13567
		x"ff",	--13568
		x"ff",	--13569
		x"ff",	--13570
		x"ff",	--13571
		x"ff",	--13572
		x"ff",	--13573
		x"ff",	--13574
		x"ff",	--13575
		x"ff",	--13576
		x"ff",	--13577
		x"ff",	--13578
		x"ff",	--13579
		x"ff",	--13580
		x"ff",	--13581
		x"ff",	--13582
		x"ff",	--13583
		x"ff",	--13584
		x"ff",	--13585
		x"ff",	--13586
		x"ff",	--13587
		x"ff",	--13588
		x"ff",	--13589
		x"ff",	--13590
		x"ff",	--13591
		x"ff",	--13592
		x"ff",	--13593
		x"ff",	--13594
		x"ff",	--13595
		x"ff",	--13596
		x"ff",	--13597
		x"ff",	--13598
		x"ff",	--13599
		x"ff",	--13600
		x"ff",	--13601
		x"ff",	--13602
		x"ff",	--13603
		x"ff",	--13604
		x"ff",	--13605
		x"ff",	--13606
		x"ff",	--13607
		x"ff",	--13608
		x"ff",	--13609
		x"ff",	--13610
		x"ff",	--13611
		x"ff",	--13612
		x"ff",	--13613
		x"ff",	--13614
		x"ff",	--13615
		x"ff",	--13616
		x"ff",	--13617
		x"ff",	--13618
		x"ff",	--13619
		x"ff",	--13620
		x"ff",	--13621
		x"ff",	--13622
		x"ff",	--13623
		x"ff",	--13624
		x"ff",	--13625
		x"ff",	--13626
		x"ff",	--13627
		x"ff",	--13628
		x"ff",	--13629
		x"ff",	--13630
		x"ff",	--13631
		x"ff",	--13632
		x"ff",	--13633
		x"ff",	--13634
		x"ff",	--13635
		x"ff",	--13636
		x"ff",	--13637
		x"ff",	--13638
		x"ff",	--13639
		x"ff",	--13640
		x"ff",	--13641
		x"ff",	--13642
		x"ff",	--13643
		x"ff",	--13644
		x"ff",	--13645
		x"ff",	--13646
		x"ff",	--13647
		x"ff",	--13648
		x"ff",	--13649
		x"ff",	--13650
		x"ff",	--13651
		x"ff",	--13652
		x"ff",	--13653
		x"ff",	--13654
		x"ff",	--13655
		x"ff",	--13656
		x"ff",	--13657
		x"ff",	--13658
		x"ff",	--13659
		x"ff",	--13660
		x"ff",	--13661
		x"ff",	--13662
		x"ff",	--13663
		x"ff",	--13664
		x"ff",	--13665
		x"ff",	--13666
		x"ff",	--13667
		x"ff",	--13668
		x"ff",	--13669
		x"ff",	--13670
		x"ff",	--13671
		x"ff",	--13672
		x"ff",	--13673
		x"ff",	--13674
		x"ff",	--13675
		x"ff",	--13676
		x"ff",	--13677
		x"ff",	--13678
		x"ff",	--13679
		x"ff",	--13680
		x"ff",	--13681
		x"ff",	--13682
		x"ff",	--13683
		x"ff",	--13684
		x"ff",	--13685
		x"ff",	--13686
		x"ff",	--13687
		x"ff",	--13688
		x"ff",	--13689
		x"ff",	--13690
		x"ff",	--13691
		x"ff",	--13692
		x"ff",	--13693
		x"ff",	--13694
		x"ff",	--13695
		x"ff",	--13696
		x"ff",	--13697
		x"ff",	--13698
		x"ff",	--13699
		x"ff",	--13700
		x"ff",	--13701
		x"ff",	--13702
		x"ff",	--13703
		x"ff",	--13704
		x"ff",	--13705
		x"ff",	--13706
		x"ff",	--13707
		x"ff",	--13708
		x"ff",	--13709
		x"ff",	--13710
		x"ff",	--13711
		x"ff",	--13712
		x"ff",	--13713
		x"ff",	--13714
		x"ff",	--13715
		x"ff",	--13716
		x"ff",	--13717
		x"ff",	--13718
		x"ff",	--13719
		x"ff",	--13720
		x"ff",	--13721
		x"ff",	--13722
		x"ff",	--13723
		x"ff",	--13724
		x"ff",	--13725
		x"ff",	--13726
		x"ff",	--13727
		x"ff",	--13728
		x"ff",	--13729
		x"ff",	--13730
		x"ff",	--13731
		x"ff",	--13732
		x"ff",	--13733
		x"ff",	--13734
		x"ff",	--13735
		x"ff",	--13736
		x"ff",	--13737
		x"ff",	--13738
		x"ff",	--13739
		x"ff",	--13740
		x"ff",	--13741
		x"ff",	--13742
		x"ff",	--13743
		x"ff",	--13744
		x"ff",	--13745
		x"ff",	--13746
		x"ff",	--13747
		x"ff",	--13748
		x"ff",	--13749
		x"ff",	--13750
		x"ff",	--13751
		x"ff",	--13752
		x"ff",	--13753
		x"ff",	--13754
		x"ff",	--13755
		x"ff",	--13756
		x"ff",	--13757
		x"ff",	--13758
		x"ff",	--13759
		x"ff",	--13760
		x"ff",	--13761
		x"ff",	--13762
		x"ff",	--13763
		x"ff",	--13764
		x"ff",	--13765
		x"ff",	--13766
		x"ff",	--13767
		x"ff",	--13768
		x"ff",	--13769
		x"ff",	--13770
		x"ff",	--13771
		x"ff",	--13772
		x"ff",	--13773
		x"ff",	--13774
		x"ff",	--13775
		x"ff",	--13776
		x"ff",	--13777
		x"ff",	--13778
		x"ff",	--13779
		x"ff",	--13780
		x"ff",	--13781
		x"ff",	--13782
		x"ff",	--13783
		x"ff",	--13784
		x"ff",	--13785
		x"ff",	--13786
		x"ff",	--13787
		x"ff",	--13788
		x"ff",	--13789
		x"ff",	--13790
		x"ff",	--13791
		x"ff",	--13792
		x"ff",	--13793
		x"ff",	--13794
		x"ff",	--13795
		x"ff",	--13796
		x"ff",	--13797
		x"ff",	--13798
		x"ff",	--13799
		x"ff",	--13800
		x"ff",	--13801
		x"ff",	--13802
		x"ff",	--13803
		x"ff",	--13804
		x"ff",	--13805
		x"ff",	--13806
		x"ff",	--13807
		x"ff",	--13808
		x"ff",	--13809
		x"ff",	--13810
		x"ff",	--13811
		x"ff",	--13812
		x"ff",	--13813
		x"ff",	--13814
		x"ff",	--13815
		x"ff",	--13816
		x"ff",	--13817
		x"ff",	--13818
		x"ff",	--13819
		x"ff",	--13820
		x"ff",	--13821
		x"ff",	--13822
		x"ff",	--13823
		x"ff",	--13824
		x"ff",	--13825
		x"ff",	--13826
		x"ff",	--13827
		x"ff",	--13828
		x"ff",	--13829
		x"ff",	--13830
		x"ff",	--13831
		x"ff",	--13832
		x"ff",	--13833
		x"ff",	--13834
		x"ff",	--13835
		x"ff",	--13836
		x"ff",	--13837
		x"ff",	--13838
		x"ff",	--13839
		x"ff",	--13840
		x"ff",	--13841
		x"ff",	--13842
		x"ff",	--13843
		x"ff",	--13844
		x"ff",	--13845
		x"ff",	--13846
		x"ff",	--13847
		x"ff",	--13848
		x"ff",	--13849
		x"ff",	--13850
		x"ff",	--13851
		x"ff",	--13852
		x"ff",	--13853
		x"ff",	--13854
		x"ff",	--13855
		x"ff",	--13856
		x"ff",	--13857
		x"ff",	--13858
		x"ff",	--13859
		x"ff",	--13860
		x"ff",	--13861
		x"ff",	--13862
		x"ff",	--13863
		x"ff",	--13864
		x"ff",	--13865
		x"ff",	--13866
		x"ff",	--13867
		x"ff",	--13868
		x"ff",	--13869
		x"ff",	--13870
		x"ff",	--13871
		x"ff",	--13872
		x"ff",	--13873
		x"ff",	--13874
		x"ff",	--13875
		x"ff",	--13876
		x"ff",	--13877
		x"ff",	--13878
		x"ff",	--13879
		x"ff",	--13880
		x"ff",	--13881
		x"ff",	--13882
		x"ff",	--13883
		x"ff",	--13884
		x"ff",	--13885
		x"ff",	--13886
		x"ff",	--13887
		x"ff",	--13888
		x"ff",	--13889
		x"ff",	--13890
		x"ff",	--13891
		x"ff",	--13892
		x"ff",	--13893
		x"ff",	--13894
		x"ff",	--13895
		x"ff",	--13896
		x"ff",	--13897
		x"ff",	--13898
		x"ff",	--13899
		x"ff",	--13900
		x"ff",	--13901
		x"ff",	--13902
		x"ff",	--13903
		x"ff",	--13904
		x"ff",	--13905
		x"ff",	--13906
		x"ff",	--13907
		x"ff",	--13908
		x"ff",	--13909
		x"ff",	--13910
		x"ff",	--13911
		x"ff",	--13912
		x"ff",	--13913
		x"ff",	--13914
		x"ff",	--13915
		x"ff",	--13916
		x"ff",	--13917
		x"ff",	--13918
		x"ff",	--13919
		x"ff",	--13920
		x"ff",	--13921
		x"ff",	--13922
		x"ff",	--13923
		x"ff",	--13924
		x"ff",	--13925
		x"ff",	--13926
		x"ff",	--13927
		x"ff",	--13928
		x"ff",	--13929
		x"ff",	--13930
		x"ff",	--13931
		x"ff",	--13932
		x"ff",	--13933
		x"ff",	--13934
		x"ff",	--13935
		x"ff",	--13936
		x"ff",	--13937
		x"ff",	--13938
		x"ff",	--13939
		x"ff",	--13940
		x"ff",	--13941
		x"ff",	--13942
		x"ff",	--13943
		x"ff",	--13944
		x"ff",	--13945
		x"ff",	--13946
		x"ff",	--13947
		x"ff",	--13948
		x"ff",	--13949
		x"ff",	--13950
		x"ff",	--13951
		x"ff",	--13952
		x"ff",	--13953
		x"ff",	--13954
		x"ff",	--13955
		x"ff",	--13956
		x"ff",	--13957
		x"ff",	--13958
		x"ff",	--13959
		x"ff",	--13960
		x"ff",	--13961
		x"ff",	--13962
		x"ff",	--13963
		x"ff",	--13964
		x"ff",	--13965
		x"ff",	--13966
		x"ff",	--13967
		x"ff",	--13968
		x"ff",	--13969
		x"ff",	--13970
		x"ff",	--13971
		x"ff",	--13972
		x"ff",	--13973
		x"ff",	--13974
		x"ff",	--13975
		x"ff",	--13976
		x"ff",	--13977
		x"ff",	--13978
		x"ff",	--13979
		x"ff",	--13980
		x"ff",	--13981
		x"ff",	--13982
		x"ff",	--13983
		x"ff",	--13984
		x"ff",	--13985
		x"ff",	--13986
		x"ff",	--13987
		x"ff",	--13988
		x"ff",	--13989
		x"ff",	--13990
		x"ff",	--13991
		x"ff",	--13992
		x"ff",	--13993
		x"ff",	--13994
		x"ff",	--13995
		x"ff",	--13996
		x"ff",	--13997
		x"ff",	--13998
		x"ff",	--13999
		x"ff",	--14000
		x"ff",	--14001
		x"ff",	--14002
		x"ff",	--14003
		x"ff",	--14004
		x"ff",	--14005
		x"ff",	--14006
		x"ff",	--14007
		x"ff",	--14008
		x"ff",	--14009
		x"ff",	--14010
		x"ff",	--14011
		x"ff",	--14012
		x"ff",	--14013
		x"ff",	--14014
		x"ff",	--14015
		x"ff",	--14016
		x"ff",	--14017
		x"ff",	--14018
		x"ff",	--14019
		x"ff",	--14020
		x"ff",	--14021
		x"ff",	--14022
		x"ff",	--14023
		x"ff",	--14024
		x"ff",	--14025
		x"ff",	--14026
		x"ff",	--14027
		x"ff",	--14028
		x"ff",	--14029
		x"ff",	--14030
		x"ff",	--14031
		x"ff",	--14032
		x"ff",	--14033
		x"ff",	--14034
		x"ff",	--14035
		x"ff",	--14036
		x"ff",	--14037
		x"ff",	--14038
		x"ff",	--14039
		x"ff",	--14040
		x"ff",	--14041
		x"ff",	--14042
		x"ff",	--14043
		x"ff",	--14044
		x"ff",	--14045
		x"ff",	--14046
		x"ff",	--14047
		x"ff",	--14048
		x"ff",	--14049
		x"ff",	--14050
		x"ff",	--14051
		x"ff",	--14052
		x"ff",	--14053
		x"ff",	--14054
		x"ff",	--14055
		x"ff",	--14056
		x"ff",	--14057
		x"ff",	--14058
		x"ff",	--14059
		x"ff",	--14060
		x"ff",	--14061
		x"ff",	--14062
		x"ff",	--14063
		x"ff",	--14064
		x"ff",	--14065
		x"ff",	--14066
		x"ff",	--14067
		x"ff",	--14068
		x"ff",	--14069
		x"ff",	--14070
		x"ff",	--14071
		x"ff",	--14072
		x"ff",	--14073
		x"ff",	--14074
		x"ff",	--14075
		x"ff",	--14076
		x"ff",	--14077
		x"ff",	--14078
		x"ff",	--14079
		x"ff",	--14080
		x"ff",	--14081
		x"ff",	--14082
		x"ff",	--14083
		x"ff",	--14084
		x"ff",	--14085
		x"ff",	--14086
		x"ff",	--14087
		x"ff",	--14088
		x"ff",	--14089
		x"ff",	--14090
		x"ff",	--14091
		x"ff",	--14092
		x"ff",	--14093
		x"ff",	--14094
		x"ff",	--14095
		x"ff",	--14096
		x"ff",	--14097
		x"ff",	--14098
		x"ff",	--14099
		x"ff",	--14100
		x"ff",	--14101
		x"ff",	--14102
		x"ff",	--14103
		x"ff",	--14104
		x"ff",	--14105
		x"ff",	--14106
		x"ff",	--14107
		x"ff",	--14108
		x"ff",	--14109
		x"ff",	--14110
		x"ff",	--14111
		x"ff",	--14112
		x"ff",	--14113
		x"ff",	--14114
		x"ff",	--14115
		x"ff",	--14116
		x"ff",	--14117
		x"ff",	--14118
		x"ff",	--14119
		x"ff",	--14120
		x"ff",	--14121
		x"ff",	--14122
		x"ff",	--14123
		x"ff",	--14124
		x"ff",	--14125
		x"ff",	--14126
		x"ff",	--14127
		x"ff",	--14128
		x"ff",	--14129
		x"ff",	--14130
		x"ff",	--14131
		x"ff",	--14132
		x"ff",	--14133
		x"ff",	--14134
		x"ff",	--14135
		x"ff",	--14136
		x"ff",	--14137
		x"ff",	--14138
		x"ff",	--14139
		x"ff",	--14140
		x"ff",	--14141
		x"ff",	--14142
		x"ff",	--14143
		x"ff",	--14144
		x"ff",	--14145
		x"ff",	--14146
		x"ff",	--14147
		x"ff",	--14148
		x"ff",	--14149
		x"ff",	--14150
		x"ff",	--14151
		x"ff",	--14152
		x"ff",	--14153
		x"ff",	--14154
		x"ff",	--14155
		x"ff",	--14156
		x"ff",	--14157
		x"ff",	--14158
		x"ff",	--14159
		x"ff",	--14160
		x"ff",	--14161
		x"ff",	--14162
		x"ff",	--14163
		x"ff",	--14164
		x"ff",	--14165
		x"ff",	--14166
		x"ff",	--14167
		x"ff",	--14168
		x"ff",	--14169
		x"ff",	--14170
		x"ff",	--14171
		x"ff",	--14172
		x"ff",	--14173
		x"ff",	--14174
		x"ff",	--14175
		x"ff",	--14176
		x"ff",	--14177
		x"ff",	--14178
		x"ff",	--14179
		x"ff",	--14180
		x"ff",	--14181
		x"ff",	--14182
		x"ff",	--14183
		x"ff",	--14184
		x"ff",	--14185
		x"ff",	--14186
		x"ff",	--14187
		x"ff",	--14188
		x"ff",	--14189
		x"ff",	--14190
		x"ff",	--14191
		x"ff",	--14192
		x"ff",	--14193
		x"ff",	--14194
		x"ff",	--14195
		x"ff",	--14196
		x"ff",	--14197
		x"ff",	--14198
		x"ff",	--14199
		x"ff",	--14200
		x"ff",	--14201
		x"ff",	--14202
		x"ff",	--14203
		x"ff",	--14204
		x"ff",	--14205
		x"ff",	--14206
		x"ff",	--14207
		x"ff",	--14208
		x"ff",	--14209
		x"ff",	--14210
		x"ff",	--14211
		x"ff",	--14212
		x"ff",	--14213
		x"ff",	--14214
		x"ff",	--14215
		x"ff",	--14216
		x"ff",	--14217
		x"ff",	--14218
		x"ff",	--14219
		x"ff",	--14220
		x"ff",	--14221
		x"ff",	--14222
		x"ff",	--14223
		x"ff",	--14224
		x"ff",	--14225
		x"ff",	--14226
		x"ff",	--14227
		x"ff",	--14228
		x"ff",	--14229
		x"ff",	--14230
		x"ff",	--14231
		x"ff",	--14232
		x"ff",	--14233
		x"ff",	--14234
		x"ff",	--14235
		x"ff",	--14236
		x"ff",	--14237
		x"ff",	--14238
		x"ff",	--14239
		x"ff",	--14240
		x"ff",	--14241
		x"ff",	--14242
		x"ff",	--14243
		x"ff",	--14244
		x"ff",	--14245
		x"ff",	--14246
		x"ff",	--14247
		x"ff",	--14248
		x"ff",	--14249
		x"ff",	--14250
		x"ff",	--14251
		x"ff",	--14252
		x"ff",	--14253
		x"ff",	--14254
		x"ff",	--14255
		x"ff",	--14256
		x"ff",	--14257
		x"ff",	--14258
		x"ff",	--14259
		x"ff",	--14260
		x"ff",	--14261
		x"ff",	--14262
		x"ff",	--14263
		x"ff",	--14264
		x"ff",	--14265
		x"ff",	--14266
		x"ff",	--14267
		x"ff",	--14268
		x"ff",	--14269
		x"ff",	--14270
		x"ff",	--14271
		x"ff",	--14272
		x"ff",	--14273
		x"ff",	--14274
		x"ff",	--14275
		x"ff",	--14276
		x"ff",	--14277
		x"ff",	--14278
		x"ff",	--14279
		x"ff",	--14280
		x"ff",	--14281
		x"ff",	--14282
		x"ff",	--14283
		x"ff",	--14284
		x"ff",	--14285
		x"ff",	--14286
		x"ff",	--14287
		x"ff",	--14288
		x"ff",	--14289
		x"ff",	--14290
		x"ff",	--14291
		x"ff",	--14292
		x"ff",	--14293
		x"ff",	--14294
		x"ff",	--14295
		x"ff",	--14296
		x"ff",	--14297
		x"ff",	--14298
		x"ff",	--14299
		x"ff",	--14300
		x"ff",	--14301
		x"ff",	--14302
		x"ff",	--14303
		x"ff",	--14304
		x"ff",	--14305
		x"ff",	--14306
		x"ff",	--14307
		x"ff",	--14308
		x"ff",	--14309
		x"ff",	--14310
		x"ff",	--14311
		x"ff",	--14312
		x"ff",	--14313
		x"ff",	--14314
		x"ff",	--14315
		x"ff",	--14316
		x"ff",	--14317
		x"ff",	--14318
		x"ff",	--14319
		x"ff",	--14320
		x"ff",	--14321
		x"ff",	--14322
		x"ff",	--14323
		x"ff",	--14324
		x"ff",	--14325
		x"ff",	--14326
		x"ff",	--14327
		x"ff",	--14328
		x"ff",	--14329
		x"ff",	--14330
		x"ff",	--14331
		x"ff",	--14332
		x"ff",	--14333
		x"ff",	--14334
		x"ff",	--14335
		x"ff",	--14336
		x"ff",	--14337
		x"ff",	--14338
		x"ff",	--14339
		x"ff",	--14340
		x"ff",	--14341
		x"ff",	--14342
		x"ff",	--14343
		x"ff",	--14344
		x"ff",	--14345
		x"ff",	--14346
		x"ff",	--14347
		x"ff",	--14348
		x"ff",	--14349
		x"ff",	--14350
		x"ff",	--14351
		x"ff",	--14352
		x"ff",	--14353
		x"ff",	--14354
		x"ff",	--14355
		x"ff",	--14356
		x"ff",	--14357
		x"ff",	--14358
		x"ff",	--14359
		x"ff",	--14360
		x"ff",	--14361
		x"ff",	--14362
		x"ff",	--14363
		x"ff",	--14364
		x"ff",	--14365
		x"ff",	--14366
		x"ff",	--14367
		x"ff",	--14368
		x"ff",	--14369
		x"ff",	--14370
		x"ff",	--14371
		x"ff",	--14372
		x"ff",	--14373
		x"ff",	--14374
		x"ff",	--14375
		x"ff",	--14376
		x"ff",	--14377
		x"ff",	--14378
		x"ff",	--14379
		x"ff",	--14380
		x"ff",	--14381
		x"ff",	--14382
		x"ff",	--14383
		x"ff",	--14384
		x"ff",	--14385
		x"ff",	--14386
		x"ff",	--14387
		x"ff",	--14388
		x"ff",	--14389
		x"ff",	--14390
		x"ff",	--14391
		x"ff",	--14392
		x"ff",	--14393
		x"ff",	--14394
		x"ff",	--14395
		x"ff",	--14396
		x"ff",	--14397
		x"ff",	--14398
		x"ff",	--14399
		x"ff",	--14400
		x"ff",	--14401
		x"ff",	--14402
		x"ff",	--14403
		x"ff",	--14404
		x"ff",	--14405
		x"ff",	--14406
		x"ff",	--14407
		x"ff",	--14408
		x"ff",	--14409
		x"ff",	--14410
		x"ff",	--14411
		x"ff",	--14412
		x"ff",	--14413
		x"ff",	--14414
		x"ff",	--14415
		x"ff",	--14416
		x"ff",	--14417
		x"ff",	--14418
		x"ff",	--14419
		x"ff",	--14420
		x"ff",	--14421
		x"ff",	--14422
		x"ff",	--14423
		x"ff",	--14424
		x"ff",	--14425
		x"ff",	--14426
		x"ff",	--14427
		x"ff",	--14428
		x"ff",	--14429
		x"ff",	--14430
		x"ff",	--14431
		x"ff",	--14432
		x"ff",	--14433
		x"ff",	--14434
		x"ff",	--14435
		x"ff",	--14436
		x"ff",	--14437
		x"ff",	--14438
		x"ff",	--14439
		x"ff",	--14440
		x"ff",	--14441
		x"ff",	--14442
		x"ff",	--14443
		x"ff",	--14444
		x"ff",	--14445
		x"ff",	--14446
		x"ff",	--14447
		x"ff",	--14448
		x"ff",	--14449
		x"ff",	--14450
		x"ff",	--14451
		x"ff",	--14452
		x"ff",	--14453
		x"ff",	--14454
		x"ff",	--14455
		x"ff",	--14456
		x"ff",	--14457
		x"ff",	--14458
		x"ff",	--14459
		x"ff",	--14460
		x"ff",	--14461
		x"ff",	--14462
		x"ff",	--14463
		x"ff",	--14464
		x"ff",	--14465
		x"ff",	--14466
		x"ff",	--14467
		x"ff",	--14468
		x"ff",	--14469
		x"ff",	--14470
		x"ff",	--14471
		x"ff",	--14472
		x"ff",	--14473
		x"ff",	--14474
		x"ff",	--14475
		x"ff",	--14476
		x"ff",	--14477
		x"ff",	--14478
		x"ff",	--14479
		x"ff",	--14480
		x"ff",	--14481
		x"ff",	--14482
		x"ff",	--14483
		x"ff",	--14484
		x"ff",	--14485
		x"ff",	--14486
		x"ff",	--14487
		x"ff",	--14488
		x"ff",	--14489
		x"ff",	--14490
		x"ff",	--14491
		x"ff",	--14492
		x"ff",	--14493
		x"ff",	--14494
		x"ff",	--14495
		x"ff",	--14496
		x"ff",	--14497
		x"ff",	--14498
		x"ff",	--14499
		x"ff",	--14500
		x"ff",	--14501
		x"ff",	--14502
		x"ff",	--14503
		x"ff",	--14504
		x"ff",	--14505
		x"ff",	--14506
		x"ff",	--14507
		x"ff",	--14508
		x"ff",	--14509
		x"ff",	--14510
		x"ff",	--14511
		x"ff",	--14512
		x"ff",	--14513
		x"ff",	--14514
		x"ff",	--14515
		x"ff",	--14516
		x"ff",	--14517
		x"ff",	--14518
		x"ff",	--14519
		x"ff",	--14520
		x"ff",	--14521
		x"ff",	--14522
		x"ff",	--14523
		x"ff",	--14524
		x"ff",	--14525
		x"ff",	--14526
		x"ff",	--14527
		x"ff",	--14528
		x"ff",	--14529
		x"ff",	--14530
		x"ff",	--14531
		x"ff",	--14532
		x"ff",	--14533
		x"ff",	--14534
		x"ff",	--14535
		x"ff",	--14536
		x"ff",	--14537
		x"ff",	--14538
		x"ff",	--14539
		x"ff",	--14540
		x"ff",	--14541
		x"ff",	--14542
		x"ff",	--14543
		x"ff",	--14544
		x"ff",	--14545
		x"ff",	--14546
		x"ff",	--14547
		x"ff",	--14548
		x"ff",	--14549
		x"ff",	--14550
		x"ff",	--14551
		x"ff",	--14552
		x"ff",	--14553
		x"ff",	--14554
		x"ff",	--14555
		x"ff",	--14556
		x"ff",	--14557
		x"ff",	--14558
		x"ff",	--14559
		x"ff",	--14560
		x"ff",	--14561
		x"ff",	--14562
		x"ff",	--14563
		x"ff",	--14564
		x"ff",	--14565
		x"ff",	--14566
		x"ff",	--14567
		x"ff",	--14568
		x"ff",	--14569
		x"ff",	--14570
		x"ff",	--14571
		x"ff",	--14572
		x"ff",	--14573
		x"ff",	--14574
		x"ff",	--14575
		x"ff",	--14576
		x"ff",	--14577
		x"ff",	--14578
		x"ff",	--14579
		x"ff",	--14580
		x"ff",	--14581
		x"ff",	--14582
		x"ff",	--14583
		x"ff",	--14584
		x"ff",	--14585
		x"ff",	--14586
		x"ff",	--14587
		x"ff",	--14588
		x"ff",	--14589
		x"ff",	--14590
		x"ff",	--14591
		x"ff",	--14592
		x"ff",	--14593
		x"ff",	--14594
		x"ff",	--14595
		x"ff",	--14596
		x"ff",	--14597
		x"ff",	--14598
		x"ff",	--14599
		x"ff",	--14600
		x"ff",	--14601
		x"ff",	--14602
		x"ff",	--14603
		x"ff",	--14604
		x"ff",	--14605
		x"ff",	--14606
		x"ff",	--14607
		x"ff",	--14608
		x"ff",	--14609
		x"ff",	--14610
		x"ff",	--14611
		x"ff",	--14612
		x"ff",	--14613
		x"ff",	--14614
		x"ff",	--14615
		x"ff",	--14616
		x"ff",	--14617
		x"ff",	--14618
		x"ff",	--14619
		x"ff",	--14620
		x"ff",	--14621
		x"ff",	--14622
		x"ff",	--14623
		x"ff",	--14624
		x"ff",	--14625
		x"ff",	--14626
		x"ff",	--14627
		x"ff",	--14628
		x"ff",	--14629
		x"ff",	--14630
		x"ff",	--14631
		x"ff",	--14632
		x"ff",	--14633
		x"ff",	--14634
		x"ff",	--14635
		x"ff",	--14636
		x"ff",	--14637
		x"ff",	--14638
		x"ff",	--14639
		x"ff",	--14640
		x"ff",	--14641
		x"ff",	--14642
		x"ff",	--14643
		x"ff",	--14644
		x"ff",	--14645
		x"ff",	--14646
		x"ff",	--14647
		x"ff",	--14648
		x"ff",	--14649
		x"ff",	--14650
		x"ff",	--14651
		x"ff",	--14652
		x"ff",	--14653
		x"ff",	--14654
		x"ff",	--14655
		x"ff",	--14656
		x"ff",	--14657
		x"ff",	--14658
		x"ff",	--14659
		x"ff",	--14660
		x"ff",	--14661
		x"ff",	--14662
		x"ff",	--14663
		x"ff",	--14664
		x"ff",	--14665
		x"ff",	--14666
		x"ff",	--14667
		x"ff",	--14668
		x"ff",	--14669
		x"ff",	--14670
		x"ff",	--14671
		x"ff",	--14672
		x"ff",	--14673
		x"ff",	--14674
		x"ff",	--14675
		x"ff",	--14676
		x"ff",	--14677
		x"ff",	--14678
		x"ff",	--14679
		x"ff",	--14680
		x"ff",	--14681
		x"ff",	--14682
		x"ff",	--14683
		x"ff",	--14684
		x"ff",	--14685
		x"ff",	--14686
		x"ff",	--14687
		x"ff",	--14688
		x"ff",	--14689
		x"ff",	--14690
		x"ff",	--14691
		x"ff",	--14692
		x"ff",	--14693
		x"ff",	--14694
		x"ff",	--14695
		x"ff",	--14696
		x"ff",	--14697
		x"ff",	--14698
		x"ff",	--14699
		x"ff",	--14700
		x"ff",	--14701
		x"ff",	--14702
		x"ff",	--14703
		x"ff",	--14704
		x"ff",	--14705
		x"ff",	--14706
		x"ff",	--14707
		x"ff",	--14708
		x"ff",	--14709
		x"ff",	--14710
		x"ff",	--14711
		x"ff",	--14712
		x"ff",	--14713
		x"ff",	--14714
		x"ff",	--14715
		x"ff",	--14716
		x"ff",	--14717
		x"ff",	--14718
		x"ff",	--14719
		x"ff",	--14720
		x"ff",	--14721
		x"ff",	--14722
		x"ff",	--14723
		x"ff",	--14724
		x"ff",	--14725
		x"ff",	--14726
		x"ff",	--14727
		x"ff",	--14728
		x"ff",	--14729
		x"ff",	--14730
		x"ff",	--14731
		x"ff",	--14732
		x"ff",	--14733
		x"ff",	--14734
		x"ff",	--14735
		x"ff",	--14736
		x"ff",	--14737
		x"ff",	--14738
		x"ff",	--14739
		x"ff",	--14740
		x"ff",	--14741
		x"ff",	--14742
		x"ff",	--14743
		x"ff",	--14744
		x"ff",	--14745
		x"ff",	--14746
		x"ff",	--14747
		x"ff",	--14748
		x"ff",	--14749
		x"ff",	--14750
		x"ff",	--14751
		x"ff",	--14752
		x"ff",	--14753
		x"ff",	--14754
		x"ff",	--14755
		x"ff",	--14756
		x"ff",	--14757
		x"ff",	--14758
		x"ff",	--14759
		x"ff",	--14760
		x"ff",	--14761
		x"ff",	--14762
		x"ff",	--14763
		x"ff",	--14764
		x"ff",	--14765
		x"ff",	--14766
		x"ff",	--14767
		x"ff",	--14768
		x"ff",	--14769
		x"ff",	--14770
		x"ff",	--14771
		x"ff",	--14772
		x"ff",	--14773
		x"ff",	--14774
		x"ff",	--14775
		x"ff",	--14776
		x"ff",	--14777
		x"ff",	--14778
		x"ff",	--14779
		x"ff",	--14780
		x"ff",	--14781
		x"ff",	--14782
		x"ff",	--14783
		x"ff",	--14784
		x"ff",	--14785
		x"ff",	--14786
		x"ff",	--14787
		x"ff",	--14788
		x"ff",	--14789
		x"ff",	--14790
		x"ff",	--14791
		x"ff",	--14792
		x"ff",	--14793
		x"ff",	--14794
		x"ff",	--14795
		x"ff",	--14796
		x"ff",	--14797
		x"ff",	--14798
		x"ff",	--14799
		x"ff",	--14800
		x"ff",	--14801
		x"ff",	--14802
		x"ff",	--14803
		x"ff",	--14804
		x"ff",	--14805
		x"ff",	--14806
		x"ff",	--14807
		x"ff",	--14808
		x"ff",	--14809
		x"ff",	--14810
		x"ff",	--14811
		x"ff",	--14812
		x"ff",	--14813
		x"ff",	--14814
		x"ff",	--14815
		x"ff",	--14816
		x"ff",	--14817
		x"ff",	--14818
		x"ff",	--14819
		x"ff",	--14820
		x"ff",	--14821
		x"ff",	--14822
		x"ff",	--14823
		x"ff",	--14824
		x"ff",	--14825
		x"ff",	--14826
		x"ff",	--14827
		x"ff",	--14828
		x"ff",	--14829
		x"ff",	--14830
		x"ff",	--14831
		x"ff",	--14832
		x"ff",	--14833
		x"ff",	--14834
		x"ff",	--14835
		x"ff",	--14836
		x"ff",	--14837
		x"ff",	--14838
		x"ff",	--14839
		x"ff",	--14840
		x"ff",	--14841
		x"ff",	--14842
		x"ff",	--14843
		x"ff",	--14844
		x"ff",	--14845
		x"ff",	--14846
		x"ff",	--14847
		x"ff",	--14848
		x"ff",	--14849
		x"ff",	--14850
		x"ff",	--14851
		x"ff",	--14852
		x"ff",	--14853
		x"ff",	--14854
		x"ff",	--14855
		x"ff",	--14856
		x"ff",	--14857
		x"ff",	--14858
		x"ff",	--14859
		x"ff",	--14860
		x"ff",	--14861
		x"ff",	--14862
		x"ff",	--14863
		x"ff",	--14864
		x"ff",	--14865
		x"ff",	--14866
		x"ff",	--14867
		x"ff",	--14868
		x"ff",	--14869
		x"ff",	--14870
		x"ff",	--14871
		x"ff",	--14872
		x"ff",	--14873
		x"ff",	--14874
		x"ff",	--14875
		x"ff",	--14876
		x"ff",	--14877
		x"ff",	--14878
		x"ff",	--14879
		x"ff",	--14880
		x"ff",	--14881
		x"ff",	--14882
		x"ff",	--14883
		x"ff",	--14884
		x"ff",	--14885
		x"ff",	--14886
		x"ff",	--14887
		x"ff",	--14888
		x"ff",	--14889
		x"ff",	--14890
		x"ff",	--14891
		x"ff",	--14892
		x"ff",	--14893
		x"ff",	--14894
		x"ff",	--14895
		x"ff",	--14896
		x"ff",	--14897
		x"ff",	--14898
		x"ff",	--14899
		x"ff",	--14900
		x"ff",	--14901
		x"ff",	--14902
		x"ff",	--14903
		x"ff",	--14904
		x"ff",	--14905
		x"ff",	--14906
		x"ff",	--14907
		x"ff",	--14908
		x"ff",	--14909
		x"ff",	--14910
		x"ff",	--14911
		x"ff",	--14912
		x"ff",	--14913
		x"ff",	--14914
		x"ff",	--14915
		x"ff",	--14916
		x"ff",	--14917
		x"ff",	--14918
		x"ff",	--14919
		x"ff",	--14920
		x"ff",	--14921
		x"ff",	--14922
		x"ff",	--14923
		x"ff",	--14924
		x"ff",	--14925
		x"ff",	--14926
		x"ff",	--14927
		x"ff",	--14928
		x"ff",	--14929
		x"ff",	--14930
		x"ff",	--14931
		x"ff",	--14932
		x"ff",	--14933
		x"ff",	--14934
		x"ff",	--14935
		x"ff",	--14936
		x"ff",	--14937
		x"ff",	--14938
		x"ff",	--14939
		x"ff",	--14940
		x"ff",	--14941
		x"ff",	--14942
		x"ff",	--14943
		x"ff",	--14944
		x"ff",	--14945
		x"ff",	--14946
		x"ff",	--14947
		x"ff",	--14948
		x"ff",	--14949
		x"ff",	--14950
		x"ff",	--14951
		x"ff",	--14952
		x"ff",	--14953
		x"ff",	--14954
		x"ff",	--14955
		x"ff",	--14956
		x"ff",	--14957
		x"ff",	--14958
		x"ff",	--14959
		x"ff",	--14960
		x"ff",	--14961
		x"ff",	--14962
		x"ff",	--14963
		x"ff",	--14964
		x"ff",	--14965
		x"ff",	--14966
		x"ff",	--14967
		x"ff",	--14968
		x"ff",	--14969
		x"ff",	--14970
		x"ff",	--14971
		x"ff",	--14972
		x"ff",	--14973
		x"ff",	--14974
		x"ff",	--14975
		x"ff",	--14976
		x"ff",	--14977
		x"ff",	--14978
		x"ff",	--14979
		x"ff",	--14980
		x"ff",	--14981
		x"ff",	--14982
		x"ff",	--14983
		x"ff",	--14984
		x"ff",	--14985
		x"ff",	--14986
		x"ff",	--14987
		x"ff",	--14988
		x"ff",	--14989
		x"ff",	--14990
		x"ff",	--14991
		x"ff",	--14992
		x"ff",	--14993
		x"ff",	--14994
		x"ff",	--14995
		x"ff",	--14996
		x"ff",	--14997
		x"ff",	--14998
		x"ff",	--14999
		x"ff",	--15000
		x"ff",	--15001
		x"ff",	--15002
		x"ff",	--15003
		x"ff",	--15004
		x"ff",	--15005
		x"ff",	--15006
		x"ff",	--15007
		x"ff",	--15008
		x"ff",	--15009
		x"ff",	--15010
		x"ff",	--15011
		x"ff",	--15012
		x"ff",	--15013
		x"ff",	--15014
		x"ff",	--15015
		x"ff",	--15016
		x"ff",	--15017
		x"ff",	--15018
		x"ff",	--15019
		x"ff",	--15020
		x"ff",	--15021
		x"ff",	--15022
		x"ff",	--15023
		x"ff",	--15024
		x"ff",	--15025
		x"ff",	--15026
		x"ff",	--15027
		x"ff",	--15028
		x"ff",	--15029
		x"ff",	--15030
		x"ff",	--15031
		x"ff",	--15032
		x"ff",	--15033
		x"ff",	--15034
		x"ff",	--15035
		x"ff",	--15036
		x"ff",	--15037
		x"ff",	--15038
		x"ff",	--15039
		x"ff",	--15040
		x"ff",	--15041
		x"ff",	--15042
		x"ff",	--15043
		x"ff",	--15044
		x"ff",	--15045
		x"ff",	--15046
		x"ff",	--15047
		x"ff",	--15048
		x"ff",	--15049
		x"ff",	--15050
		x"ff",	--15051
		x"ff",	--15052
		x"ff",	--15053
		x"ff",	--15054
		x"ff",	--15055
		x"ff",	--15056
		x"ff",	--15057
		x"ff",	--15058
		x"ff",	--15059
		x"ff",	--15060
		x"ff",	--15061
		x"ff",	--15062
		x"ff",	--15063
		x"ff",	--15064
		x"ff",	--15065
		x"ff",	--15066
		x"ff",	--15067
		x"ff",	--15068
		x"ff",	--15069
		x"ff",	--15070
		x"ff",	--15071
		x"ff",	--15072
		x"ff",	--15073
		x"ff",	--15074
		x"ff",	--15075
		x"ff",	--15076
		x"ff",	--15077
		x"ff",	--15078
		x"ff",	--15079
		x"ff",	--15080
		x"ff",	--15081
		x"ff",	--15082
		x"ff",	--15083
		x"ff",	--15084
		x"ff",	--15085
		x"ff",	--15086
		x"ff",	--15087
		x"ff",	--15088
		x"ff",	--15089
		x"ff",	--15090
		x"ff",	--15091
		x"ff",	--15092
		x"ff",	--15093
		x"ff",	--15094
		x"ff",	--15095
		x"ff",	--15096
		x"ff",	--15097
		x"ff",	--15098
		x"ff",	--15099
		x"ff",	--15100
		x"ff",	--15101
		x"ff",	--15102
		x"ff",	--15103
		x"ff",	--15104
		x"ff",	--15105
		x"ff",	--15106
		x"ff",	--15107
		x"ff",	--15108
		x"ff",	--15109
		x"ff",	--15110
		x"ff",	--15111
		x"ff",	--15112
		x"ff",	--15113
		x"ff",	--15114
		x"ff",	--15115
		x"ff",	--15116
		x"ff",	--15117
		x"ff",	--15118
		x"ff",	--15119
		x"ff",	--15120
		x"ff",	--15121
		x"ff",	--15122
		x"ff",	--15123
		x"ff",	--15124
		x"ff",	--15125
		x"ff",	--15126
		x"ff",	--15127
		x"ff",	--15128
		x"ff",	--15129
		x"ff",	--15130
		x"ff",	--15131
		x"ff",	--15132
		x"ff",	--15133
		x"ff",	--15134
		x"ff",	--15135
		x"ff",	--15136
		x"ff",	--15137
		x"ff",	--15138
		x"ff",	--15139
		x"ff",	--15140
		x"ff",	--15141
		x"ff",	--15142
		x"ff",	--15143
		x"ff",	--15144
		x"ff",	--15145
		x"ff",	--15146
		x"ff",	--15147
		x"ff",	--15148
		x"ff",	--15149
		x"ff",	--15150
		x"ff",	--15151
		x"ff",	--15152
		x"ff",	--15153
		x"ff",	--15154
		x"ff",	--15155
		x"ff",	--15156
		x"ff",	--15157
		x"ff",	--15158
		x"ff",	--15159
		x"ff",	--15160
		x"ff",	--15161
		x"ff",	--15162
		x"ff",	--15163
		x"ff",	--15164
		x"ff",	--15165
		x"ff",	--15166
		x"ff",	--15167
		x"ff",	--15168
		x"ff",	--15169
		x"ff",	--15170
		x"ff",	--15171
		x"ff",	--15172
		x"ff",	--15173
		x"ff",	--15174
		x"ff",	--15175
		x"ff",	--15176
		x"ff",	--15177
		x"ff",	--15178
		x"ff",	--15179
		x"ff",	--15180
		x"ff",	--15181
		x"ff",	--15182
		x"ff",	--15183
		x"ff",	--15184
		x"ff",	--15185
		x"ff",	--15186
		x"ff",	--15187
		x"ff",	--15188
		x"ff",	--15189
		x"ff",	--15190
		x"ff",	--15191
		x"ff",	--15192
		x"ff",	--15193
		x"ff",	--15194
		x"ff",	--15195
		x"ff",	--15196
		x"ff",	--15197
		x"ff",	--15198
		x"ff",	--15199
		x"ff",	--15200
		x"ff",	--15201
		x"ff",	--15202
		x"ff",	--15203
		x"ff",	--15204
		x"ff",	--15205
		x"ff",	--15206
		x"ff",	--15207
		x"ff",	--15208
		x"ff",	--15209
		x"ff",	--15210
		x"ff",	--15211
		x"ff",	--15212
		x"ff",	--15213
		x"ff",	--15214
		x"ff",	--15215
		x"ff",	--15216
		x"ff",	--15217
		x"ff",	--15218
		x"ff",	--15219
		x"ff",	--15220
		x"ff",	--15221
		x"ff",	--15222
		x"ff",	--15223
		x"ff",	--15224
		x"ff",	--15225
		x"ff",	--15226
		x"ff",	--15227
		x"ff",	--15228
		x"ff",	--15229
		x"ff",	--15230
		x"ff",	--15231
		x"ff",	--15232
		x"ff",	--15233
		x"ff",	--15234
		x"ff",	--15235
		x"ff",	--15236
		x"ff",	--15237
		x"ff",	--15238
		x"ff",	--15239
		x"ff",	--15240
		x"ff",	--15241
		x"ff",	--15242
		x"ff",	--15243
		x"ff",	--15244
		x"ff",	--15245
		x"ff",	--15246
		x"ff",	--15247
		x"ff",	--15248
		x"ff",	--15249
		x"ff",	--15250
		x"ff",	--15251
		x"ff",	--15252
		x"ff",	--15253
		x"ff",	--15254
		x"ff",	--15255
		x"ff",	--15256
		x"ff",	--15257
		x"ff",	--15258
		x"ff",	--15259
		x"ff",	--15260
		x"ff",	--15261
		x"ff",	--15262
		x"ff",	--15263
		x"ff",	--15264
		x"ff",	--15265
		x"ff",	--15266
		x"ff",	--15267
		x"ff",	--15268
		x"ff",	--15269
		x"ff",	--15270
		x"ff",	--15271
		x"ff",	--15272
		x"ff",	--15273
		x"ff",	--15274
		x"ff",	--15275
		x"ff",	--15276
		x"ff",	--15277
		x"ff",	--15278
		x"ff",	--15279
		x"ff",	--15280
		x"ff",	--15281
		x"ff",	--15282
		x"ff",	--15283
		x"ff",	--15284
		x"ff",	--15285
		x"ff",	--15286
		x"ff",	--15287
		x"ff",	--15288
		x"ff",	--15289
		x"ff",	--15290
		x"ff",	--15291
		x"ff",	--15292
		x"ff",	--15293
		x"ff",	--15294
		x"ff",	--15295
		x"ff",	--15296
		x"ff",	--15297
		x"ff",	--15298
		x"ff",	--15299
		x"ff",	--15300
		x"ff",	--15301
		x"ff",	--15302
		x"ff",	--15303
		x"ff",	--15304
		x"ff",	--15305
		x"ff",	--15306
		x"ff",	--15307
		x"ff",	--15308
		x"ff",	--15309
		x"ff",	--15310
		x"ff",	--15311
		x"ff",	--15312
		x"ff",	--15313
		x"ff",	--15314
		x"ff",	--15315
		x"ff",	--15316
		x"ff",	--15317
		x"ff",	--15318
		x"ff",	--15319
		x"ff",	--15320
		x"ff",	--15321
		x"ff",	--15322
		x"ff",	--15323
		x"ff",	--15324
		x"ff",	--15325
		x"ff",	--15326
		x"ff",	--15327
		x"ff",	--15328
		x"ff",	--15329
		x"ff",	--15330
		x"ff",	--15331
		x"ff",	--15332
		x"ff",	--15333
		x"ff",	--15334
		x"ff",	--15335
		x"ff",	--15336
		x"ff",	--15337
		x"ff",	--15338
		x"ff",	--15339
		x"ff",	--15340
		x"ff",	--15341
		x"ff",	--15342
		x"ff",	--15343
		x"ff",	--15344
		x"ff",	--15345
		x"ff",	--15346
		x"ff",	--15347
		x"ff",	--15348
		x"ff",	--15349
		x"ff",	--15350
		x"ff",	--15351
		x"ff",	--15352
		x"ff",	--15353
		x"ff",	--15354
		x"ff",	--15355
		x"ff",	--15356
		x"ff",	--15357
		x"ff",	--15358
		x"ff",	--15359
		x"ff",	--15360
		x"ff",	--15361
		x"ff",	--15362
		x"ff",	--15363
		x"ff",	--15364
		x"ff",	--15365
		x"ff",	--15366
		x"ff",	--15367
		x"ff",	--15368
		x"ff",	--15369
		x"ff",	--15370
		x"ff",	--15371
		x"ff",	--15372
		x"ff",	--15373
		x"ff",	--15374
		x"ff",	--15375
		x"ff",	--15376
		x"ff",	--15377
		x"ff",	--15378
		x"ff",	--15379
		x"ff",	--15380
		x"ff",	--15381
		x"ff",	--15382
		x"ff",	--15383
		x"ff",	--15384
		x"ff",	--15385
		x"ff",	--15386
		x"ff",	--15387
		x"ff",	--15388
		x"ff",	--15389
		x"ff",	--15390
		x"ff",	--15391
		x"ff",	--15392
		x"ff",	--15393
		x"ff",	--15394
		x"ff",	--15395
		x"ff",	--15396
		x"ff",	--15397
		x"ff",	--15398
		x"ff",	--15399
		x"ff",	--15400
		x"ff",	--15401
		x"ff",	--15402
		x"ff",	--15403
		x"ff",	--15404
		x"ff",	--15405
		x"ff",	--15406
		x"ff",	--15407
		x"ff",	--15408
		x"ff",	--15409
		x"ff",	--15410
		x"ff",	--15411
		x"ff",	--15412
		x"ff",	--15413
		x"ff",	--15414
		x"ff",	--15415
		x"ff",	--15416
		x"ff",	--15417
		x"ff",	--15418
		x"ff",	--15419
		x"ff",	--15420
		x"ff",	--15421
		x"ff",	--15422
		x"ff",	--15423
		x"ff",	--15424
		x"ff",	--15425
		x"ff",	--15426
		x"ff",	--15427
		x"ff",	--15428
		x"ff",	--15429
		x"ff",	--15430
		x"ff",	--15431
		x"ff",	--15432
		x"ff",	--15433
		x"ff",	--15434
		x"ff",	--15435
		x"ff",	--15436
		x"ff",	--15437
		x"ff",	--15438
		x"ff",	--15439
		x"ff",	--15440
		x"ff",	--15441
		x"ff",	--15442
		x"ff",	--15443
		x"ff",	--15444
		x"ff",	--15445
		x"ff",	--15446
		x"ff",	--15447
		x"ff",	--15448
		x"ff",	--15449
		x"ff",	--15450
		x"ff",	--15451
		x"ff",	--15452
		x"ff",	--15453
		x"ff",	--15454
		x"ff",	--15455
		x"ff",	--15456
		x"ff",	--15457
		x"ff",	--15458
		x"ff",	--15459
		x"ff",	--15460
		x"ff",	--15461
		x"ff",	--15462
		x"ff",	--15463
		x"ff",	--15464
		x"ff",	--15465
		x"ff",	--15466
		x"ff",	--15467
		x"ff",	--15468
		x"ff",	--15469
		x"ff",	--15470
		x"ff",	--15471
		x"ff",	--15472
		x"ff",	--15473
		x"ff",	--15474
		x"ff",	--15475
		x"ff",	--15476
		x"ff",	--15477
		x"ff",	--15478
		x"ff",	--15479
		x"ff",	--15480
		x"ff",	--15481
		x"ff",	--15482
		x"ff",	--15483
		x"ff",	--15484
		x"ff",	--15485
		x"ff",	--15486
		x"ff",	--15487
		x"ff",	--15488
		x"ff",	--15489
		x"ff",	--15490
		x"ff",	--15491
		x"ff",	--15492
		x"ff",	--15493
		x"ff",	--15494
		x"ff",	--15495
		x"ff",	--15496
		x"ff",	--15497
		x"ff",	--15498
		x"ff",	--15499
		x"ff",	--15500
		x"ff",	--15501
		x"ff",	--15502
		x"ff",	--15503
		x"ff",	--15504
		x"ff",	--15505
		x"ff",	--15506
		x"ff",	--15507
		x"ff",	--15508
		x"ff",	--15509
		x"ff",	--15510
		x"ff",	--15511
		x"ff",	--15512
		x"ff",	--15513
		x"ff",	--15514
		x"ff",	--15515
		x"ff",	--15516
		x"ff",	--15517
		x"ff",	--15518
		x"ff",	--15519
		x"ff",	--15520
		x"ff",	--15521
		x"ff",	--15522
		x"ff",	--15523
		x"ff",	--15524
		x"ff",	--15525
		x"ff",	--15526
		x"ff",	--15527
		x"ff",	--15528
		x"ff",	--15529
		x"ff",	--15530
		x"ff",	--15531
		x"ff",	--15532
		x"ff",	--15533
		x"ff",	--15534
		x"ff",	--15535
		x"ff",	--15536
		x"ff",	--15537
		x"ff",	--15538
		x"ff",	--15539
		x"ff",	--15540
		x"ff",	--15541
		x"ff",	--15542
		x"ff",	--15543
		x"ff",	--15544
		x"ff",	--15545
		x"ff",	--15546
		x"ff",	--15547
		x"ff",	--15548
		x"ff",	--15549
		x"ff",	--15550
		x"ff",	--15551
		x"ff",	--15552
		x"ff",	--15553
		x"ff",	--15554
		x"ff",	--15555
		x"ff",	--15556
		x"ff",	--15557
		x"ff",	--15558
		x"ff",	--15559
		x"ff",	--15560
		x"ff",	--15561
		x"ff",	--15562
		x"ff",	--15563
		x"ff",	--15564
		x"ff",	--15565
		x"ff",	--15566
		x"ff",	--15567
		x"ff",	--15568
		x"ff",	--15569
		x"ff",	--15570
		x"ff",	--15571
		x"ff",	--15572
		x"ff",	--15573
		x"ff",	--15574
		x"ff",	--15575
		x"ff",	--15576
		x"ff",	--15577
		x"ff",	--15578
		x"ff",	--15579
		x"ff",	--15580
		x"ff",	--15581
		x"ff",	--15582
		x"ff",	--15583
		x"ff",	--15584
		x"ff",	--15585
		x"ff",	--15586
		x"ff",	--15587
		x"ff",	--15588
		x"ff",	--15589
		x"ff",	--15590
		x"ff",	--15591
		x"ff",	--15592
		x"ff",	--15593
		x"ff",	--15594
		x"ff",	--15595
		x"ff",	--15596
		x"ff",	--15597
		x"ff",	--15598
		x"ff",	--15599
		x"ff",	--15600
		x"ff",	--15601
		x"ff",	--15602
		x"ff",	--15603
		x"ff",	--15604
		x"ff",	--15605
		x"ff",	--15606
		x"ff",	--15607
		x"ff",	--15608
		x"ff",	--15609
		x"ff",	--15610
		x"ff",	--15611
		x"ff",	--15612
		x"ff",	--15613
		x"ff",	--15614
		x"ff",	--15615
		x"ff",	--15616
		x"ff",	--15617
		x"ff",	--15618
		x"ff",	--15619
		x"ff",	--15620
		x"ff",	--15621
		x"ff",	--15622
		x"ff",	--15623
		x"ff",	--15624
		x"ff",	--15625
		x"ff",	--15626
		x"ff",	--15627
		x"ff",	--15628
		x"ff",	--15629
		x"ff",	--15630
		x"ff",	--15631
		x"ff",	--15632
		x"ff",	--15633
		x"ff",	--15634
		x"ff",	--15635
		x"ff",	--15636
		x"ff",	--15637
		x"ff",	--15638
		x"ff",	--15639
		x"ff",	--15640
		x"ff",	--15641
		x"ff",	--15642
		x"ff",	--15643
		x"ff",	--15644
		x"ff",	--15645
		x"ff",	--15646
		x"ff",	--15647
		x"ff",	--15648
		x"ff",	--15649
		x"ff",	--15650
		x"ff",	--15651
		x"ff",	--15652
		x"ff",	--15653
		x"ff",	--15654
		x"ff",	--15655
		x"ff",	--15656
		x"ff",	--15657
		x"ff",	--15658
		x"ff",	--15659
		x"ff",	--15660
		x"ff",	--15661
		x"ff",	--15662
		x"ff",	--15663
		x"ff",	--15664
		x"ff",	--15665
		x"ff",	--15666
		x"ff",	--15667
		x"ff",	--15668
		x"ff",	--15669
		x"ff",	--15670
		x"ff",	--15671
		x"ff",	--15672
		x"ff",	--15673
		x"ff",	--15674
		x"ff",	--15675
		x"ff",	--15676
		x"ff",	--15677
		x"ff",	--15678
		x"ff",	--15679
		x"ff",	--15680
		x"ff",	--15681
		x"ff",	--15682
		x"ff",	--15683
		x"ff",	--15684
		x"ff",	--15685
		x"ff",	--15686
		x"ff",	--15687
		x"ff",	--15688
		x"ff",	--15689
		x"ff",	--15690
		x"ff",	--15691
		x"ff",	--15692
		x"ff",	--15693
		x"ff",	--15694
		x"ff",	--15695
		x"ff",	--15696
		x"ff",	--15697
		x"ff",	--15698
		x"ff",	--15699
		x"ff",	--15700
		x"ff",	--15701
		x"ff",	--15702
		x"ff",	--15703
		x"ff",	--15704
		x"ff",	--15705
		x"ff",	--15706
		x"ff",	--15707
		x"ff",	--15708
		x"ff",	--15709
		x"ff",	--15710
		x"ff",	--15711
		x"ff",	--15712
		x"ff",	--15713
		x"ff",	--15714
		x"ff",	--15715
		x"ff",	--15716
		x"ff",	--15717
		x"ff",	--15718
		x"ff",	--15719
		x"ff",	--15720
		x"ff",	--15721
		x"ff",	--15722
		x"ff",	--15723
		x"ff",	--15724
		x"ff",	--15725
		x"ff",	--15726
		x"ff",	--15727
		x"ff",	--15728
		x"ff",	--15729
		x"ff",	--15730
		x"ff",	--15731
		x"ff",	--15732
		x"ff",	--15733
		x"ff",	--15734
		x"ff",	--15735
		x"ff",	--15736
		x"ff",	--15737
		x"ff",	--15738
		x"ff",	--15739
		x"ff",	--15740
		x"ff",	--15741
		x"ff",	--15742
		x"ff",	--15743
		x"ff",	--15744
		x"ff",	--15745
		x"ff",	--15746
		x"ff",	--15747
		x"ff",	--15748
		x"ff",	--15749
		x"ff",	--15750
		x"ff",	--15751
		x"ff",	--15752
		x"ff",	--15753
		x"ff",	--15754
		x"ff",	--15755
		x"ff",	--15756
		x"ff",	--15757
		x"ff",	--15758
		x"ff",	--15759
		x"ff",	--15760
		x"ff",	--15761
		x"ff",	--15762
		x"ff",	--15763
		x"ff",	--15764
		x"ff",	--15765
		x"ff",	--15766
		x"ff",	--15767
		x"ff",	--15768
		x"ff",	--15769
		x"ff",	--15770
		x"ff",	--15771
		x"ff",	--15772
		x"ff",	--15773
		x"ff",	--15774
		x"ff",	--15775
		x"ff",	--15776
		x"ff",	--15777
		x"ff",	--15778
		x"ff",	--15779
		x"ff",	--15780
		x"ff",	--15781
		x"ff",	--15782
		x"ff",	--15783
		x"ff",	--15784
		x"ff",	--15785
		x"ff",	--15786
		x"ff",	--15787
		x"ff",	--15788
		x"ff",	--15789
		x"ff",	--15790
		x"ff",	--15791
		x"ff",	--15792
		x"ff",	--15793
		x"ff",	--15794
		x"ff",	--15795
		x"ff",	--15796
		x"ff",	--15797
		x"ff",	--15798
		x"ff",	--15799
		x"ff",	--15800
		x"ff",	--15801
		x"ff",	--15802
		x"ff",	--15803
		x"ff",	--15804
		x"ff",	--15805
		x"ff",	--15806
		x"ff",	--15807
		x"ff",	--15808
		x"ff",	--15809
		x"ff",	--15810
		x"ff",	--15811
		x"ff",	--15812
		x"ff",	--15813
		x"ff",	--15814
		x"ff",	--15815
		x"ff",	--15816
		x"ff",	--15817
		x"ff",	--15818
		x"ff",	--15819
		x"ff",	--15820
		x"ff",	--15821
		x"ff",	--15822
		x"ff",	--15823
		x"ff",	--15824
		x"ff",	--15825
		x"ff",	--15826
		x"ff",	--15827
		x"ff",	--15828
		x"ff",	--15829
		x"ff",	--15830
		x"ff",	--15831
		x"ff",	--15832
		x"ff",	--15833
		x"ff",	--15834
		x"ff",	--15835
		x"ff",	--15836
		x"ff",	--15837
		x"ff",	--15838
		x"ff",	--15839
		x"ff",	--15840
		x"ff",	--15841
		x"ff",	--15842
		x"ff",	--15843
		x"ff",	--15844
		x"ff",	--15845
		x"ff",	--15846
		x"ff",	--15847
		x"ff",	--15848
		x"ff",	--15849
		x"ff",	--15850
		x"ff",	--15851
		x"ff",	--15852
		x"ff",	--15853
		x"ff",	--15854
		x"ff",	--15855
		x"ff",	--15856
		x"ff",	--15857
		x"ff",	--15858
		x"ff",	--15859
		x"ff",	--15860
		x"ff",	--15861
		x"ff",	--15862
		x"ff",	--15863
		x"ff",	--15864
		x"ff",	--15865
		x"ff",	--15866
		x"ff",	--15867
		x"ff",	--15868
		x"ff",	--15869
		x"ff",	--15870
		x"ff",	--15871
		x"ff",	--15872
		x"ff",	--15873
		x"ff",	--15874
		x"ff",	--15875
		x"ff",	--15876
		x"ff",	--15877
		x"ff",	--15878
		x"ff",	--15879
		x"ff",	--15880
		x"ff",	--15881
		x"ff",	--15882
		x"ff",	--15883
		x"ff",	--15884
		x"ff",	--15885
		x"ff",	--15886
		x"ff",	--15887
		x"ff",	--15888
		x"ff",	--15889
		x"ff",	--15890
		x"ff",	--15891
		x"ff",	--15892
		x"ff",	--15893
		x"ff",	--15894
		x"ff",	--15895
		x"ff",	--15896
		x"ff",	--15897
		x"ff",	--15898
		x"ff",	--15899
		x"ff",	--15900
		x"ff",	--15901
		x"ff",	--15902
		x"ff",	--15903
		x"ff",	--15904
		x"ff",	--15905
		x"ff",	--15906
		x"ff",	--15907
		x"ff",	--15908
		x"ff",	--15909
		x"ff",	--15910
		x"ff",	--15911
		x"ff",	--15912
		x"ff",	--15913
		x"ff",	--15914
		x"ff",	--15915
		x"ff",	--15916
		x"ff",	--15917
		x"ff",	--15918
		x"ff",	--15919
		x"ff",	--15920
		x"ff",	--15921
		x"ff",	--15922
		x"ff",	--15923
		x"ff",	--15924
		x"ff",	--15925
		x"ff",	--15926
		x"ff",	--15927
		x"ff",	--15928
		x"ff",	--15929
		x"ff",	--15930
		x"ff",	--15931
		x"ff",	--15932
		x"ff",	--15933
		x"ff",	--15934
		x"ff",	--15935
		x"ff",	--15936
		x"ff",	--15937
		x"ff",	--15938
		x"ff",	--15939
		x"ff",	--15940
		x"ff",	--15941
		x"ff",	--15942
		x"ff",	--15943
		x"ff",	--15944
		x"ff",	--15945
		x"ff",	--15946
		x"ff",	--15947
		x"ff",	--15948
		x"ff",	--15949
		x"ff",	--15950
		x"ff",	--15951
		x"ff",	--15952
		x"ff",	--15953
		x"ff",	--15954
		x"ff",	--15955
		x"ff",	--15956
		x"ff",	--15957
		x"ff",	--15958
		x"ff",	--15959
		x"ff",	--15960
		x"ff",	--15961
		x"ff",	--15962
		x"ff",	--15963
		x"ff",	--15964
		x"ff",	--15965
		x"ff",	--15966
		x"ff",	--15967
		x"ff",	--15968
		x"ff",	--15969
		x"ff",	--15970
		x"ff",	--15971
		x"ff",	--15972
		x"ff",	--15973
		x"ff",	--15974
		x"ff",	--15975
		x"ff",	--15976
		x"ff",	--15977
		x"ff",	--15978
		x"ff",	--15979
		x"ff",	--15980
		x"ff",	--15981
		x"ff",	--15982
		x"ff",	--15983
		x"ff",	--15984
		x"ff",	--15985
		x"ff",	--15986
		x"ff",	--15987
		x"ff",	--15988
		x"ff",	--15989
		x"ff",	--15990
		x"ff",	--15991
		x"ff",	--15992
		x"ff",	--15993
		x"ff",	--15994
		x"ff",	--15995
		x"ff",	--15996
		x"ff",	--15997
		x"ff",	--15998
		x"ff",	--15999
		x"ff",	--16000
		x"ff",	--16001
		x"ff",	--16002
		x"ff",	--16003
		x"ff",	--16004
		x"ff",	--16005
		x"ff",	--16006
		x"ff",	--16007
		x"ff",	--16008
		x"ff",	--16009
		x"ff",	--16010
		x"ff",	--16011
		x"ff",	--16012
		x"ff",	--16013
		x"ff",	--16014
		x"ff",	--16015
		x"ff",	--16016
		x"ff",	--16017
		x"ff",	--16018
		x"ff",	--16019
		x"ff",	--16020
		x"ff",	--16021
		x"ff",	--16022
		x"ff",	--16023
		x"ff",	--16024
		x"ff",	--16025
		x"ff",	--16026
		x"ff",	--16027
		x"ff",	--16028
		x"ff",	--16029
		x"ff",	--16030
		x"ff",	--16031
		x"ff",	--16032
		x"ff",	--16033
		x"ff",	--16034
		x"ff",	--16035
		x"ff",	--16036
		x"ff",	--16037
		x"ff",	--16038
		x"ff",	--16039
		x"ff",	--16040
		x"ff",	--16041
		x"ff",	--16042
		x"ff",	--16043
		x"ff",	--16044
		x"ff",	--16045
		x"ff",	--16046
		x"ff",	--16047
		x"ff",	--16048
		x"ff",	--16049
		x"ff",	--16050
		x"ff",	--16051
		x"ff",	--16052
		x"ff",	--16053
		x"ff",	--16054
		x"ff",	--16055
		x"ff",	--16056
		x"ff",	--16057
		x"ff",	--16058
		x"ff",	--16059
		x"ff",	--16060
		x"ff",	--16061
		x"ff",	--16062
		x"ff",	--16063
		x"ff",	--16064
		x"ff",	--16065
		x"ff",	--16066
		x"ff",	--16067
		x"ff",	--16068
		x"ff",	--16069
		x"ff",	--16070
		x"ff",	--16071
		x"ff",	--16072
		x"ff",	--16073
		x"ff",	--16074
		x"ff",	--16075
		x"ff",	--16076
		x"ff",	--16077
		x"ff",	--16078
		x"ff",	--16079
		x"ff",	--16080
		x"ff",	--16081
		x"ff",	--16082
		x"ff",	--16083
		x"ff",	--16084
		x"ff",	--16085
		x"ff",	--16086
		x"ff",	--16087
		x"ff",	--16088
		x"ff",	--16089
		x"ff",	--16090
		x"ff",	--16091
		x"ff",	--16092
		x"ff",	--16093
		x"ff",	--16094
		x"ff",	--16095
		x"ff",	--16096
		x"ff",	--16097
		x"ff",	--16098
		x"ff",	--16099
		x"ff",	--16100
		x"ff",	--16101
		x"ff",	--16102
		x"ff",	--16103
		x"ff",	--16104
		x"ff",	--16105
		x"ff",	--16106
		x"ff",	--16107
		x"ff",	--16108
		x"ff",	--16109
		x"ff",	--16110
		x"ff",	--16111
		x"ff",	--16112
		x"ff",	--16113
		x"ff",	--16114
		x"ff",	--16115
		x"ff",	--16116
		x"ff",	--16117
		x"ff",	--16118
		x"ff",	--16119
		x"ff",	--16120
		x"ff",	--16121
		x"ff",	--16122
		x"ff",	--16123
		x"ff",	--16124
		x"ff",	--16125
		x"ff",	--16126
		x"ff",	--16127
		x"ff",	--16128
		x"ff",	--16129
		x"ff",	--16130
		x"ff",	--16131
		x"ff",	--16132
		x"ff",	--16133
		x"ff",	--16134
		x"ff",	--16135
		x"ff",	--16136
		x"ff",	--16137
		x"ff",	--16138
		x"ff",	--16139
		x"ff",	--16140
		x"ff",	--16141
		x"ff",	--16142
		x"ff",	--16143
		x"ff",	--16144
		x"ff",	--16145
		x"ff",	--16146
		x"ff",	--16147
		x"ff",	--16148
		x"ff",	--16149
		x"ff",	--16150
		x"ff",	--16151
		x"ff",	--16152
		x"ff",	--16153
		x"ff",	--16154
		x"ff",	--16155
		x"ff",	--16156
		x"ff",	--16157
		x"ff",	--16158
		x"ff",	--16159
		x"ff",	--16160
		x"ff",	--16161
		x"ff",	--16162
		x"ff",	--16163
		x"ff",	--16164
		x"ff",	--16165
		x"ff",	--16166
		x"ff",	--16167
		x"ff",	--16168
		x"ff",	--16169
		x"ff",	--16170
		x"ff",	--16171
		x"ff",	--16172
		x"ff",	--16173
		x"ff",	--16174
		x"ff",	--16175
		x"ff",	--16176
		x"ff",	--16177
		x"ff",	--16178
		x"ff",	--16179
		x"ff",	--16180
		x"ff",	--16181
		x"ff",	--16182
		x"ff",	--16183
		x"ff",	--16184
		x"ff",	--16185
		x"ff",	--16186
		x"ff",	--16187
		x"ff",	--16188
		x"ff",	--16189
		x"ff",	--16190
		x"ff",	--16191
		x"ff",	--16192
		x"ff",	--16193
		x"ff",	--16194
		x"ff",	--16195
		x"ff",	--16196
		x"ff",	--16197
		x"ff",	--16198
		x"ff",	--16199
		x"ff",	--16200
		x"ff",	--16201
		x"ff",	--16202
		x"ff",	--16203
		x"ff",	--16204
		x"ff",	--16205
		x"ff",	--16206
		x"ff",	--16207
		x"ff",	--16208
		x"ff",	--16209
		x"ff",	--16210
		x"ff",	--16211
		x"ff",	--16212
		x"ff",	--16213
		x"ff",	--16214
		x"ff",	--16215
		x"ff",	--16216
		x"ff",	--16217
		x"ff",	--16218
		x"ff",	--16219
		x"ff",	--16220
		x"ff",	--16221
		x"ff",	--16222
		x"ff",	--16223
		x"ff",	--16224
		x"ff",	--16225
		x"ff",	--16226
		x"ff",	--16227
		x"ff",	--16228
		x"ff",	--16229
		x"ff",	--16230
		x"ff",	--16231
		x"ff",	--16232
		x"ff",	--16233
		x"ff",	--16234
		x"ff",	--16235
		x"ff",	--16236
		x"ff",	--16237
		x"ff",	--16238
		x"ff",	--16239
		x"ff",	--16240
		x"ff",	--16241
		x"ff",	--16242
		x"ff",	--16243
		x"ff",	--16244
		x"ff",	--16245
		x"ff",	--16246
		x"ff",	--16247
		x"ff",	--16248
		x"ff",	--16249
		x"ff",	--16250
		x"ff",	--16251
		x"ff",	--16252
		x"ff",	--16253
		x"ff",	--16254
		x"ff",	--16255
		x"ff",	--16256
		x"ff",	--16257
		x"ff",	--16258
		x"ff",	--16259
		x"ff",	--16260
		x"ff",	--16261
		x"ff",	--16262
		x"ff",	--16263
		x"ff",	--16264
		x"ff",	--16265
		x"ff",	--16266
		x"ff",	--16267
		x"ff",	--16268
		x"ff",	--16269
		x"ff",	--16270
		x"ff",	--16271
		x"ff",	--16272
		x"ff",	--16273
		x"ff",	--16274
		x"ff",	--16275
		x"ff",	--16276
		x"ff",	--16277
		x"ff",	--16278
		x"ff",	--16279
		x"ff",	--16280
		x"ff",	--16281
		x"ff",	--16282
		x"ff",	--16283
		x"ff",	--16284
		x"ff",	--16285
		x"ff",	--16286
		x"ff",	--16287
		x"ff",	--16288
		x"ff",	--16289
		x"ff",	--16290
		x"ff",	--16291
		x"ff",	--16292
		x"ff",	--16293
		x"ff",	--16294
		x"ff",	--16295
		x"ff",	--16296
		x"ff",	--16297
		x"ff",	--16298
		x"ff",	--16299
		x"ff",	--16300
		x"ff",	--16301
		x"ff",	--16302
		x"ff",	--16303
		x"ff",	--16304
		x"ff",	--16305
		x"ff",	--16306
		x"ff",	--16307
		x"ff",	--16308
		x"ff",	--16309
		x"ff",	--16310
		x"ff",	--16311
		x"ff",	--16312
		x"ff",	--16313
		x"ff",	--16314
		x"ff",	--16315
		x"ff",	--16316
		x"ff",	--16317
		x"ff",	--16318
		x"ff",	--16319
		x"ff",	--16320
		x"ff",	--16321
		x"ff",	--16322
		x"ff",	--16323
		x"ff",	--16324
		x"ff",	--16325
		x"ff",	--16326
		x"ff",	--16327
		x"ff",	--16328
		x"ff",	--16329
		x"ff",	--16330
		x"ff",	--16331
		x"ff",	--16332
		x"ff",	--16333
		x"ff",	--16334
		x"ff",	--16335
		x"ff",	--16336
		x"ff",	--16337
		x"ff",	--16338
		x"ff",	--16339
		x"ff",	--16340
		x"ff",	--16341
		x"ff",	--16342
		x"ff",	--16343
		x"ff",	--16344
		x"ff",	--16345
		x"ff",	--16346
		x"ff",	--16347
		x"ff",	--16348
		x"ff",	--16349
		x"ff",	--16350
		x"ff",	--16351
		x"ff",	--16352
		x"ff",	--16353
		x"ff",	--16354
		x"ff",	--16355
		x"ff",	--16356
		x"ff",	--16357
		x"ff",	--16358
		x"ff",	--16359
		x"ff",	--16360
		x"ff",	--16361
		x"ff",	--16362
		x"ff",	--16363
		x"ff",	--16364
		x"ff",	--16365
		x"ff",	--16366
		x"ff",	--16367
		x"fc",	--16368
		x"fc",	--16369
		x"fc",	--16370
		x"fc",	--16371
		x"fc",	--16372
		x"fc",	--16373
		x"fc",	--16374
		x"32",	--16375
		x"84",	--16376
		x"fc",	--16377
		x"fc",	--16378
		x"fc",	--16379
		x"fc",	--16380
		x"fc",	--16381
		x"fc",	--16382
		x"00");	--16383
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"dd",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"9d",	--44
		x"12",	--45
		x"97",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"d4",	--50
		x"12",	--51
		x"9c",	--52
		x"53",	--53
		x"40",	--54
		x"d4",	--55
		x"40",	--56
		x"85",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"97",	--61
		x"40",	--62
		x"d4",	--63
		x"40",	--64
		x"91",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"97",	--69
		x"40",	--70
		x"d4",	--71
		x"40",	--72
		x"92",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"97",	--77
		x"40",	--78
		x"d4",	--79
		x"40",	--80
		x"85",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"97",	--85
		x"40",	--86
		x"d4",	--87
		x"40",	--88
		x"8a",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"97",	--93
		x"40",	--94
		x"d4",	--95
		x"40",	--96
		x"8b",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"97",	--101
		x"40",	--102
		x"d4",	--103
		x"40",	--104
		x"86",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"97",	--109
		x"40",	--110
		x"d4",	--111
		x"40",	--112
		x"84",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"97",	--117
		x"40",	--118
		x"d4",	--119
		x"40",	--120
		x"87",	--121
		x"40",	--122
		x"00",	--123
		x"12",	--124
		x"97",	--125
		x"40",	--126
		x"d5",	--127
		x"40",	--128
		x"84",	--129
		x"40",	--130
		x"00",	--131
		x"12",	--132
		x"97",	--133
		x"40",	--134
		x"d5",	--135
		x"40",	--136
		x"8f",	--137
		x"40",	--138
		x"00",	--139
		x"12",	--140
		x"97",	--141
		x"40",	--142
		x"d5",	--143
		x"40",	--144
		x"87",	--145
		x"40",	--146
		x"00",	--147
		x"12",	--148
		x"97",	--149
		x"43",	--150
		x"43",	--151
		x"12",	--152
		x"97",	--153
		x"43",	--154
		x"40",	--155
		x"4e",	--156
		x"40",	--157
		x"01",	--158
		x"41",	--159
		x"50",	--160
		x"00",	--161
		x"12",	--162
		x"96",	--163
		x"41",	--164
		x"50",	--165
		x"00",	--166
		x"12",	--167
		x"96",	--168
		x"43",	--169
		x"40",	--170
		x"4e",	--171
		x"40",	--172
		x"01",	--173
		x"41",	--174
		x"52",	--175
		x"12",	--176
		x"96",	--177
		x"41",	--178
		x"52",	--179
		x"12",	--180
		x"96",	--181
		x"41",	--182
		x"52",	--183
		x"41",	--184
		x"50",	--185
		x"00",	--186
		x"12",	--187
		x"8a",	--188
		x"40",	--189
		x"01",	--190
		x"41",	--191
		x"50",	--192
		x"00",	--193
		x"12",	--194
		x"9a",	--195
		x"40",	--196
		x"01",	--197
		x"41",	--198
		x"52",	--199
		x"12",	--200
		x"9a",	--201
		x"41",	--202
		x"52",	--203
		x"41",	--204
		x"50",	--205
		x"00",	--206
		x"12",	--207
		x"8b",	--208
		x"41",	--209
		x"52",	--210
		x"41",	--211
		x"50",	--212
		x"00",	--213
		x"12",	--214
		x"8b",	--215
		x"12",	--216
		x"98",	--217
		x"40",	--218
		x"01",	--219
		x"41",	--220
		x"53",	--221
		x"12",	--222
		x"9a",	--223
		x"41",	--224
		x"53",	--225
		x"12",	--226
		x"85",	--227
		x"40",	--228
		x"00",	--229
		x"40",	--230
		x"11",	--231
		x"41",	--232
		x"53",	--233
		x"12",	--234
		x"9a",	--235
		x"40",	--236
		x"01",	--237
		x"41",	--238
		x"12",	--239
		x"98",	--240
		x"41",	--241
		x"12",	--242
		x"84",	--243
		x"12",	--244
		x"40",	--245
		x"12",	--246
		x"12",	--247
		x"12",	--248
		x"12",	--249
		x"39",	--250
		x"12",	--251
		x"b7",	--252
		x"12",	--253
		x"3a",	--254
		x"12",	--255
		x"49",	--256
		x"40",	--257
		x"00",	--258
		x"41",	--259
		x"50",	--260
		x"00",	--261
		x"41",	--262
		x"50",	--263
		x"00",	--264
		x"41",	--265
		x"50",	--266
		x"00",	--267
		x"12",	--268
		x"89",	--269
		x"50",	--270
		x"00",	--271
		x"12",	--272
		x"40",	--273
		x"12",	--274
		x"12",	--275
		x"12",	--276
		x"12",	--277
		x"39",	--278
		x"12",	--279
		x"b7",	--280
		x"12",	--281
		x"3a",	--282
		x"12",	--283
		x"49",	--284
		x"40",	--285
		x"00",	--286
		x"41",	--287
		x"50",	--288
		x"00",	--289
		x"41",	--290
		x"50",	--291
		x"00",	--292
		x"41",	--293
		x"50",	--294
		x"00",	--295
		x"12",	--296
		x"89",	--297
		x"50",	--298
		x"00",	--299
		x"41",	--300
		x"50",	--301
		x"00",	--302
		x"41",	--303
		x"50",	--304
		x"00",	--305
		x"12",	--306
		x"86",	--307
		x"41",	--308
		x"12",	--309
		x"86",	--310
		x"12",	--311
		x"86",	--312
		x"12",	--313
		x"04",	--314
		x"12",	--315
		x"3e",	--316
		x"12",	--317
		x"99",	--318
		x"40",	--319
		x"c2",	--320
		x"40",	--321
		x"3d",	--322
		x"41",	--323
		x"50",	--324
		x"00",	--325
		x"12",	--326
		x"93",	--327
		x"50",	--328
		x"00",	--329
		x"41",	--330
		x"50",	--331
		x"00",	--332
		x"41",	--333
		x"52",	--334
		x"41",	--335
		x"50",	--336
		x"00",	--337
		x"12",	--338
		x"93",	--339
		x"40",	--340
		x"00",	--341
		x"41",	--342
		x"50",	--343
		x"00",	--344
		x"12",	--345
		x"96",	--346
		x"41",	--347
		x"50",	--348
		x"00",	--349
		x"12",	--350
		x"84",	--351
		x"41",	--352
		x"50",	--353
		x"00",	--354
		x"41",	--355
		x"50",	--356
		x"00",	--357
		x"12",	--358
		x"8f",	--359
		x"41",	--360
		x"12",	--361
		x"8f",	--362
		x"40",	--363
		x"00",	--364
		x"12",	--365
		x"8f",	--366
		x"40",	--367
		x"ff",	--368
		x"00",	--369
		x"d2",	--370
		x"43",	--371
		x"43",	--372
		x"3c",	--373
		x"43",	--374
		x"3c",	--375
		x"43",	--376
		x"3c",	--377
		x"43",	--378
		x"12",	--379
		x"9d",	--380
		x"93",	--381
		x"27",	--382
		x"12",	--383
		x"9d",	--384
		x"93",	--385
		x"20",	--386
		x"90",	--387
		x"00",	--388
		x"24",	--389
		x"90",	--390
		x"00",	--391
		x"27",	--392
		x"92",	--393
		x"20",	--394
		x"3c",	--395
		x"12",	--396
		x"d5",	--397
		x"12",	--398
		x"9c",	--399
		x"53",	--400
		x"40",	--401
		x"00",	--402
		x"51",	--403
		x"5f",	--404
		x"43",	--405
		x"00",	--406
		x"4f",	--407
		x"41",	--408
		x"00",	--409
		x"12",	--410
		x"98",	--411
		x"43",	--412
		x"3f",	--413
		x"93",	--414
		x"27",	--415
		x"53",	--416
		x"12",	--417
		x"d5",	--418
		x"12",	--419
		x"9c",	--420
		x"53",	--421
		x"3f",	--422
		x"90",	--423
		x"00",	--424
		x"2f",	--425
		x"93",	--426
		x"02",	--427
		x"24",	--428
		x"4f",	--429
		x"11",	--430
		x"12",	--431
		x"12",	--432
		x"d5",	--433
		x"4f",	--434
		x"00",	--435
		x"12",	--436
		x"9c",	--437
		x"52",	--438
		x"41",	--439
		x"00",	--440
		x"40",	--441
		x"00",	--442
		x"51",	--443
		x"5a",	--444
		x"4f",	--445
		x"00",	--446
		x"53",	--447
		x"3f",	--448
		x"93",	--449
		x"20",	--450
		x"90",	--451
		x"00",	--452
		x"23",	--453
		x"3f",	--454
		x"93",	--455
		x"23",	--456
		x"90",	--457
		x"00",	--458
		x"24",	--459
		x"90",	--460
		x"00",	--461
		x"34",	--462
		x"90",	--463
		x"00",	--464
		x"23",	--465
		x"3c",	--466
		x"90",	--467
		x"00",	--468
		x"24",	--469
		x"90",	--470
		x"00",	--471
		x"23",	--472
		x"3c",	--473
		x"12",	--474
		x"d5",	--475
		x"12",	--476
		x"9c",	--477
		x"53",	--478
		x"12",	--479
		x"86",	--480
		x"43",	--481
		x"3f",	--482
		x"12",	--483
		x"d5",	--484
		x"12",	--485
		x"9c",	--486
		x"53",	--487
		x"12",	--488
		x"87",	--489
		x"43",	--490
		x"3f",	--491
		x"12",	--492
		x"d5",	--493
		x"12",	--494
		x"9c",	--495
		x"53",	--496
		x"12",	--497
		x"87",	--498
		x"43",	--499
		x"3f",	--500
		x"12",	--501
		x"d5",	--502
		x"12",	--503
		x"9c",	--504
		x"53",	--505
		x"12",	--506
		x"87",	--507
		x"43",	--508
		x"3f",	--509
		x"40",	--510
		x"d4",	--511
		x"4f",	--512
		x"02",	--513
		x"41",	--514
		x"12",	--515
		x"12",	--516
		x"d4",	--517
		x"12",	--518
		x"9c",	--519
		x"53",	--520
		x"42",	--521
		x"02",	--522
		x"43",	--523
		x"40",	--524
		x"44",	--525
		x"4b",	--526
		x"00",	--527
		x"4b",	--528
		x"00",	--529
		x"12",	--530
		x"be",	--531
		x"12",	--532
		x"c4",	--533
		x"12",	--534
		x"43",	--535
		x"40",	--536
		x"44",	--537
		x"4b",	--538
		x"00",	--539
		x"4b",	--540
		x"00",	--541
		x"12",	--542
		x"be",	--543
		x"12",	--544
		x"c4",	--545
		x"12",	--546
		x"43",	--547
		x"40",	--548
		x"44",	--549
		x"4b",	--550
		x"00",	--551
		x"4b",	--552
		x"00",	--553
		x"12",	--554
		x"be",	--555
		x"12",	--556
		x"c4",	--557
		x"12",	--558
		x"12",	--559
		x"d4",	--560
		x"12",	--561
		x"02",	--562
		x"12",	--563
		x"c9",	--564
		x"50",	--565
		x"00",	--566
		x"12",	--567
		x"02",	--568
		x"12",	--569
		x"d4",	--570
		x"12",	--571
		x"9c",	--572
		x"52",	--573
		x"43",	--574
		x"41",	--575
		x"41",	--576
		x"12",	--577
		x"12",	--578
		x"d4",	--579
		x"12",	--580
		x"9c",	--581
		x"53",	--582
		x"43",	--583
		x"4b",	--584
		x"42",	--585
		x"02",	--586
		x"12",	--587
		x"98",	--588
		x"12",	--589
		x"12",	--590
		x"d4",	--591
		x"12",	--592
		x"9c",	--593
		x"52",	--594
		x"53",	--595
		x"90",	--596
		x"00",	--597
		x"23",	--598
		x"12",	--599
		x"d4",	--600
		x"12",	--601
		x"9c",	--602
		x"53",	--603
		x"41",	--604
		x"41",	--605
		x"4f",	--606
		x"02",	--607
		x"41",	--608
		x"12",	--609
		x"83",	--610
		x"4e",	--611
		x"43",	--612
		x"00",	--613
		x"93",	--614
		x"24",	--615
		x"93",	--616
		x"02",	--617
		x"24",	--618
		x"43",	--619
		x"02",	--620
		x"41",	--621
		x"4b",	--622
		x"00",	--623
		x"12",	--624
		x"87",	--625
		x"43",	--626
		x"4f",	--627
		x"42",	--628
		x"02",	--629
		x"12",	--630
		x"99",	--631
		x"43",	--632
		x"53",	--633
		x"41",	--634
		x"41",	--635
		x"93",	--636
		x"02",	--637
		x"24",	--638
		x"43",	--639
		x"02",	--640
		x"42",	--641
		x"02",	--642
		x"12",	--643
		x"99",	--644
		x"43",	--645
		x"53",	--646
		x"41",	--647
		x"41",	--648
		x"43",	--649
		x"12",	--650
		x"84",	--651
		x"43",	--652
		x"53",	--653
		x"41",	--654
		x"41",	--655
		x"43",	--656
		x"40",	--657
		x"84",	--658
		x"12",	--659
		x"99",	--660
		x"4f",	--661
		x"02",	--662
		x"3f",	--663
		x"4f",	--664
		x"02",	--665
		x"41",	--666
		x"12",	--667
		x"12",	--668
		x"82",	--669
		x"4f",	--670
		x"4e",	--671
		x"93",	--672
		x"38",	--673
		x"41",	--674
		x"4b",	--675
		x"00",	--676
		x"12",	--677
		x"87",	--678
		x"4f",	--679
		x"93",	--680
		x"24",	--681
		x"41",	--682
		x"4b",	--683
		x"00",	--684
		x"4d",	--685
		x"00",	--686
		x"12",	--687
		x"87",	--688
		x"4f",	--689
		x"41",	--690
		x"00",	--691
		x"42",	--692
		x"02",	--693
		x"12",	--694
		x"9a",	--695
		x"43",	--696
		x"52",	--697
		x"41",	--698
		x"41",	--699
		x"41",	--700
		x"40",	--701
		x"00",	--702
		x"40",	--703
		x"11",	--704
		x"3f",	--705
		x"40",	--706
		x"11",	--707
		x"3f",	--708
		x"43",	--709
		x"93",	--710
		x"02",	--711
		x"24",	--712
		x"43",	--713
		x"4f",	--714
		x"02",	--715
		x"43",	--716
		x"41",	--717
		x"42",	--718
		x"00",	--719
		x"4e",	--720
		x"be",	--721
		x"20",	--722
		x"df",	--723
		x"00",	--724
		x"41",	--725
		x"cf",	--726
		x"00",	--727
		x"41",	--728
		x"42",	--729
		x"02",	--730
		x"92",	--731
		x"2c",	--732
		x"4e",	--733
		x"5f",	--734
		x"4f",	--735
		x"d4",	--736
		x"43",	--737
		x"00",	--738
		x"90",	--739
		x"00",	--740
		x"38",	--741
		x"43",	--742
		x"02",	--743
		x"41",	--744
		x"53",	--745
		x"4e",	--746
		x"02",	--747
		x"41",	--748
		x"40",	--749
		x"00",	--750
		x"00",	--751
		x"3f",	--752
		x"40",	--753
		x"00",	--754
		x"00",	--755
		x"3f",	--756
		x"42",	--757
		x"00",	--758
		x"3f",	--759
		x"40",	--760
		x"00",	--761
		x"00",	--762
		x"3f",	--763
		x"40",	--764
		x"00",	--765
		x"00",	--766
		x"3f",	--767
		x"40",	--768
		x"00",	--769
		x"00",	--770
		x"3f",	--771
		x"40",	--772
		x"00",	--773
		x"00",	--774
		x"3f",	--775
		x"43",	--776
		x"42",	--777
		x"02",	--778
		x"12",	--779
		x"8a",	--780
		x"43",	--781
		x"42",	--782
		x"02",	--783
		x"12",	--784
		x"8a",	--785
		x"12",	--786
		x"d5",	--787
		x"12",	--788
		x"9c",	--789
		x"53",	--790
		x"41",	--791
		x"93",	--792
		x"02",	--793
		x"24",	--794
		x"42",	--795
		x"02",	--796
		x"12",	--797
		x"89",	--798
		x"42",	--799
		x"02",	--800
		x"12",	--801
		x"89",	--802
		x"41",	--803
		x"43",	--804
		x"40",	--805
		x"86",	--806
		x"12",	--807
		x"99",	--808
		x"4f",	--809
		x"02",	--810
		x"3f",	--811
		x"4f",	--812
		x"02",	--813
		x"4e",	--814
		x"02",	--815
		x"41",	--816
		x"4f",	--817
		x"02",	--818
		x"41",	--819
		x"12",	--820
		x"12",	--821
		x"83",	--822
		x"4e",	--823
		x"90",	--824
		x"00",	--825
		x"38",	--826
		x"20",	--827
		x"41",	--828
		x"4b",	--829
		x"00",	--830
		x"12",	--831
		x"88",	--832
		x"4f",	--833
		x"41",	--834
		x"4b",	--835
		x"00",	--836
		x"12",	--837
		x"88",	--838
		x"4f",	--839
		x"12",	--840
		x"12",	--841
		x"12",	--842
		x"d5",	--843
		x"12",	--844
		x"9c",	--845
		x"50",	--846
		x"00",	--847
		x"4a",	--848
		x"42",	--849
		x"02",	--850
		x"12",	--851
		x"8a",	--852
		x"4b",	--853
		x"42",	--854
		x"02",	--855
		x"12",	--856
		x"8a",	--857
		x"43",	--858
		x"53",	--859
		x"41",	--860
		x"41",	--861
		x"41",	--862
		x"41",	--863
		x"4b",	--864
		x"00",	--865
		x"12",	--866
		x"87",	--867
		x"43",	--868
		x"4f",	--869
		x"42",	--870
		x"02",	--871
		x"12",	--872
		x"99",	--873
		x"3f",	--874
		x"12",	--875
		x"d5",	--876
		x"12",	--877
		x"9c",	--878
		x"4b",	--879
		x"00",	--880
		x"12",	--881
		x"d5",	--882
		x"12",	--883
		x"9c",	--884
		x"52",	--885
		x"43",	--886
		x"3f",	--887
		x"40",	--888
		x"00",	--889
		x"42",	--890
		x"02",	--891
		x"12",	--892
		x"8a",	--893
		x"40",	--894
		x"ff",	--895
		x"42",	--896
		x"02",	--897
		x"12",	--898
		x"8a",	--899
		x"43",	--900
		x"40",	--901
		x"00",	--902
		x"42",	--903
		x"02",	--904
		x"12",	--905
		x"99",	--906
		x"41",	--907
		x"40",	--908
		x"ff",	--909
		x"42",	--910
		x"02",	--911
		x"12",	--912
		x"8a",	--913
		x"40",	--914
		x"00",	--915
		x"42",	--916
		x"02",	--917
		x"12",	--918
		x"8a",	--919
		x"43",	--920
		x"40",	--921
		x"00",	--922
		x"42",	--923
		x"02",	--924
		x"12",	--925
		x"99",	--926
		x"41",	--927
		x"40",	--928
		x"ff",	--929
		x"42",	--930
		x"02",	--931
		x"12",	--932
		x"8a",	--933
		x"40",	--934
		x"ff",	--935
		x"42",	--936
		x"02",	--937
		x"12",	--938
		x"8a",	--939
		x"43",	--940
		x"40",	--941
		x"00",	--942
		x"42",	--943
		x"02",	--944
		x"12",	--945
		x"99",	--946
		x"41",	--947
		x"40",	--948
		x"00",	--949
		x"42",	--950
		x"02",	--951
		x"12",	--952
		x"8a",	--953
		x"40",	--954
		x"00",	--955
		x"42",	--956
		x"02",	--957
		x"12",	--958
		x"8a",	--959
		x"43",	--960
		x"40",	--961
		x"00",	--962
		x"42",	--963
		x"02",	--964
		x"12",	--965
		x"99",	--966
		x"41",	--967
		x"12",	--968
		x"d5",	--969
		x"12",	--970
		x"9c",	--971
		x"53",	--972
		x"43",	--973
		x"41",	--974
		x"40",	--975
		x"80",	--976
		x"01",	--977
		x"40",	--978
		x"00",	--979
		x"01",	--980
		x"40",	--981
		x"02",	--982
		x"01",	--983
		x"12",	--984
		x"d5",	--985
		x"12",	--986
		x"9c",	--987
		x"43",	--988
		x"01",	--989
		x"40",	--990
		x"d5",	--991
		x"00",	--992
		x"12",	--993
		x"9c",	--994
		x"53",	--995
		x"43",	--996
		x"41",	--997
		x"12",	--998
		x"12",	--999
		x"43",	--1000
		x"00",	--1001
		x"4f",	--1002
		x"93",	--1003
		x"24",	--1004
		x"53",	--1005
		x"43",	--1006
		x"43",	--1007
		x"3c",	--1008
		x"90",	--1009
		x"00",	--1010
		x"2c",	--1011
		x"5c",	--1012
		x"5c",	--1013
		x"5c",	--1014
		x"5c",	--1015
		x"11",	--1016
		x"5d",	--1017
		x"50",	--1018
		x"ff",	--1019
		x"43",	--1020
		x"4f",	--1021
		x"93",	--1022
		x"24",	--1023
		x"90",	--1024
		x"00",	--1025
		x"24",	--1026
		x"4d",	--1027
		x"50",	--1028
		x"ff",	--1029
		x"93",	--1030
		x"23",	--1031
		x"90",	--1032
		x"00",	--1033
		x"2c",	--1034
		x"5c",	--1035
		x"4c",	--1036
		x"5b",	--1037
		x"5b",	--1038
		x"5b",	--1039
		x"11",	--1040
		x"5d",	--1041
		x"50",	--1042
		x"ff",	--1043
		x"4f",	--1044
		x"93",	--1045
		x"23",	--1046
		x"43",	--1047
		x"00",	--1048
		x"4c",	--1049
		x"41",	--1050
		x"41",	--1051
		x"41",	--1052
		x"43",	--1053
		x"3f",	--1054
		x"4d",	--1055
		x"50",	--1056
		x"ff",	--1057
		x"90",	--1058
		x"00",	--1059
		x"2c",	--1060
		x"5c",	--1061
		x"5c",	--1062
		x"5c",	--1063
		x"5c",	--1064
		x"11",	--1065
		x"5d",	--1066
		x"50",	--1067
		x"ff",	--1068
		x"43",	--1069
		x"3f",	--1070
		x"4d",	--1071
		x"50",	--1072
		x"ff",	--1073
		x"90",	--1074
		x"00",	--1075
		x"2c",	--1076
		x"5c",	--1077
		x"5c",	--1078
		x"5c",	--1079
		x"5c",	--1080
		x"11",	--1081
		x"5d",	--1082
		x"50",	--1083
		x"ff",	--1084
		x"43",	--1085
		x"3f",	--1086
		x"11",	--1087
		x"12",	--1088
		x"12",	--1089
		x"d5",	--1090
		x"12",	--1091
		x"9c",	--1092
		x"52",	--1093
		x"43",	--1094
		x"4c",	--1095
		x"41",	--1096
		x"41",	--1097
		x"41",	--1098
		x"43",	--1099
		x"3f",	--1100
		x"12",	--1101
		x"12",	--1102
		x"43",	--1103
		x"00",	--1104
		x"4f",	--1105
		x"93",	--1106
		x"24",	--1107
		x"53",	--1108
		x"43",	--1109
		x"43",	--1110
		x"3c",	--1111
		x"4b",	--1112
		x"50",	--1113
		x"ff",	--1114
		x"90",	--1115
		x"00",	--1116
		x"2c",	--1117
		x"5c",	--1118
		x"4c",	--1119
		x"5d",	--1120
		x"5d",	--1121
		x"5d",	--1122
		x"11",	--1123
		x"5b",	--1124
		x"50",	--1125
		x"ff",	--1126
		x"4f",	--1127
		x"93",	--1128
		x"24",	--1129
		x"90",	--1130
		x"00",	--1131
		x"23",	--1132
		x"43",	--1133
		x"4f",	--1134
		x"93",	--1135
		x"23",	--1136
		x"12",	--1137
		x"c2",	--1138
		x"43",	--1139
		x"4a",	--1140
		x"01",	--1141
		x"4c",	--1142
		x"01",	--1143
		x"42",	--1144
		x"01",	--1145
		x"41",	--1146
		x"43",	--1147
		x"00",	--1148
		x"41",	--1149
		x"41",	--1150
		x"41",	--1151
		x"11",	--1152
		x"12",	--1153
		x"12",	--1154
		x"d5",	--1155
		x"12",	--1156
		x"9c",	--1157
		x"52",	--1158
		x"43",	--1159
		x"41",	--1160
		x"41",	--1161
		x"41",	--1162
		x"43",	--1163
		x"3f",	--1164
		x"12",	--1165
		x"12",	--1166
		x"12",	--1167
		x"4f",	--1168
		x"4f",	--1169
		x"00",	--1170
		x"12",	--1171
		x"9a",	--1172
		x"4e",	--1173
		x"4f",	--1174
		x"89",	--1175
		x"00",	--1176
		x"79",	--1177
		x"00",	--1178
		x"12",	--1179
		x"c3",	--1180
		x"4a",	--1181
		x"00",	--1182
		x"4b",	--1183
		x"00",	--1184
		x"4e",	--1185
		x"4f",	--1186
		x"49",	--1187
		x"12",	--1188
		x"90",	--1189
		x"43",	--1190
		x"40",	--1191
		x"3f",	--1192
		x"12",	--1193
		x"bd",	--1194
		x"4e",	--1195
		x"4f",	--1196
		x"40",	--1197
		x"66",	--1198
		x"40",	--1199
		x"3f",	--1200
		x"12",	--1201
		x"c2",	--1202
		x"93",	--1203
		x"24",	--1204
		x"34",	--1205
		x"40",	--1206
		x"cc",	--1207
		x"40",	--1208
		x"3d",	--1209
		x"4a",	--1210
		x"4b",	--1211
		x"12",	--1212
		x"c2",	--1213
		x"93",	--1214
		x"34",	--1215
		x"40",	--1216
		x"cc",	--1217
		x"40",	--1218
		x"3d",	--1219
		x"4a",	--1220
		x"4b",	--1221
		x"49",	--1222
		x"00",	--1223
		x"12",	--1224
		x"97",	--1225
		x"41",	--1226
		x"41",	--1227
		x"41",	--1228
		x"41",	--1229
		x"40",	--1230
		x"66",	--1231
		x"40",	--1232
		x"3f",	--1233
		x"3f",	--1234
		x"12",	--1235
		x"12",	--1236
		x"4f",	--1237
		x"4c",	--1238
		x"4e",	--1239
		x"00",	--1240
		x"4d",	--1241
		x"00",	--1242
		x"12",	--1243
		x"00",	--1244
		x"12",	--1245
		x"00",	--1246
		x"12",	--1247
		x"00",	--1248
		x"12",	--1249
		x"00",	--1250
		x"12",	--1251
		x"00",	--1252
		x"12",	--1253
		x"00",	--1254
		x"41",	--1255
		x"00",	--1256
		x"41",	--1257
		x"00",	--1258
		x"12",	--1259
		x"90",	--1260
		x"50",	--1261
		x"00",	--1262
		x"4a",	--1263
		x"00",	--1264
		x"4b",	--1265
		x"40",	--1266
		x"89",	--1267
		x"12",	--1268
		x"99",	--1269
		x"4f",	--1270
		x"00",	--1271
		x"41",	--1272
		x"41",	--1273
		x"41",	--1274
		x"12",	--1275
		x"4f",	--1276
		x"4f",	--1277
		x"00",	--1278
		x"12",	--1279
		x"9a",	--1280
		x"4e",	--1281
		x"00",	--1282
		x"4f",	--1283
		x"00",	--1284
		x"43",	--1285
		x"4b",	--1286
		x"00",	--1287
		x"4b",	--1288
		x"00",	--1289
		x"12",	--1290
		x"99",	--1291
		x"41",	--1292
		x"41",	--1293
		x"12",	--1294
		x"4f",	--1295
		x"43",	--1296
		x"40",	--1297
		x"3f",	--1298
		x"4f",	--1299
		x"00",	--1300
		x"12",	--1301
		x"97",	--1302
		x"4b",	--1303
		x"00",	--1304
		x"12",	--1305
		x"99",	--1306
		x"41",	--1307
		x"41",	--1308
		x"12",	--1309
		x"4f",	--1310
		x"4e",	--1311
		x"10",	--1312
		x"11",	--1313
		x"10",	--1314
		x"11",	--1315
		x"4d",	--1316
		x"12",	--1317
		x"c3",	--1318
		x"4e",	--1319
		x"4f",	--1320
		x"4b",	--1321
		x"12",	--1322
		x"90",	--1323
		x"41",	--1324
		x"41",	--1325
		x"12",	--1326
		x"12",	--1327
		x"43",	--1328
		x"40",	--1329
		x"3f",	--1330
		x"4a",	--1331
		x"4b",	--1332
		x"42",	--1333
		x"02",	--1334
		x"12",	--1335
		x"97",	--1336
		x"4a",	--1337
		x"4b",	--1338
		x"42",	--1339
		x"02",	--1340
		x"12",	--1341
		x"97",	--1342
		x"12",	--1343
		x"d5",	--1344
		x"12",	--1345
		x"9c",	--1346
		x"53",	--1347
		x"41",	--1348
		x"41",	--1349
		x"41",	--1350
		x"4f",	--1351
		x"02",	--1352
		x"4e",	--1353
		x"02",	--1354
		x"41",	--1355
		x"12",	--1356
		x"12",	--1357
		x"83",	--1358
		x"4f",	--1359
		x"4e",	--1360
		x"93",	--1361
		x"02",	--1362
		x"24",	--1363
		x"90",	--1364
		x"00",	--1365
		x"38",	--1366
		x"20",	--1367
		x"41",	--1368
		x"4b",	--1369
		x"00",	--1370
		x"12",	--1371
		x"87",	--1372
		x"4f",	--1373
		x"41",	--1374
		x"4b",	--1375
		x"00",	--1376
		x"12",	--1377
		x"87",	--1378
		x"4f",	--1379
		x"12",	--1380
		x"12",	--1381
		x"12",	--1382
		x"d6",	--1383
		x"12",	--1384
		x"9c",	--1385
		x"50",	--1386
		x"00",	--1387
		x"4a",	--1388
		x"43",	--1389
		x"12",	--1390
		x"c4",	--1391
		x"43",	--1392
		x"40",	--1393
		x"42",	--1394
		x"12",	--1395
		x"c0",	--1396
		x"4e",	--1397
		x"4f",	--1398
		x"43",	--1399
		x"40",	--1400
		x"3f",	--1401
		x"12",	--1402
		x"be",	--1403
		x"4e",	--1404
		x"4f",	--1405
		x"42",	--1406
		x"02",	--1407
		x"12",	--1408
		x"97",	--1409
		x"4b",	--1410
		x"43",	--1411
		x"12",	--1412
		x"c4",	--1413
		x"43",	--1414
		x"40",	--1415
		x"42",	--1416
		x"12",	--1417
		x"c0",	--1418
		x"4e",	--1419
		x"4f",	--1420
		x"42",	--1421
		x"02",	--1422
		x"12",	--1423
		x"97",	--1424
		x"43",	--1425
		x"53",	--1426
		x"41",	--1427
		x"41",	--1428
		x"41",	--1429
		x"41",	--1430
		x"4b",	--1431
		x"00",	--1432
		x"12",	--1433
		x"87",	--1434
		x"43",	--1435
		x"4f",	--1436
		x"42",	--1437
		x"02",	--1438
		x"12",	--1439
		x"99",	--1440
		x"3f",	--1441
		x"43",	--1442
		x"40",	--1443
		x"8a",	--1444
		x"12",	--1445
		x"99",	--1446
		x"4f",	--1447
		x"02",	--1448
		x"3f",	--1449
		x"12",	--1450
		x"d5",	--1451
		x"12",	--1452
		x"9c",	--1453
		x"40",	--1454
		x"d6",	--1455
		x"00",	--1456
		x"12",	--1457
		x"9c",	--1458
		x"4b",	--1459
		x"00",	--1460
		x"12",	--1461
		x"d6",	--1462
		x"12",	--1463
		x"9c",	--1464
		x"52",	--1465
		x"43",	--1466
		x"3f",	--1467
		x"12",	--1468
		x"12",	--1469
		x"42",	--1470
		x"02",	--1471
		x"12",	--1472
		x"9a",	--1473
		x"4e",	--1474
		x"4f",	--1475
		x"42",	--1476
		x"02",	--1477
		x"12",	--1478
		x"9a",	--1479
		x"12",	--1480
		x"12",	--1481
		x"e3",	--1482
		x"e3",	--1483
		x"53",	--1484
		x"63",	--1485
		x"12",	--1486
		x"12",	--1487
		x"12",	--1488
		x"d6",	--1489
		x"12",	--1490
		x"02",	--1491
		x"12",	--1492
		x"c9",	--1493
		x"50",	--1494
		x"00",	--1495
		x"12",	--1496
		x"02",	--1497
		x"12",	--1498
		x"d6",	--1499
		x"12",	--1500
		x"9c",	--1501
		x"52",	--1502
		x"41",	--1503
		x"41",	--1504
		x"41",	--1505
		x"4f",	--1506
		x"02",	--1507
		x"4e",	--1508
		x"02",	--1509
		x"41",	--1510
		x"4f",	--1511
		x"02",	--1512
		x"4e",	--1513
		x"02",	--1514
		x"41",	--1515
		x"12",	--1516
		x"12",	--1517
		x"12",	--1518
		x"12",	--1519
		x"83",	--1520
		x"4f",	--1521
		x"4e",	--1522
		x"43",	--1523
		x"00",	--1524
		x"93",	--1525
		x"24",	--1526
		x"93",	--1527
		x"02",	--1528
		x"24",	--1529
		x"43",	--1530
		x"02",	--1531
		x"41",	--1532
		x"4b",	--1533
		x"00",	--1534
		x"12",	--1535
		x"87",	--1536
		x"4f",	--1537
		x"90",	--1538
		x"00",	--1539
		x"34",	--1540
		x"43",	--1541
		x"49",	--1542
		x"48",	--1543
		x"42",	--1544
		x"02",	--1545
		x"12",	--1546
		x"99",	--1547
		x"43",	--1548
		x"53",	--1549
		x"41",	--1550
		x"41",	--1551
		x"41",	--1552
		x"41",	--1553
		x"41",	--1554
		x"93",	--1555
		x"02",	--1556
		x"24",	--1557
		x"43",	--1558
		x"02",	--1559
		x"42",	--1560
		x"02",	--1561
		x"12",	--1562
		x"99",	--1563
		x"43",	--1564
		x"53",	--1565
		x"41",	--1566
		x"41",	--1567
		x"41",	--1568
		x"41",	--1569
		x"41",	--1570
		x"41",	--1571
		x"4b",	--1572
		x"00",	--1573
		x"12",	--1574
		x"87",	--1575
		x"4f",	--1576
		x"90",	--1577
		x"00",	--1578
		x"3b",	--1579
		x"41",	--1580
		x"4b",	--1581
		x"00",	--1582
		x"12",	--1583
		x"87",	--1584
		x"4f",	--1585
		x"41",	--1586
		x"4b",	--1587
		x"00",	--1588
		x"12",	--1589
		x"87",	--1590
		x"4f",	--1591
		x"12",	--1592
		x"12",	--1593
		x"12",	--1594
		x"d6",	--1595
		x"12",	--1596
		x"9c",	--1597
		x"50",	--1598
		x"00",	--1599
		x"4a",	--1600
		x"43",	--1601
		x"12",	--1602
		x"c4",	--1603
		x"43",	--1604
		x"40",	--1605
		x"42",	--1606
		x"12",	--1607
		x"c0",	--1608
		x"4e",	--1609
		x"4f",	--1610
		x"42",	--1611
		x"02",	--1612
		x"12",	--1613
		x"97",	--1614
		x"4b",	--1615
		x"43",	--1616
		x"12",	--1617
		x"c4",	--1618
		x"43",	--1619
		x"40",	--1620
		x"42",	--1621
		x"12",	--1622
		x"c0",	--1623
		x"4e",	--1624
		x"4f",	--1625
		x"42",	--1626
		x"02",	--1627
		x"12",	--1628
		x"97",	--1629
		x"3f",	--1630
		x"43",	--1631
		x"12",	--1632
		x"8b",	--1633
		x"43",	--1634
		x"53",	--1635
		x"41",	--1636
		x"41",	--1637
		x"41",	--1638
		x"41",	--1639
		x"41",	--1640
		x"43",	--1641
		x"40",	--1642
		x"8b",	--1643
		x"12",	--1644
		x"99",	--1645
		x"4f",	--1646
		x"02",	--1647
		x"3f",	--1648
		x"12",	--1649
		x"12",	--1650
		x"12",	--1651
		x"12",	--1652
		x"4f",	--1653
		x"40",	--1654
		x"d7",	--1655
		x"43",	--1656
		x"43",	--1657
		x"4b",	--1658
		x"48",	--1659
		x"12",	--1660
		x"98",	--1661
		x"9a",	--1662
		x"2c",	--1663
		x"43",	--1664
		x"4b",	--1665
		x"f0",	--1666
		x"00",	--1667
		x"24",	--1668
		x"5e",	--1669
		x"53",	--1670
		x"23",	--1671
		x"5e",	--1672
		x"53",	--1673
		x"53",	--1674
		x"90",	--1675
		x"00",	--1676
		x"23",	--1677
		x"49",	--1678
		x"41",	--1679
		x"41",	--1680
		x"41",	--1681
		x"41",	--1682
		x"41",	--1683
		x"12",	--1684
		x"12",	--1685
		x"93",	--1686
		x"02",	--1687
		x"20",	--1688
		x"41",	--1689
		x"41",	--1690
		x"41",	--1691
		x"42",	--1692
		x"02",	--1693
		x"12",	--1694
		x"8c",	--1695
		x"4f",	--1696
		x"43",	--1697
		x"4b",	--1698
		x"42",	--1699
		x"02",	--1700
		x"12",	--1701
		x"98",	--1702
		x"12",	--1703
		x"12",	--1704
		x"d6",	--1705
		x"12",	--1706
		x"9c",	--1707
		x"52",	--1708
		x"53",	--1709
		x"90",	--1710
		x"00",	--1711
		x"23",	--1712
		x"12",	--1713
		x"d6",	--1714
		x"12",	--1715
		x"9c",	--1716
		x"53",	--1717
		x"42",	--1718
		x"02",	--1719
		x"93",	--1720
		x"20",	--1721
		x"93",	--1722
		x"24",	--1723
		x"b2",	--1724
		x"20",	--1725
		x"b3",	--1726
		x"20",	--1727
		x"b3",	--1728
		x"20",	--1729
		x"b2",	--1730
		x"24",	--1731
		x"43",	--1732
		x"02",	--1733
		x"43",	--1734
		x"42",	--1735
		x"02",	--1736
		x"12",	--1737
		x"8a",	--1738
		x"43",	--1739
		x"42",	--1740
		x"02",	--1741
		x"12",	--1742
		x"8a",	--1743
		x"40",	--1744
		x"00",	--1745
		x"02",	--1746
		x"40",	--1747
		x"00",	--1748
		x"02",	--1749
		x"12",	--1750
		x"d6",	--1751
		x"12",	--1752
		x"9c",	--1753
		x"53",	--1754
		x"3f",	--1755
		x"93",	--1756
		x"02",	--1757
		x"20",	--1758
		x"42",	--1759
		x"02",	--1760
		x"93",	--1761
		x"24",	--1762
		x"93",	--1763
		x"24",	--1764
		x"93",	--1765
		x"24",	--1766
		x"90",	--1767
		x"00",	--1768
		x"24",	--1769
		x"53",	--1770
		x"4e",	--1771
		x"02",	--1772
		x"3f",	--1773
		x"43",	--1774
		x"02",	--1775
		x"3f",	--1776
		x"43",	--1777
		x"42",	--1778
		x"02",	--1779
		x"12",	--1780
		x"8a",	--1781
		x"43",	--1782
		x"42",	--1783
		x"02",	--1784
		x"12",	--1785
		x"8a",	--1786
		x"12",	--1787
		x"d6",	--1788
		x"12",	--1789
		x"9c",	--1790
		x"53",	--1791
		x"53",	--1792
		x"02",	--1793
		x"93",	--1794
		x"23",	--1795
		x"43",	--1796
		x"02",	--1797
		x"43",	--1798
		x"02",	--1799
		x"43",	--1800
		x"02",	--1801
		x"3f",	--1802
		x"43",	--1803
		x"42",	--1804
		x"02",	--1805
		x"12",	--1806
		x"8a",	--1807
		x"43",	--1808
		x"42",	--1809
		x"02",	--1810
		x"12",	--1811
		x"8a",	--1812
		x"12",	--1813
		x"12",	--1814
		x"d6",	--1815
		x"12",	--1816
		x"9c",	--1817
		x"52",	--1818
		x"3f",	--1819
		x"40",	--1820
		x"00",	--1821
		x"42",	--1822
		x"02",	--1823
		x"12",	--1824
		x"8a",	--1825
		x"40",	--1826
		x"00",	--1827
		x"42",	--1828
		x"02",	--1829
		x"12",	--1830
		x"8a",	--1831
		x"12",	--1832
		x"d6",	--1833
		x"12",	--1834
		x"9c",	--1835
		x"53",	--1836
		x"42",	--1837
		x"02",	--1838
		x"3f",	--1839
		x"40",	--1840
		x"00",	--1841
		x"42",	--1842
		x"02",	--1843
		x"12",	--1844
		x"8a",	--1845
		x"40",	--1846
		x"ff",	--1847
		x"42",	--1848
		x"02",	--1849
		x"12",	--1850
		x"8a",	--1851
		x"3f",	--1852
		x"12",	--1853
		x"d6",	--1854
		x"12",	--1855
		x"9c",	--1856
		x"53",	--1857
		x"3f",	--1858
		x"43",	--1859
		x"02",	--1860
		x"43",	--1861
		x"42",	--1862
		x"02",	--1863
		x"12",	--1864
		x"8a",	--1865
		x"43",	--1866
		x"42",	--1867
		x"02",	--1868
		x"12",	--1869
		x"8a",	--1870
		x"40",	--1871
		x"00",	--1872
		x"02",	--1873
		x"40",	--1874
		x"00",	--1875
		x"02",	--1876
		x"12",	--1877
		x"d6",	--1878
		x"12",	--1879
		x"9c",	--1880
		x"53",	--1881
		x"3f",	--1882
		x"40",	--1883
		x"00",	--1884
		x"02",	--1885
		x"43",	--1886
		x"42",	--1887
		x"02",	--1888
		x"12",	--1889
		x"8a",	--1890
		x"43",	--1891
		x"42",	--1892
		x"02",	--1893
		x"12",	--1894
		x"8a",	--1895
		x"40",	--1896
		x"00",	--1897
		x"02",	--1898
		x"40",	--1899
		x"00",	--1900
		x"02",	--1901
		x"12",	--1902
		x"d6",	--1903
		x"12",	--1904
		x"9c",	--1905
		x"53",	--1906
		x"3f",	--1907
		x"43",	--1908
		x"42",	--1909
		x"02",	--1910
		x"12",	--1911
		x"98",	--1912
		x"4f",	--1913
		x"43",	--1914
		x"42",	--1915
		x"02",	--1916
		x"12",	--1917
		x"98",	--1918
		x"9f",	--1919
		x"2c",	--1920
		x"40",	--1921
		x"00",	--1922
		x"42",	--1923
		x"02",	--1924
		x"12",	--1925
		x"8a",	--1926
		x"40",	--1927
		x"00",	--1928
		x"42",	--1929
		x"02",	--1930
		x"12",	--1931
		x"8a",	--1932
		x"12",	--1933
		x"d6",	--1934
		x"12",	--1935
		x"9c",	--1936
		x"53",	--1937
		x"42",	--1938
		x"02",	--1939
		x"3f",	--1940
		x"40",	--1941
		x"ff",	--1942
		x"42",	--1943
		x"02",	--1944
		x"12",	--1945
		x"8a",	--1946
		x"40",	--1947
		x"ff",	--1948
		x"42",	--1949
		x"02",	--1950
		x"12",	--1951
		x"8a",	--1952
		x"12",	--1953
		x"d6",	--1954
		x"12",	--1955
		x"9c",	--1956
		x"53",	--1957
		x"42",	--1958
		x"02",	--1959
		x"3f",	--1960
		x"40",	--1961
		x"ff",	--1962
		x"42",	--1963
		x"02",	--1964
		x"12",	--1965
		x"8a",	--1966
		x"40",	--1967
		x"ff",	--1968
		x"42",	--1969
		x"02",	--1970
		x"12",	--1971
		x"8a",	--1972
		x"3f",	--1973
		x"4f",	--1974
		x"02",	--1975
		x"4e",	--1976
		x"02",	--1977
		x"41",	--1978
		x"4f",	--1979
		x"02",	--1980
		x"41",	--1981
		x"12",	--1982
		x"4f",	--1983
		x"43",	--1984
		x"40",	--1985
		x"8d",	--1986
		x"12",	--1987
		x"99",	--1988
		x"4f",	--1989
		x"02",	--1990
		x"43",	--1991
		x"4b",	--1992
		x"12",	--1993
		x"99",	--1994
		x"41",	--1995
		x"41",	--1996
		x"12",	--1997
		x"4e",	--1998
		x"93",	--1999
		x"24",	--2000
		x"93",	--2001
		x"20",	--2002
		x"4e",	--2003
		x"00",	--2004
		x"4f",	--2005
		x"90",	--2006
		x"00",	--2007
		x"24",	--2008
		x"90",	--2009
		x"00",	--2010
		x"24",	--2011
		x"43",	--2012
		x"41",	--2013
		x"41",	--2014
		x"93",	--2015
		x"02",	--2016
		x"20",	--2017
		x"4f",	--2018
		x"02",	--2019
		x"93",	--2020
		x"24",	--2021
		x"12",	--2022
		x"d6",	--2023
		x"12",	--2024
		x"9c",	--2025
		x"53",	--2026
		x"43",	--2027
		x"41",	--2028
		x"41",	--2029
		x"43",	--2030
		x"42",	--2031
		x"02",	--2032
		x"12",	--2033
		x"8a",	--2034
		x"43",	--2035
		x"42",	--2036
		x"02",	--2037
		x"12",	--2038
		x"8a",	--2039
		x"12",	--2040
		x"d6",	--2041
		x"12",	--2042
		x"9c",	--2043
		x"53",	--2044
		x"43",	--2045
		x"41",	--2046
		x"41",	--2047
		x"43",	--2048
		x"4f",	--2049
		x"02",	--2050
		x"93",	--2051
		x"27",	--2052
		x"3f",	--2053
		x"43",	--2054
		x"02",	--2055
		x"3f",	--2056
		x"43",	--2057
		x"02",	--2058
		x"12",	--2059
		x"d6",	--2060
		x"12",	--2061
		x"9c",	--2062
		x"53",	--2063
		x"43",	--2064
		x"42",	--2065
		x"02",	--2066
		x"12",	--2067
		x"8a",	--2068
		x"43",	--2069
		x"42",	--2070
		x"02",	--2071
		x"12",	--2072
		x"8a",	--2073
		x"4b",	--2074
		x"00",	--2075
		x"4f",	--2076
		x"3f",	--2077
		x"4d",	--2078
		x"00",	--2079
		x"4e",	--2080
		x"00",	--2081
		x"41",	--2082
		x"00",	--2083
		x"00",	--2084
		x"41",	--2085
		x"00",	--2086
		x"00",	--2087
		x"41",	--2088
		x"00",	--2089
		x"00",	--2090
		x"41",	--2091
		x"00",	--2092
		x"00",	--2093
		x"41",	--2094
		x"00",	--2095
		x"00",	--2096
		x"41",	--2097
		x"00",	--2098
		x"00",	--2099
		x"43",	--2100
		x"00",	--2101
		x"43",	--2102
		x"00",	--2103
		x"43",	--2104
		x"00",	--2105
		x"43",	--2106
		x"00",	--2107
		x"43",	--2108
		x"00",	--2109
		x"43",	--2110
		x"00",	--2111
		x"43",	--2112
		x"00",	--2113
		x"43",	--2114
		x"00",	--2115
		x"41",	--2116
		x"43",	--2117
		x"00",	--2118
		x"43",	--2119
		x"00",	--2120
		x"43",	--2121
		x"00",	--2122
		x"43",	--2123
		x"00",	--2124
		x"43",	--2125
		x"00",	--2126
		x"43",	--2127
		x"00",	--2128
		x"41",	--2129
		x"4d",	--2130
		x"00",	--2131
		x"4e",	--2132
		x"00",	--2133
		x"41",	--2134
		x"4d",	--2135
		x"00",	--2136
		x"4e",	--2137
		x"00",	--2138
		x"41",	--2139
		x"4d",	--2140
		x"00",	--2141
		x"4e",	--2142
		x"00",	--2143
		x"41",	--2144
		x"4d",	--2145
		x"00",	--2146
		x"4e",	--2147
		x"00",	--2148
		x"41",	--2149
		x"4d",	--2150
		x"00",	--2151
		x"4e",	--2152
		x"00",	--2153
		x"41",	--2154
		x"12",	--2155
		x"12",	--2156
		x"12",	--2157
		x"12",	--2158
		x"12",	--2159
		x"12",	--2160
		x"12",	--2161
		x"4f",	--2162
		x"4d",	--2163
		x"4e",	--2164
		x"4f",	--2165
		x"00",	--2166
		x"4f",	--2167
		x"00",	--2168
		x"4f",	--2169
		x"00",	--2170
		x"4f",	--2171
		x"00",	--2172
		x"4a",	--2173
		x"4b",	--2174
		x"46",	--2175
		x"47",	--2176
		x"12",	--2177
		x"c2",	--2178
		x"49",	--2179
		x"00",	--2180
		x"49",	--2181
		x"00",	--2182
		x"93",	--2183
		x"34",	--2184
		x"46",	--2185
		x"47",	--2186
		x"12",	--2187
		x"bd",	--2188
		x"4e",	--2189
		x"4f",	--2190
		x"4e",	--2191
		x"00",	--2192
		x"4f",	--2193
		x"00",	--2194
		x"4e",	--2195
		x"4f",	--2196
		x"4a",	--2197
		x"4b",	--2198
		x"12",	--2199
		x"c2",	--2200
		x"93",	--2201
		x"34",	--2202
		x"4a",	--2203
		x"00",	--2204
		x"4b",	--2205
		x"00",	--2206
		x"44",	--2207
		x"45",	--2208
		x"4a",	--2209
		x"4b",	--2210
		x"12",	--2211
		x"be",	--2212
		x"4e",	--2213
		x"4f",	--2214
		x"49",	--2215
		x"00",	--2216
		x"49",	--2217
		x"00",	--2218
		x"12",	--2219
		x"bd",	--2220
		x"4e",	--2221
		x"4f",	--2222
		x"4e",	--2223
		x"00",	--2224
		x"4f",	--2225
		x"00",	--2226
		x"49",	--2227
		x"49",	--2228
		x"00",	--2229
		x"4a",	--2230
		x"4b",	--2231
		x"12",	--2232
		x"be",	--2233
		x"4e",	--2234
		x"4f",	--2235
		x"49",	--2236
		x"00",	--2237
		x"49",	--2238
		x"00",	--2239
		x"46",	--2240
		x"47",	--2241
		x"12",	--2242
		x"be",	--2243
		x"44",	--2244
		x"45",	--2245
		x"12",	--2246
		x"bd",	--2247
		x"4e",	--2248
		x"4f",	--2249
		x"49",	--2250
		x"00",	--2251
		x"49",	--2252
		x"00",	--2253
		x"4a",	--2254
		x"4b",	--2255
		x"12",	--2256
		x"be",	--2257
		x"49",	--2258
		x"00",	--2259
		x"49",	--2260
		x"00",	--2261
		x"12",	--2262
		x"be",	--2263
		x"46",	--2264
		x"47",	--2265
		x"12",	--2266
		x"bd",	--2267
		x"41",	--2268
		x"41",	--2269
		x"41",	--2270
		x"41",	--2271
		x"41",	--2272
		x"41",	--2273
		x"41",	--2274
		x"41",	--2275
		x"46",	--2276
		x"47",	--2277
		x"12",	--2278
		x"be",	--2279
		x"4e",	--2280
		x"4f",	--2281
		x"4e",	--2282
		x"00",	--2283
		x"4f",	--2284
		x"00",	--2285
		x"4e",	--2286
		x"4f",	--2287
		x"4a",	--2288
		x"4b",	--2289
		x"12",	--2290
		x"c2",	--2291
		x"93",	--2292
		x"24",	--2293
		x"37",	--2294
		x"46",	--2295
		x"47",	--2296
		x"3f",	--2297
		x"12",	--2298
		x"12",	--2299
		x"83",	--2300
		x"4f",	--2301
		x"4e",	--2302
		x"12",	--2303
		x"d7",	--2304
		x"12",	--2305
		x"9c",	--2306
		x"53",	--2307
		x"90",	--2308
		x"00",	--2309
		x"38",	--2310
		x"41",	--2311
		x"4b",	--2312
		x"00",	--2313
		x"12",	--2314
		x"87",	--2315
		x"4f",	--2316
		x"41",	--2317
		x"4b",	--2318
		x"00",	--2319
		x"12",	--2320
		x"87",	--2321
		x"4f",	--2322
		x"12",	--2323
		x"12",	--2324
		x"12",	--2325
		x"d7",	--2326
		x"12",	--2327
		x"9c",	--2328
		x"50",	--2329
		x"00",	--2330
		x"4b",	--2331
		x"00",	--2332
		x"43",	--2333
		x"53",	--2334
		x"41",	--2335
		x"41",	--2336
		x"41",	--2337
		x"12",	--2338
		x"d7",	--2339
		x"12",	--2340
		x"9c",	--2341
		x"40",	--2342
		x"d7",	--2343
		x"00",	--2344
		x"12",	--2345
		x"9c",	--2346
		x"4b",	--2347
		x"00",	--2348
		x"12",	--2349
		x"d7",	--2350
		x"12",	--2351
		x"9c",	--2352
		x"52",	--2353
		x"43",	--2354
		x"3f",	--2355
		x"12",	--2356
		x"83",	--2357
		x"4e",	--2358
		x"93",	--2359
		x"24",	--2360
		x"38",	--2361
		x"12",	--2362
		x"d7",	--2363
		x"12",	--2364
		x"9c",	--2365
		x"53",	--2366
		x"41",	--2367
		x"4b",	--2368
		x"00",	--2369
		x"12",	--2370
		x"87",	--2371
		x"12",	--2372
		x"12",	--2373
		x"12",	--2374
		x"d7",	--2375
		x"12",	--2376
		x"9c",	--2377
		x"50",	--2378
		x"00",	--2379
		x"43",	--2380
		x"53",	--2381
		x"41",	--2382
		x"41",	--2383
		x"12",	--2384
		x"d7",	--2385
		x"12",	--2386
		x"9c",	--2387
		x"40",	--2388
		x"d7",	--2389
		x"00",	--2390
		x"12",	--2391
		x"9c",	--2392
		x"4b",	--2393
		x"00",	--2394
		x"12",	--2395
		x"d7",	--2396
		x"12",	--2397
		x"9c",	--2398
		x"52",	--2399
		x"43",	--2400
		x"3f",	--2401
		x"12",	--2402
		x"12",	--2403
		x"12",	--2404
		x"12",	--2405
		x"12",	--2406
		x"12",	--2407
		x"4e",	--2408
		x"4f",	--2409
		x"4c",	--2410
		x"4d",	--2411
		x"12",	--2412
		x"bd",	--2413
		x"4e",	--2414
		x"4f",	--2415
		x"40",	--2416
		x"0f",	--2417
		x"40",	--2418
		x"c0",	--2419
		x"12",	--2420
		x"c3",	--2421
		x"93",	--2422
		x"24",	--2423
		x"38",	--2424
		x"40",	--2425
		x"0f",	--2426
		x"40",	--2427
		x"40",	--2428
		x"4a",	--2429
		x"4b",	--2430
		x"12",	--2431
		x"c2",	--2432
		x"93",	--2433
		x"24",	--2434
		x"34",	--2435
		x"4a",	--2436
		x"4b",	--2437
		x"41",	--2438
		x"41",	--2439
		x"41",	--2440
		x"41",	--2441
		x"41",	--2442
		x"41",	--2443
		x"41",	--2444
		x"40",	--2445
		x"0f",	--2446
		x"40",	--2447
		x"40",	--2448
		x"4a",	--2449
		x"4b",	--2450
		x"12",	--2451
		x"be",	--2452
		x"4e",	--2453
		x"4f",	--2454
		x"3f",	--2455
		x"40",	--2456
		x"0f",	--2457
		x"40",	--2458
		x"40",	--2459
		x"46",	--2460
		x"47",	--2461
		x"12",	--2462
		x"bd",	--2463
		x"48",	--2464
		x"49",	--2465
		x"12",	--2466
		x"bd",	--2467
		x"4e",	--2468
		x"4f",	--2469
		x"3f",	--2470
		x"12",	--2471
		x"4f",	--2472
		x"43",	--2473
		x"00",	--2474
		x"43",	--2475
		x"00",	--2476
		x"43",	--2477
		x"00",	--2478
		x"43",	--2479
		x"00",	--2480
		x"43",	--2481
		x"00",	--2482
		x"43",	--2483
		x"00",	--2484
		x"4d",	--2485
		x"00",	--2486
		x"4e",	--2487
		x"00",	--2488
		x"41",	--2489
		x"00",	--2490
		x"00",	--2491
		x"41",	--2492
		x"00",	--2493
		x"00",	--2494
		x"41",	--2495
		x"00",	--2496
		x"00",	--2497
		x"43",	--2498
		x"00",	--2499
		x"43",	--2500
		x"00",	--2501
		x"43",	--2502
		x"00",	--2503
		x"43",	--2504
		x"00",	--2505
		x"4f",	--2506
		x"40",	--2507
		x"96",	--2508
		x"12",	--2509
		x"99",	--2510
		x"4f",	--2511
		x"00",	--2512
		x"41",	--2513
		x"41",	--2514
		x"4e",	--2515
		x"00",	--2516
		x"4d",	--2517
		x"00",	--2518
		x"41",	--2519
		x"12",	--2520
		x"12",	--2521
		x"12",	--2522
		x"12",	--2523
		x"12",	--2524
		x"12",	--2525
		x"12",	--2526
		x"50",	--2527
		x"ff",	--2528
		x"4f",	--2529
		x"4d",	--2530
		x"00",	--2531
		x"4e",	--2532
		x"00",	--2533
		x"40",	--2534
		x"0f",	--2535
		x"40",	--2536
		x"40",	--2537
		x"4f",	--2538
		x"4f",	--2539
		x"00",	--2540
		x"12",	--2541
		x"be",	--2542
		x"4e",	--2543
		x"4f",	--2544
		x"47",	--2545
		x"00",	--2546
		x"4e",	--2547
		x"10",	--2548
		x"11",	--2549
		x"10",	--2550
		x"11",	--2551
		x"12",	--2552
		x"c3",	--2553
		x"4e",	--2554
		x"4f",	--2555
		x"4a",	--2556
		x"4b",	--2557
		x"12",	--2558
		x"c0",	--2559
		x"4e",	--2560
		x"4f",	--2561
		x"41",	--2562
		x"00",	--2563
		x"41",	--2564
		x"00",	--2565
		x"87",	--2566
		x"00",	--2567
		x"77",	--2568
		x"00",	--2569
		x"41",	--2570
		x"00",	--2571
		x"41",	--2572
		x"00",	--2573
		x"87",	--2574
		x"00",	--2575
		x"77",	--2576
		x"00",	--2577
		x"48",	--2578
		x"49",	--2579
		x"12",	--2580
		x"c3",	--2581
		x"4a",	--2582
		x"4b",	--2583
		x"12",	--2584
		x"be",	--2585
		x"4e",	--2586
		x"00",	--2587
		x"4f",	--2588
		x"00",	--2589
		x"44",	--2590
		x"45",	--2591
		x"12",	--2592
		x"c3",	--2593
		x"4a",	--2594
		x"4b",	--2595
		x"12",	--2596
		x"be",	--2597
		x"4e",	--2598
		x"4f",	--2599
		x"4e",	--2600
		x"4f",	--2601
		x"41",	--2602
		x"41",	--2603
		x"00",	--2604
		x"12",	--2605
		x"bd",	--2606
		x"4e",	--2607
		x"00",	--2608
		x"4f",	--2609
		x"00",	--2610
		x"93",	--2611
		x"20",	--2612
		x"93",	--2613
		x"20",	--2614
		x"93",	--2615
		x"20",	--2616
		x"40",	--2617
		x"96",	--2618
		x"47",	--2619
		x"00",	--2620
		x"47",	--2621
		x"00",	--2622
		x"41",	--2623
		x"41",	--2624
		x"00",	--2625
		x"4a",	--2626
		x"4b",	--2627
		x"12",	--2628
		x"be",	--2629
		x"4e",	--2630
		x"4f",	--2631
		x"48",	--2632
		x"49",	--2633
		x"41",	--2634
		x"00",	--2635
		x"41",	--2636
		x"00",	--2637
		x"12",	--2638
		x"be",	--2639
		x"4a",	--2640
		x"4b",	--2641
		x"12",	--2642
		x"c0",	--2643
		x"4e",	--2644
		x"4f",	--2645
		x"48",	--2646
		x"49",	--2647
		x"48",	--2648
		x"49",	--2649
		x"12",	--2650
		x"bd",	--2651
		x"4e",	--2652
		x"4f",	--2653
		x"4a",	--2654
		x"4b",	--2655
		x"12",	--2656
		x"c0",	--2657
		x"12",	--2658
		x"a1",	--2659
		x"4e",	--2660
		x"00",	--2661
		x"4f",	--2662
		x"00",	--2663
		x"47",	--2664
		x"00",	--2665
		x"47",	--2666
		x"00",	--2667
		x"4a",	--2668
		x"4b",	--2669
		x"12",	--2670
		x"a1",	--2671
		x"44",	--2672
		x"45",	--2673
		x"12",	--2674
		x"be",	--2675
		x"4e",	--2676
		x"4f",	--2677
		x"47",	--2678
		x"00",	--2679
		x"47",	--2680
		x"00",	--2681
		x"12",	--2682
		x"be",	--2683
		x"4e",	--2684
		x"00",	--2685
		x"4f",	--2686
		x"00",	--2687
		x"4a",	--2688
		x"4b",	--2689
		x"12",	--2690
		x"b6",	--2691
		x"44",	--2692
		x"45",	--2693
		x"12",	--2694
		x"be",	--2695
		x"47",	--2696
		x"00",	--2697
		x"47",	--2698
		x"00",	--2699
		x"12",	--2700
		x"bd",	--2701
		x"4e",	--2702
		x"4f",	--2703
		x"41",	--2704
		x"41",	--2705
		x"00",	--2706
		x"4a",	--2707
		x"4b",	--2708
		x"12",	--2709
		x"92",	--2710
		x"4e",	--2711
		x"4f",	--2712
		x"4e",	--2713
		x"00",	--2714
		x"4f",	--2715
		x"00",	--2716
		x"12",	--2717
		x"a1",	--2718
		x"44",	--2719
		x"45",	--2720
		x"12",	--2721
		x"be",	--2722
		x"41",	--2723
		x"00",	--2724
		x"41",	--2725
		x"00",	--2726
		x"12",	--2727
		x"bd",	--2728
		x"4e",	--2729
		x"00",	--2730
		x"4f",	--2731
		x"00",	--2732
		x"4a",	--2733
		x"4b",	--2734
		x"12",	--2735
		x"b6",	--2736
		x"44",	--2737
		x"45",	--2738
		x"12",	--2739
		x"be",	--2740
		x"4e",	--2741
		x"4f",	--2742
		x"48",	--2743
		x"49",	--2744
		x"12",	--2745
		x"be",	--2746
		x"4e",	--2747
		x"00",	--2748
		x"4f",	--2749
		x"00",	--2750
		x"41",	--2751
		x"00",	--2752
		x"00",	--2753
		x"41",	--2754
		x"00",	--2755
		x"00",	--2756
		x"41",	--2757
		x"00",	--2758
		x"00",	--2759
		x"41",	--2760
		x"00",	--2761
		x"00",	--2762
		x"50",	--2763
		x"00",	--2764
		x"41",	--2765
		x"41",	--2766
		x"41",	--2767
		x"41",	--2768
		x"41",	--2769
		x"41",	--2770
		x"41",	--2771
		x"41",	--2772
		x"94",	--2773
		x"23",	--2774
		x"95",	--2775
		x"23",	--2776
		x"43",	--2777
		x"40",	--2778
		x"3f",	--2779
		x"41",	--2780
		x"00",	--2781
		x"41",	--2782
		x"00",	--2783
		x"12",	--2784
		x"be",	--2785
		x"4e",	--2786
		x"4f",	--2787
		x"47",	--2788
		x"00",	--2789
		x"47",	--2790
		x"00",	--2791
		x"48",	--2792
		x"49",	--2793
		x"12",	--2794
		x"b6",	--2795
		x"4a",	--2796
		x"4b",	--2797
		x"12",	--2798
		x"be",	--2799
		x"4e",	--2800
		x"4f",	--2801
		x"47",	--2802
		x"00",	--2803
		x"47",	--2804
		x"00",	--2805
		x"12",	--2806
		x"bd",	--2807
		x"4e",	--2808
		x"00",	--2809
		x"4f",	--2810
		x"00",	--2811
		x"48",	--2812
		x"49",	--2813
		x"12",	--2814
		x"a1",	--2815
		x"4a",	--2816
		x"4b",	--2817
		x"12",	--2818
		x"be",	--2819
		x"4e",	--2820
		x"4f",	--2821
		x"47",	--2822
		x"00",	--2823
		x"47",	--2824
		x"00",	--2825
		x"12",	--2826
		x"bd",	--2827
		x"4e",	--2828
		x"00",	--2829
		x"4f",	--2830
		x"00",	--2831
		x"3f",	--2832
		x"93",	--2833
		x"27",	--2834
		x"40",	--2835
		x"94",	--2836
		x"12",	--2837
		x"12",	--2838
		x"12",	--2839
		x"4f",	--2840
		x"4f",	--2841
		x"00",	--2842
		x"12",	--2843
		x"9a",	--2844
		x"4e",	--2845
		x"4f",	--2846
		x"49",	--2847
		x"00",	--2848
		x"12",	--2849
		x"9a",	--2850
		x"4a",	--2851
		x"4b",	--2852
		x"e3",	--2853
		x"e3",	--2854
		x"53",	--2855
		x"63",	--2856
		x"12",	--2857
		x"12",	--2858
		x"4e",	--2859
		x"4f",	--2860
		x"49",	--2861
		x"12",	--2862
		x"93",	--2863
		x"52",	--2864
		x"41",	--2865
		x"41",	--2866
		x"41",	--2867
		x"41",	--2868
		x"43",	--2869
		x"4f",	--2870
		x"00",	--2871
		x"12",	--2872
		x"99",	--2873
		x"41",	--2874
		x"4f",	--2875
		x"00",	--2876
		x"12",	--2877
		x"99",	--2878
		x"41",	--2879
		x"12",	--2880
		x"12",	--2881
		x"4e",	--2882
		x"4c",	--2883
		x"4e",	--2884
		x"00",	--2885
		x"4d",	--2886
		x"00",	--2887
		x"4c",	--2888
		x"00",	--2889
		x"4d",	--2890
		x"43",	--2891
		x"40",	--2892
		x"36",	--2893
		x"40",	--2894
		x"01",	--2895
		x"12",	--2896
		x"d2",	--2897
		x"4e",	--2898
		x"00",	--2899
		x"12",	--2900
		x"c2",	--2901
		x"43",	--2902
		x"4a",	--2903
		x"01",	--2904
		x"40",	--2905
		x"00",	--2906
		x"01",	--2907
		x"42",	--2908
		x"01",	--2909
		x"00",	--2910
		x"41",	--2911
		x"43",	--2912
		x"41",	--2913
		x"41",	--2914
		x"41",	--2915
		x"12",	--2916
		x"12",	--2917
		x"12",	--2918
		x"43",	--2919
		x"00",	--2920
		x"40",	--2921
		x"3f",	--2922
		x"00",	--2923
		x"4f",	--2924
		x"4b",	--2925
		x"00",	--2926
		x"43",	--2927
		x"12",	--2928
		x"c4",	--2929
		x"43",	--2930
		x"40",	--2931
		x"3f",	--2932
		x"12",	--2933
		x"be",	--2934
		x"4e",	--2935
		x"4f",	--2936
		x"4b",	--2937
		x"00",	--2938
		x"43",	--2939
		x"12",	--2940
		x"c4",	--2941
		x"4e",	--2942
		x"4f",	--2943
		x"48",	--2944
		x"49",	--2945
		x"12",	--2946
		x"be",	--2947
		x"12",	--2948
		x"ba",	--2949
		x"4e",	--2950
		x"00",	--2951
		x"43",	--2952
		x"00",	--2953
		x"41",	--2954
		x"41",	--2955
		x"41",	--2956
		x"41",	--2957
		x"12",	--2958
		x"12",	--2959
		x"12",	--2960
		x"4d",	--2961
		x"4e",	--2962
		x"4d",	--2963
		x"00",	--2964
		x"4e",	--2965
		x"00",	--2966
		x"4f",	--2967
		x"49",	--2968
		x"00",	--2969
		x"43",	--2970
		x"12",	--2971
		x"c4",	--2972
		x"4e",	--2973
		x"4f",	--2974
		x"4a",	--2975
		x"4b",	--2976
		x"12",	--2977
		x"be",	--2978
		x"4e",	--2979
		x"4f",	--2980
		x"49",	--2981
		x"00",	--2982
		x"43",	--2983
		x"12",	--2984
		x"c4",	--2985
		x"4e",	--2986
		x"4f",	--2987
		x"4a",	--2988
		x"4b",	--2989
		x"12",	--2990
		x"be",	--2991
		x"12",	--2992
		x"ba",	--2993
		x"4e",	--2994
		x"00",	--2995
		x"41",	--2996
		x"41",	--2997
		x"41",	--2998
		x"41",	--2999
		x"4f",	--3000
		x"4e",	--3001
		x"00",	--3002
		x"41",	--3003
		x"12",	--3004
		x"12",	--3005
		x"93",	--3006
		x"02",	--3007
		x"38",	--3008
		x"40",	--3009
		x"02",	--3010
		x"43",	--3011
		x"12",	--3012
		x"4b",	--3013
		x"ff",	--3014
		x"11",	--3015
		x"12",	--3016
		x"12",	--3017
		x"d7",	--3018
		x"12",	--3019
		x"9c",	--3020
		x"50",	--3021
		x"00",	--3022
		x"53",	--3023
		x"50",	--3024
		x"00",	--3025
		x"92",	--3026
		x"02",	--3027
		x"3b",	--3028
		x"43",	--3029
		x"41",	--3030
		x"41",	--3031
		x"41",	--3032
		x"42",	--3033
		x"02",	--3034
		x"90",	--3035
		x"00",	--3036
		x"34",	--3037
		x"4e",	--3038
		x"5f",	--3039
		x"5e",	--3040
		x"5f",	--3041
		x"50",	--3042
		x"02",	--3043
		x"40",	--3044
		x"00",	--3045
		x"00",	--3046
		x"40",	--3047
		x"97",	--3048
		x"00",	--3049
		x"40",	--3050
		x"02",	--3051
		x"00",	--3052
		x"53",	--3053
		x"4e",	--3054
		x"02",	--3055
		x"41",	--3056
		x"12",	--3057
		x"42",	--3058
		x"02",	--3059
		x"90",	--3060
		x"00",	--3061
		x"34",	--3062
		x"4b",	--3063
		x"5c",	--3064
		x"5b",	--3065
		x"5c",	--3066
		x"50",	--3067
		x"02",	--3068
		x"4f",	--3069
		x"00",	--3070
		x"4e",	--3071
		x"00",	--3072
		x"4d",	--3073
		x"00",	--3074
		x"53",	--3075
		x"4b",	--3076
		x"02",	--3077
		x"43",	--3078
		x"41",	--3079
		x"41",	--3080
		x"43",	--3081
		x"3f",	--3082
		x"12",	--3083
		x"50",	--3084
		x"ff",	--3085
		x"42",	--3086
		x"02",	--3087
		x"93",	--3088
		x"38",	--3089
		x"92",	--3090
		x"02",	--3091
		x"24",	--3092
		x"40",	--3093
		x"02",	--3094
		x"43",	--3095
		x"3c",	--3096
		x"50",	--3097
		x"00",	--3098
		x"9f",	--3099
		x"ff",	--3100
		x"24",	--3101
		x"53",	--3102
		x"9b",	--3103
		x"23",	--3104
		x"12",	--3105
		x"d7",	--3106
		x"12",	--3107
		x"9c",	--3108
		x"53",	--3109
		x"43",	--3110
		x"50",	--3111
		x"00",	--3112
		x"41",	--3113
		x"41",	--3114
		x"43",	--3115
		x"4e",	--3116
		x"00",	--3117
		x"4e",	--3118
		x"93",	--3119
		x"24",	--3120
		x"53",	--3121
		x"43",	--3122
		x"3c",	--3123
		x"4e",	--3124
		x"93",	--3125
		x"24",	--3126
		x"53",	--3127
		x"92",	--3128
		x"34",	--3129
		x"90",	--3130
		x"00",	--3131
		x"23",	--3132
		x"43",	--3133
		x"ff",	--3134
		x"4f",	--3135
		x"5d",	--3136
		x"51",	--3137
		x"4e",	--3138
		x"00",	--3139
		x"53",	--3140
		x"4e",	--3141
		x"93",	--3142
		x"23",	--3143
		x"4c",	--3144
		x"5e",	--3145
		x"5e",	--3146
		x"5c",	--3147
		x"50",	--3148
		x"02",	--3149
		x"41",	--3150
		x"12",	--3151
		x"00",	--3152
		x"50",	--3153
		x"00",	--3154
		x"41",	--3155
		x"41",	--3156
		x"43",	--3157
		x"3f",	--3158
		x"4e",	--3159
		x"00",	--3160
		x"43",	--3161
		x"41",	--3162
		x"5e",	--3163
		x"5f",	--3164
		x"4e",	--3165
		x"41",	--3166
		x"12",	--3167
		x"12",	--3168
		x"5e",	--3169
		x"5f",	--3170
		x"4e",	--3171
		x"43",	--3172
		x"4c",	--3173
		x"4d",	--3174
		x"5e",	--3175
		x"6f",	--3176
		x"4e",	--3177
		x"4f",	--3178
		x"5a",	--3179
		x"6b",	--3180
		x"5a",	--3181
		x"6b",	--3182
		x"40",	--3183
		x"00",	--3184
		x"43",	--3185
		x"5a",	--3186
		x"6b",	--3187
		x"12",	--3188
		x"d2",	--3189
		x"4e",	--3190
		x"41",	--3191
		x"41",	--3192
		x"41",	--3193
		x"d0",	--3194
		x"02",	--3195
		x"01",	--3196
		x"40",	--3197
		x"0b",	--3198
		x"01",	--3199
		x"43",	--3200
		x"41",	--3201
		x"12",	--3202
		x"4f",	--3203
		x"42",	--3204
		x"02",	--3205
		x"90",	--3206
		x"00",	--3207
		x"34",	--3208
		x"4f",	--3209
		x"5c",	--3210
		x"4c",	--3211
		x"5d",	--3212
		x"5d",	--3213
		x"5d",	--3214
		x"8c",	--3215
		x"50",	--3216
		x"03",	--3217
		x"43",	--3218
		x"00",	--3219
		x"43",	--3220
		x"00",	--3221
		x"43",	--3222
		x"00",	--3223
		x"4b",	--3224
		x"00",	--3225
		x"4e",	--3226
		x"00",	--3227
		x"4f",	--3228
		x"53",	--3229
		x"4e",	--3230
		x"02",	--3231
		x"41",	--3232
		x"41",	--3233
		x"43",	--3234
		x"3f",	--3235
		x"5f",	--3236
		x"4f",	--3237
		x"5c",	--3238
		x"5c",	--3239
		x"5c",	--3240
		x"8f",	--3241
		x"50",	--3242
		x"03",	--3243
		x"43",	--3244
		x"00",	--3245
		x"4e",	--3246
		x"00",	--3247
		x"43",	--3248
		x"00",	--3249
		x"4d",	--3250
		x"00",	--3251
		x"43",	--3252
		x"00",	--3253
		x"43",	--3254
		x"41",	--3255
		x"5f",	--3256
		x"4f",	--3257
		x"5e",	--3258
		x"5e",	--3259
		x"5e",	--3260
		x"8f",	--3261
		x"43",	--3262
		x"03",	--3263
		x"43",	--3264
		x"41",	--3265
		x"12",	--3266
		x"12",	--3267
		x"12",	--3268
		x"12",	--3269
		x"12",	--3270
		x"12",	--3271
		x"12",	--3272
		x"12",	--3273
		x"12",	--3274
		x"93",	--3275
		x"02",	--3276
		x"38",	--3277
		x"40",	--3278
		x"03",	--3279
		x"4a",	--3280
		x"53",	--3281
		x"4a",	--3282
		x"52",	--3283
		x"4a",	--3284
		x"50",	--3285
		x"00",	--3286
		x"43",	--3287
		x"3c",	--3288
		x"53",	--3289
		x"4f",	--3290
		x"00",	--3291
		x"53",	--3292
		x"50",	--3293
		x"00",	--3294
		x"50",	--3295
		x"00",	--3296
		x"50",	--3297
		x"00",	--3298
		x"50",	--3299
		x"00",	--3300
		x"92",	--3301
		x"02",	--3302
		x"34",	--3303
		x"93",	--3304
		x"00",	--3305
		x"27",	--3306
		x"4b",	--3307
		x"9b",	--3308
		x"00",	--3309
		x"2b",	--3310
		x"43",	--3311
		x"00",	--3312
		x"4b",	--3313
		x"00",	--3314
		x"12",	--3315
		x"00",	--3316
		x"93",	--3317
		x"00",	--3318
		x"27",	--3319
		x"47",	--3320
		x"53",	--3321
		x"4f",	--3322
		x"00",	--3323
		x"98",	--3324
		x"2b",	--3325
		x"43",	--3326
		x"00",	--3327
		x"3f",	--3328
		x"f0",	--3329
		x"ff",	--3330
		x"01",	--3331
		x"41",	--3332
		x"41",	--3333
		x"41",	--3334
		x"41",	--3335
		x"41",	--3336
		x"41",	--3337
		x"41",	--3338
		x"41",	--3339
		x"41",	--3340
		x"13",	--3341
		x"4e",	--3342
		x"00",	--3343
		x"43",	--3344
		x"41",	--3345
		x"4f",	--3346
		x"4f",	--3347
		x"4f",	--3348
		x"00",	--3349
		x"41",	--3350
		x"43",	--3351
		x"00",	--3352
		x"41",	--3353
		x"4e",	--3354
		x"00",	--3355
		x"40",	--3356
		x"9a",	--3357
		x"12",	--3358
		x"99",	--3359
		x"4f",	--3360
		x"02",	--3361
		x"43",	--3362
		x"41",	--3363
		x"4d",	--3364
		x"4f",	--3365
		x"4e",	--3366
		x"00",	--3367
		x"43",	--3368
		x"4c",	--3369
		x"42",	--3370
		x"02",	--3371
		x"12",	--3372
		x"99",	--3373
		x"41",	--3374
		x"42",	--3375
		x"00",	--3376
		x"f2",	--3377
		x"23",	--3378
		x"4f",	--3379
		x"00",	--3380
		x"43",	--3381
		x"41",	--3382
		x"f0",	--3383
		x"00",	--3384
		x"4f",	--3385
		x"d8",	--3386
		x"11",	--3387
		x"12",	--3388
		x"9a",	--3389
		x"41",	--3390
		x"12",	--3391
		x"4f",	--3392
		x"4f",	--3393
		x"11",	--3394
		x"11",	--3395
		x"11",	--3396
		x"11",	--3397
		x"4e",	--3398
		x"12",	--3399
		x"9a",	--3400
		x"4b",	--3401
		x"12",	--3402
		x"9a",	--3403
		x"41",	--3404
		x"41",	--3405
		x"12",	--3406
		x"12",	--3407
		x"4f",	--3408
		x"40",	--3409
		x"00",	--3410
		x"4a",	--3411
		x"4b",	--3412
		x"f0",	--3413
		x"00",	--3414
		x"24",	--3415
		x"11",	--3416
		x"53",	--3417
		x"23",	--3418
		x"f3",	--3419
		x"24",	--3420
		x"40",	--3421
		x"00",	--3422
		x"12",	--3423
		x"9a",	--3424
		x"53",	--3425
		x"93",	--3426
		x"23",	--3427
		x"41",	--3428
		x"41",	--3429
		x"41",	--3430
		x"40",	--3431
		x"00",	--3432
		x"3f",	--3433
		x"12",	--3434
		x"4f",	--3435
		x"4f",	--3436
		x"10",	--3437
		x"11",	--3438
		x"4e",	--3439
		x"12",	--3440
		x"9a",	--3441
		x"4b",	--3442
		x"12",	--3443
		x"9a",	--3444
		x"41",	--3445
		x"41",	--3446
		x"12",	--3447
		x"12",	--3448
		x"4e",	--3449
		x"4f",	--3450
		x"4f",	--3451
		x"10",	--3452
		x"11",	--3453
		x"4d",	--3454
		x"12",	--3455
		x"9a",	--3456
		x"4b",	--3457
		x"12",	--3458
		x"9a",	--3459
		x"4b",	--3460
		x"4a",	--3461
		x"10",	--3462
		x"10",	--3463
		x"ec",	--3464
		x"ec",	--3465
		x"4d",	--3466
		x"12",	--3467
		x"9a",	--3468
		x"4a",	--3469
		x"12",	--3470
		x"9a",	--3471
		x"41",	--3472
		x"41",	--3473
		x"41",	--3474
		x"12",	--3475
		x"12",	--3476
		x"12",	--3477
		x"4f",	--3478
		x"93",	--3479
		x"24",	--3480
		x"4e",	--3481
		x"53",	--3482
		x"43",	--3483
		x"4a",	--3484
		x"5b",	--3485
		x"4d",	--3486
		x"11",	--3487
		x"12",	--3488
		x"9a",	--3489
		x"99",	--3490
		x"24",	--3491
		x"53",	--3492
		x"b0",	--3493
		x"00",	--3494
		x"20",	--3495
		x"40",	--3496
		x"00",	--3497
		x"12",	--3498
		x"9a",	--3499
		x"3f",	--3500
		x"40",	--3501
		x"00",	--3502
		x"12",	--3503
		x"9a",	--3504
		x"3f",	--3505
		x"41",	--3506
		x"41",	--3507
		x"41",	--3508
		x"41",	--3509
		x"12",	--3510
		x"12",	--3511
		x"12",	--3512
		x"4f",	--3513
		x"93",	--3514
		x"24",	--3515
		x"4e",	--3516
		x"53",	--3517
		x"43",	--3518
		x"4a",	--3519
		x"11",	--3520
		x"12",	--3521
		x"9a",	--3522
		x"99",	--3523
		x"24",	--3524
		x"53",	--3525
		x"b0",	--3526
		x"00",	--3527
		x"23",	--3528
		x"40",	--3529
		x"00",	--3530
		x"12",	--3531
		x"9a",	--3532
		x"4a",	--3533
		x"11",	--3534
		x"12",	--3535
		x"9a",	--3536
		x"99",	--3537
		x"23",	--3538
		x"41",	--3539
		x"41",	--3540
		x"41",	--3541
		x"41",	--3542
		x"12",	--3543
		x"12",	--3544
		x"12",	--3545
		x"50",	--3546
		x"ff",	--3547
		x"4f",	--3548
		x"93",	--3549
		x"38",	--3550
		x"90",	--3551
		x"00",	--3552
		x"38",	--3553
		x"43",	--3554
		x"41",	--3555
		x"59",	--3556
		x"40",	--3557
		x"00",	--3558
		x"4b",	--3559
		x"12",	--3560
		x"d2",	--3561
		x"50",	--3562
		x"00",	--3563
		x"4f",	--3564
		x"00",	--3565
		x"53",	--3566
		x"40",	--3567
		x"00",	--3568
		x"4b",	--3569
		x"12",	--3570
		x"d2",	--3571
		x"4f",	--3572
		x"90",	--3573
		x"00",	--3574
		x"37",	--3575
		x"49",	--3576
		x"53",	--3577
		x"51",	--3578
		x"40",	--3579
		x"00",	--3580
		x"4b",	--3581
		x"12",	--3582
		x"d2",	--3583
		x"50",	--3584
		x"00",	--3585
		x"4f",	--3586
		x"00",	--3587
		x"53",	--3588
		x"41",	--3589
		x"5a",	--3590
		x"4f",	--3591
		x"11",	--3592
		x"12",	--3593
		x"9a",	--3594
		x"93",	--3595
		x"23",	--3596
		x"50",	--3597
		x"00",	--3598
		x"41",	--3599
		x"41",	--3600
		x"41",	--3601
		x"41",	--3602
		x"40",	--3603
		x"00",	--3604
		x"12",	--3605
		x"9a",	--3606
		x"e3",	--3607
		x"53",	--3608
		x"3f",	--3609
		x"43",	--3610
		x"43",	--3611
		x"3f",	--3612
		x"12",	--3613
		x"12",	--3614
		x"12",	--3615
		x"41",	--3616
		x"52",	--3617
		x"4b",	--3618
		x"49",	--3619
		x"93",	--3620
		x"20",	--3621
		x"3c",	--3622
		x"11",	--3623
		x"12",	--3624
		x"9a",	--3625
		x"49",	--3626
		x"4a",	--3627
		x"53",	--3628
		x"4a",	--3629
		x"00",	--3630
		x"93",	--3631
		x"24",	--3632
		x"90",	--3633
		x"00",	--3634
		x"23",	--3635
		x"49",	--3636
		x"53",	--3637
		x"49",	--3638
		x"00",	--3639
		x"50",	--3640
		x"ff",	--3641
		x"90",	--3642
		x"00",	--3643
		x"2f",	--3644
		x"4f",	--3645
		x"5f",	--3646
		x"4f",	--3647
		x"d7",	--3648
		x"41",	--3649
		x"41",	--3650
		x"41",	--3651
		x"41",	--3652
		x"4b",	--3653
		x"52",	--3654
		x"4b",	--3655
		x"00",	--3656
		x"4b",	--3657
		x"12",	--3658
		x"9b",	--3659
		x"49",	--3660
		x"3f",	--3661
		x"4b",	--3662
		x"53",	--3663
		x"4b",	--3664
		x"12",	--3665
		x"9a",	--3666
		x"49",	--3667
		x"3f",	--3668
		x"4b",	--3669
		x"53",	--3670
		x"4f",	--3671
		x"49",	--3672
		x"93",	--3673
		x"27",	--3674
		x"53",	--3675
		x"11",	--3676
		x"12",	--3677
		x"9a",	--3678
		x"49",	--3679
		x"93",	--3680
		x"23",	--3681
		x"3f",	--3682
		x"4b",	--3683
		x"52",	--3684
		x"4b",	--3685
		x"00",	--3686
		x"4b",	--3687
		x"12",	--3688
		x"9b",	--3689
		x"49",	--3690
		x"3f",	--3691
		x"4b",	--3692
		x"53",	--3693
		x"4b",	--3694
		x"4e",	--3695
		x"10",	--3696
		x"11",	--3697
		x"10",	--3698
		x"11",	--3699
		x"12",	--3700
		x"9a",	--3701
		x"49",	--3702
		x"3f",	--3703
		x"4b",	--3704
		x"53",	--3705
		x"4b",	--3706
		x"12",	--3707
		x"9b",	--3708
		x"49",	--3709
		x"3f",	--3710
		x"4b",	--3711
		x"53",	--3712
		x"4b",	--3713
		x"12",	--3714
		x"9a",	--3715
		x"49",	--3716
		x"3f",	--3717
		x"4b",	--3718
		x"53",	--3719
		x"4b",	--3720
		x"12",	--3721
		x"9a",	--3722
		x"49",	--3723
		x"3f",	--3724
		x"4b",	--3725
		x"53",	--3726
		x"4b",	--3727
		x"12",	--3728
		x"9a",	--3729
		x"49",	--3730
		x"3f",	--3731
		x"40",	--3732
		x"00",	--3733
		x"12",	--3734
		x"9a",	--3735
		x"3f",	--3736
		x"12",	--3737
		x"12",	--3738
		x"42",	--3739
		x"02",	--3740
		x"42",	--3741
		x"00",	--3742
		x"05",	--3743
		x"42",	--3744
		x"02",	--3745
		x"90",	--3746
		x"00",	--3747
		x"34",	--3748
		x"53",	--3749
		x"02",	--3750
		x"42",	--3751
		x"02",	--3752
		x"42",	--3753
		x"02",	--3754
		x"9f",	--3755
		x"20",	--3756
		x"53",	--3757
		x"02",	--3758
		x"40",	--3759
		x"00",	--3760
		x"00",	--3761
		x"41",	--3762
		x"41",	--3763
		x"c0",	--3764
		x"00",	--3765
		x"00",	--3766
		x"13",	--3767
		x"43",	--3768
		x"02",	--3769
		x"3f",	--3770
		x"4e",	--3771
		x"4f",	--3772
		x"40",	--3773
		x"36",	--3774
		x"40",	--3775
		x"01",	--3776
		x"12",	--3777
		x"d2",	--3778
		x"53",	--3779
		x"4e",	--3780
		x"00",	--3781
		x"40",	--3782
		x"00",	--3783
		x"00",	--3784
		x"41",	--3785
		x"42",	--3786
		x"02",	--3787
		x"42",	--3788
		x"02",	--3789
		x"9f",	--3790
		x"38",	--3791
		x"42",	--3792
		x"02",	--3793
		x"82",	--3794
		x"02",	--3795
		x"41",	--3796
		x"42",	--3797
		x"02",	--3798
		x"42",	--3799
		x"02",	--3800
		x"40",	--3801
		x"00",	--3802
		x"8d",	--3803
		x"8e",	--3804
		x"41",	--3805
		x"42",	--3806
		x"02",	--3807
		x"4f",	--3808
		x"05",	--3809
		x"42",	--3810
		x"02",	--3811
		x"42",	--3812
		x"02",	--3813
		x"9e",	--3814
		x"24",	--3815
		x"42",	--3816
		x"02",	--3817
		x"90",	--3818
		x"00",	--3819
		x"38",	--3820
		x"43",	--3821
		x"02",	--3822
		x"41",	--3823
		x"53",	--3824
		x"02",	--3825
		x"41",	--3826
		x"43",	--3827
		x"41",	--3828
		x"12",	--3829
		x"12",	--3830
		x"12",	--3831
		x"12",	--3832
		x"12",	--3833
		x"12",	--3834
		x"12",	--3835
		x"12",	--3836
		x"82",	--3837
		x"4e",	--3838
		x"4f",	--3839
		x"4e",	--3840
		x"00",	--3841
		x"4f",	--3842
		x"00",	--3843
		x"4e",	--3844
		x"4f",	--3845
		x"f3",	--3846
		x"f0",	--3847
		x"7f",	--3848
		x"90",	--3849
		x"50",	--3850
		x"38",	--3851
		x"90",	--3852
		x"7f",	--3853
		x"38",	--3854
		x"20",	--3855
		x"93",	--3856
		x"28",	--3857
		x"44",	--3858
		x"45",	--3859
		x"44",	--3860
		x"45",	--3861
		x"12",	--3862
		x"bd",	--3863
		x"40",	--3864
		x"a0",	--3865
		x"93",	--3866
		x"00",	--3867
		x"34",	--3868
		x"40",	--3869
		x"a1",	--3870
		x"20",	--3871
		x"93",	--3872
		x"00",	--3873
		x"2c",	--3874
		x"40",	--3875
		x"a1",	--3876
		x"40",	--3877
		x"0f",	--3878
		x"40",	--3879
		x"3f",	--3880
		x"40",	--3881
		x"a1",	--3882
		x"90",	--3883
		x"3e",	--3884
		x"38",	--3885
		x"4e",	--3886
		x"4f",	--3887
		x"f0",	--3888
		x"7f",	--3889
		x"90",	--3890
		x"3f",	--3891
		x"38",	--3892
		x"3c",	--3893
		x"90",	--3894
		x"31",	--3895
		x"34",	--3896
		x"40",	--3897
		x"f2",	--3898
		x"40",	--3899
		x"71",	--3900
		x"12",	--3901
		x"bd",	--3902
		x"43",	--3903
		x"40",	--3904
		x"3f",	--3905
		x"12",	--3906
		x"c2",	--3907
		x"93",	--3908
		x"24",	--3909
		x"38",	--3910
		x"40",	--3911
		x"a1",	--3912
		x"43",	--3913
		x"43",	--3914
		x"3c",	--3915
		x"90",	--3916
		x"40",	--3917
		x"38",	--3918
		x"3c",	--3919
		x"90",	--3920
		x"3f",	--3921
		x"38",	--3922
		x"43",	--3923
		x"40",	--3924
		x"3f",	--3925
		x"4a",	--3926
		x"4b",	--3927
		x"12",	--3928
		x"be",	--3929
		x"4e",	--3930
		x"4f",	--3931
		x"43",	--3932
		x"40",	--3933
		x"3f",	--3934
		x"4a",	--3935
		x"4b",	--3936
		x"12",	--3937
		x"bd",	--3938
		x"4e",	--3939
		x"4f",	--3940
		x"48",	--3941
		x"49",	--3942
		x"12",	--3943
		x"c0",	--3944
		x"4e",	--3945
		x"4f",	--3946
		x"43",	--3947
		x"43",	--3948
		x"3c",	--3949
		x"4a",	--3950
		x"4b",	--3951
		x"4a",	--3952
		x"4b",	--3953
		x"12",	--3954
		x"bd",	--3955
		x"43",	--3956
		x"40",	--3957
		x"3f",	--3958
		x"12",	--3959
		x"be",	--3960
		x"4e",	--3961
		x"4f",	--3962
		x"43",	--3963
		x"40",	--3964
		x"40",	--3965
		x"4a",	--3966
		x"4b",	--3967
		x"12",	--3968
		x"bd",	--3969
		x"4e",	--3970
		x"4f",	--3971
		x"48",	--3972
		x"49",	--3973
		x"12",	--3974
		x"c0",	--3975
		x"4e",	--3976
		x"4f",	--3977
		x"43",	--3978
		x"43",	--3979
		x"3c",	--3980
		x"4a",	--3981
		x"4b",	--3982
		x"43",	--3983
		x"40",	--3984
		x"bf",	--3985
		x"12",	--3986
		x"c0",	--3987
		x"4e",	--3988
		x"4f",	--3989
		x"40",	--3990
		x"00",	--3991
		x"43",	--3992
		x"3c",	--3993
		x"43",	--3994
		x"40",	--3995
		x"3f",	--3996
		x"4a",	--3997
		x"4b",	--3998
		x"12",	--3999
		x"be",	--4000
		x"4e",	--4001
		x"4f",	--4002
		x"43",	--4003
		x"40",	--4004
		x"3f",	--4005
		x"4a",	--4006
		x"4b",	--4007
		x"12",	--4008
		x"be",	--4009
		x"43",	--4010
		x"40",	--4011
		x"3f",	--4012
		x"12",	--4013
		x"bd",	--4014
		x"4e",	--4015
		x"4f",	--4016
		x"48",	--4017
		x"49",	--4018
		x"12",	--4019
		x"c0",	--4020
		x"4e",	--4021
		x"4f",	--4022
		x"43",	--4023
		x"43",	--4024
		x"44",	--4025
		x"45",	--4026
		x"44",	--4027
		x"45",	--4028
		x"12",	--4029
		x"be",	--4030
		x"4e",	--4031
		x"4f",	--4032
		x"4e",	--4033
		x"4f",	--4034
		x"12",	--4035
		x"be",	--4036
		x"4e",	--4037
		x"4f",	--4038
		x"40",	--4039
		x"69",	--4040
		x"40",	--4041
		x"3c",	--4042
		x"12",	--4043
		x"be",	--4044
		x"40",	--4045
		x"da",	--4046
		x"40",	--4047
		x"3d",	--4048
		x"12",	--4049
		x"bd",	--4050
		x"4e",	--4051
		x"4f",	--4052
		x"4a",	--4053
		x"4b",	--4054
		x"12",	--4055
		x"be",	--4056
		x"40",	--4057
		x"6b",	--4058
		x"40",	--4059
		x"3d",	--4060
		x"12",	--4061
		x"bd",	--4062
		x"4e",	--4063
		x"4f",	--4064
		x"4a",	--4065
		x"4b",	--4066
		x"12",	--4067
		x"be",	--4068
		x"40",	--4069
		x"2e",	--4070
		x"40",	--4071
		x"3d",	--4072
		x"12",	--4073
		x"bd",	--4074
		x"4e",	--4075
		x"4f",	--4076
		x"4a",	--4077
		x"4b",	--4078
		x"12",	--4079
		x"be",	--4080
		x"40",	--4081
		x"49",	--4082
		x"40",	--4083
		x"3e",	--4084
		x"12",	--4085
		x"bd",	--4086
		x"4e",	--4087
		x"4f",	--4088
		x"4a",	--4089
		x"4b",	--4090
		x"12",	--4091
		x"be",	--4092
		x"40",	--4093
		x"aa",	--4094
		x"40",	--4095
		x"3e",	--4096
		x"12",	--4097
		x"bd",	--4098
		x"4e",	--4099
		x"4f",	--4100
		x"48",	--4101
		x"49",	--4102
		x"12",	--4103
		x"be",	--4104
		x"4e",	--4105
		x"00",	--4106
		x"4f",	--4107
		x"00",	--4108
		x"40",	--4109
		x"a2",	--4110
		x"40",	--4111
		x"bd",	--4112
		x"4a",	--4113
		x"4b",	--4114
		x"12",	--4115
		x"be",	--4116
		x"40",	--4117
		x"f1",	--4118
		x"40",	--4119
		x"3d",	--4120
		x"12",	--4121
		x"be",	--4122
		x"4e",	--4123
		x"4f",	--4124
		x"4a",	--4125
		x"4b",	--4126
		x"12",	--4127
		x"be",	--4128
		x"40",	--4129
		x"87",	--4130
		x"40",	--4131
		x"3d",	--4132
		x"12",	--4133
		x"be",	--4134
		x"4e",	--4135
		x"4f",	--4136
		x"4a",	--4137
		x"4b",	--4138
		x"12",	--4139
		x"be",	--4140
		x"40",	--4141
		x"8e",	--4142
		x"40",	--4143
		x"3d",	--4144
		x"12",	--4145
		x"be",	--4146
		x"4e",	--4147
		x"4f",	--4148
		x"4a",	--4149
		x"4b",	--4150
		x"12",	--4151
		x"be",	--4152
		x"40",	--4153
		x"cc",	--4154
		x"40",	--4155
		x"3e",	--4156
		x"12",	--4157
		x"be",	--4158
		x"4e",	--4159
		x"4f",	--4160
		x"4a",	--4161
		x"4b",	--4162
		x"12",	--4163
		x"be",	--4164
		x"4e",	--4165
		x"4f",	--4166
		x"93",	--4167
		x"20",	--4168
		x"93",	--4169
		x"20",	--4170
		x"4e",	--4171
		x"4f",	--4172
		x"41",	--4173
		x"00",	--4174
		x"41",	--4175
		x"00",	--4176
		x"12",	--4177
		x"bd",	--4178
		x"4e",	--4179
		x"4f",	--4180
		x"44",	--4181
		x"45",	--4182
		x"12",	--4183
		x"be",	--4184
		x"4e",	--4185
		x"4f",	--4186
		x"44",	--4187
		x"45",	--4188
		x"12",	--4189
		x"be",	--4190
		x"4e",	--4191
		x"4f",	--4192
		x"3c",	--4193
		x"46",	--4194
		x"5b",	--4195
		x"5b",	--4196
		x"4b",	--4197
		x"50",	--4198
		x"d8",	--4199
		x"48",	--4200
		x"49",	--4201
		x"41",	--4202
		x"00",	--4203
		x"41",	--4204
		x"00",	--4205
		x"12",	--4206
		x"bd",	--4207
		x"4e",	--4208
		x"4f",	--4209
		x"44",	--4210
		x"45",	--4211
		x"12",	--4212
		x"be",	--4213
		x"4b",	--4214
		x"d8",	--4215
		x"4b",	--4216
		x"d8",	--4217
		x"12",	--4218
		x"be",	--4219
		x"44",	--4220
		x"45",	--4221
		x"12",	--4222
		x"be",	--4223
		x"4e",	--4224
		x"4f",	--4225
		x"47",	--4226
		x"47",	--4227
		x"00",	--4228
		x"12",	--4229
		x"be",	--4230
		x"4e",	--4231
		x"4f",	--4232
		x"93",	--4233
		x"00",	--4234
		x"34",	--4235
		x"e0",	--4236
		x"80",	--4237
		x"3c",	--4238
		x"40",	--4239
		x"0f",	--4240
		x"40",	--4241
		x"bf",	--4242
		x"44",	--4243
		x"45",	--4244
		x"52",	--4245
		x"41",	--4246
		x"41",	--4247
		x"41",	--4248
		x"41",	--4249
		x"41",	--4250
		x"41",	--4251
		x"41",	--4252
		x"41",	--4253
		x"41",	--4254
		x"12",	--4255
		x"9d",	--4256
		x"41",	--4257
		x"12",	--4258
		x"12",	--4259
		x"82",	--4260
		x"4e",	--4261
		x"4f",	--4262
		x"f3",	--4263
		x"f0",	--4264
		x"7f",	--4265
		x"90",	--4266
		x"3f",	--4267
		x"38",	--4268
		x"90",	--4269
		x"3f",	--4270
		x"34",	--4271
		x"90",	--4272
		x"0f",	--4273
		x"2c",	--4274
		x"12",	--4275
		x"43",	--4276
		x"43",	--4277
		x"3c",	--4278
		x"90",	--4279
		x"7f",	--4280
		x"38",	--4281
		x"4e",	--4282
		x"4f",	--4283
		x"12",	--4284
		x"be",	--4285
		x"3c",	--4286
		x"41",	--4287
		x"12",	--4288
		x"a3",	--4289
		x"4e",	--4290
		x"4f",	--4291
		x"f0",	--4292
		x"00",	--4293
		x"f3",	--4294
		x"41",	--4295
		x"00",	--4296
		x"41",	--4297
		x"00",	--4298
		x"41",	--4299
		x"41",	--4300
		x"00",	--4301
		x"93",	--4302
		x"20",	--4303
		x"93",	--4304
		x"24",	--4305
		x"93",	--4306
		x"20",	--4307
		x"93",	--4308
		x"24",	--4309
		x"41",	--4310
		x"41",	--4311
		x"00",	--4312
		x"93",	--4313
		x"20",	--4314
		x"93",	--4315
		x"20",	--4316
		x"12",	--4317
		x"12",	--4318
		x"b6",	--4319
		x"53",	--4320
		x"3c",	--4321
		x"12",	--4322
		x"a1",	--4323
		x"3c",	--4324
		x"12",	--4325
		x"12",	--4326
		x"b6",	--4327
		x"53",	--4328
		x"3c",	--4329
		x"12",	--4330
		x"a1",	--4331
		x"e0",	--4332
		x"80",	--4333
		x"52",	--4334
		x"41",	--4335
		x"41",	--4336
		x"41",	--4337
		x"12",	--4338
		x"a1",	--4339
		x"41",	--4340
		x"12",	--4341
		x"12",	--4342
		x"12",	--4343
		x"12",	--4344
		x"12",	--4345
		x"12",	--4346
		x"12",	--4347
		x"12",	--4348
		x"82",	--4349
		x"4e",	--4350
		x"4f",	--4351
		x"4c",	--4352
		x"4d",	--4353
		x"4e",	--4354
		x"4f",	--4355
		x"f3",	--4356
		x"f0",	--4357
		x"7f",	--4358
		x"90",	--4359
		x"32",	--4360
		x"34",	--4361
		x"12",	--4362
		x"c4",	--4363
		x"93",	--4364
		x"24",	--4365
		x"46",	--4366
		x"47",	--4367
		x"46",	--4368
		x"47",	--4369
		x"12",	--4370
		x"be",	--4371
		x"4e",	--4372
		x"4f",	--4373
		x"40",	--4374
		x"d7",	--4375
		x"40",	--4376
		x"ad",	--4377
		x"12",	--4378
		x"be",	--4379
		x"40",	--4380
		x"74",	--4381
		x"40",	--4382
		x"31",	--4383
		x"12",	--4384
		x"bd",	--4385
		x"4e",	--4386
		x"4f",	--4387
		x"48",	--4388
		x"49",	--4389
		x"12",	--4390
		x"be",	--4391
		x"40",	--4392
		x"f2",	--4393
		x"40",	--4394
		x"34",	--4395
		x"12",	--4396
		x"be",	--4397
		x"4e",	--4398
		x"4f",	--4399
		x"48",	--4400
		x"49",	--4401
		x"12",	--4402
		x"be",	--4403
		x"40",	--4404
		x"0d",	--4405
		x"40",	--4406
		x"37",	--4407
		x"12",	--4408
		x"bd",	--4409
		x"4e",	--4410
		x"4f",	--4411
		x"48",	--4412
		x"49",	--4413
		x"12",	--4414
		x"be",	--4415
		x"40",	--4416
		x"0b",	--4417
		x"40",	--4418
		x"3a",	--4419
		x"12",	--4420
		x"be",	--4421
		x"4e",	--4422
		x"4f",	--4423
		x"48",	--4424
		x"49",	--4425
		x"12",	--4426
		x"be",	--4427
		x"40",	--4428
		x"aa",	--4429
		x"40",	--4430
		x"3d",	--4431
		x"12",	--4432
		x"bd",	--4433
		x"4e",	--4434
		x"4f",	--4435
		x"48",	--4436
		x"49",	--4437
		x"12",	--4438
		x"be",	--4439
		x"4e",	--4440
		x"00",	--4441
		x"4f",	--4442
		x"00",	--4443
		x"90",	--4444
		x"3e",	--4445
		x"38",	--4446
		x"90",	--4447
		x"3e",	--4448
		x"34",	--4449
		x"90",	--4450
		x"99",	--4451
		x"2c",	--4452
		x"43",	--4453
		x"40",	--4454
		x"3f",	--4455
		x"48",	--4456
		x"49",	--4457
		x"12",	--4458
		x"be",	--4459
		x"4e",	--4460
		x"4f",	--4461
		x"41",	--4462
		x"41",	--4463
		x"00",	--4464
		x"48",	--4465
		x"49",	--4466
		x"12",	--4467
		x"be",	--4468
		x"4e",	--4469
		x"4f",	--4470
		x"44",	--4471
		x"45",	--4472
		x"46",	--4473
		x"47",	--4474
		x"12",	--4475
		x"be",	--4476
		x"4e",	--4477
		x"4f",	--4478
		x"48",	--4479
		x"49",	--4480
		x"12",	--4481
		x"be",	--4482
		x"4e",	--4483
		x"4f",	--4484
		x"4a",	--4485
		x"4b",	--4486
		x"12",	--4487
		x"be",	--4488
		x"4e",	--4489
		x"4f",	--4490
		x"43",	--4491
		x"40",	--4492
		x"3f",	--4493
		x"3c",	--4494
		x"90",	--4495
		x"3f",	--4496
		x"38",	--4497
		x"90",	--4498
		x"3f",	--4499
		x"34",	--4500
		x"93",	--4501
		x"2c",	--4502
		x"53",	--4503
		x"60",	--4504
		x"ff",	--4505
		x"3c",	--4506
		x"43",	--4507
		x"40",	--4508
		x"3e",	--4509
		x"4a",	--4510
		x"4b",	--4511
		x"43",	--4512
		x"40",	--4513
		x"3f",	--4514
		x"12",	--4515
		x"be",	--4516
		x"4e",	--4517
		x"00",	--4518
		x"4f",	--4519
		x"00",	--4520
		x"43",	--4521
		x"40",	--4522
		x"3f",	--4523
		x"48",	--4524
		x"49",	--4525
		x"12",	--4526
		x"be",	--4527
		x"4a",	--4528
		x"4b",	--4529
		x"12",	--4530
		x"be",	--4531
		x"4e",	--4532
		x"4f",	--4533
		x"41",	--4534
		x"41",	--4535
		x"00",	--4536
		x"48",	--4537
		x"49",	--4538
		x"12",	--4539
		x"be",	--4540
		x"4e",	--4541
		x"4f",	--4542
		x"44",	--4543
		x"45",	--4544
		x"46",	--4545
		x"47",	--4546
		x"12",	--4547
		x"be",	--4548
		x"4e",	--4549
		x"4f",	--4550
		x"48",	--4551
		x"49",	--4552
		x"12",	--4553
		x"be",	--4554
		x"4e",	--4555
		x"4f",	--4556
		x"4a",	--4557
		x"4b",	--4558
		x"12",	--4559
		x"be",	--4560
		x"4e",	--4561
		x"4f",	--4562
		x"41",	--4563
		x"00",	--4564
		x"41",	--4565
		x"00",	--4566
		x"12",	--4567
		x"be",	--4568
		x"3c",	--4569
		x"43",	--4570
		x"40",	--4571
		x"3f",	--4572
		x"52",	--4573
		x"41",	--4574
		x"41",	--4575
		x"41",	--4576
		x"41",	--4577
		x"41",	--4578
		x"41",	--4579
		x"41",	--4580
		x"41",	--4581
		x"41",	--4582
		x"12",	--4583
		x"12",	--4584
		x"12",	--4585
		x"12",	--4586
		x"12",	--4587
		x"12",	--4588
		x"12",	--4589
		x"12",	--4590
		x"50",	--4591
		x"ff",	--4592
		x"4d",	--4593
		x"00",	--4594
		x"4e",	--4595
		x"00",	--4596
		x"4f",	--4597
		x"00",	--4598
		x"4e",	--4599
		x"4f",	--4600
		x"f3",	--4601
		x"f0",	--4602
		x"7f",	--4603
		x"90",	--4604
		x"3f",	--4605
		x"38",	--4606
		x"90",	--4607
		x"3f",	--4608
		x"34",	--4609
		x"90",	--4610
		x"0f",	--4611
		x"2c",	--4612
		x"41",	--4613
		x"00",	--4614
		x"4e",	--4615
		x"00",	--4616
		x"4f",	--4617
		x"00",	--4618
		x"43",	--4619
		x"00",	--4620
		x"43",	--4621
		x"00",	--4622
		x"40",	--4623
		x"a8",	--4624
		x"90",	--4625
		x"40",	--4626
		x"38",	--4627
		x"90",	--4628
		x"40",	--4629
		x"34",	--4630
		x"90",	--4631
		x"cb",	--4632
		x"2c",	--4633
		x"93",	--4634
		x"00",	--4635
		x"38",	--4636
		x"20",	--4637
		x"93",	--4638
		x"00",	--4639
		x"28",	--4640
		x"40",	--4641
		x"0f",	--4642
		x"40",	--4643
		x"3f",	--4644
		x"12",	--4645
		x"be",	--4646
		x"4e",	--4647
		x"4f",	--4648
		x"f0",	--4649
		x"ff",	--4650
		x"f3",	--4651
		x"90",	--4652
		x"0f",	--4653
		x"20",	--4654
		x"90",	--4655
		x"3f",	--4656
		x"24",	--4657
		x"40",	--4658
		x"44",	--4659
		x"40",	--4660
		x"37",	--4661
		x"48",	--4662
		x"49",	--4663
		x"12",	--4664
		x"be",	--4665
		x"4e",	--4666
		x"4f",	--4667
		x"41",	--4668
		x"00",	--4669
		x"4c",	--4670
		x"00",	--4671
		x"4d",	--4672
		x"00",	--4673
		x"48",	--4674
		x"49",	--4675
		x"12",	--4676
		x"be",	--4677
		x"40",	--4678
		x"44",	--4679
		x"40",	--4680
		x"37",	--4681
		x"3c",	--4682
		x"40",	--4683
		x"44",	--4684
		x"40",	--4685
		x"37",	--4686
		x"12",	--4687
		x"be",	--4688
		x"4e",	--4689
		x"4f",	--4690
		x"40",	--4691
		x"a3",	--4692
		x"40",	--4693
		x"2e",	--4694
		x"12",	--4695
		x"be",	--4696
		x"4e",	--4697
		x"4f",	--4698
		x"41",	--4699
		x"00",	--4700
		x"4c",	--4701
		x"00",	--4702
		x"4d",	--4703
		x"00",	--4704
		x"4a",	--4705
		x"4b",	--4706
		x"12",	--4707
		x"be",	--4708
		x"40",	--4709
		x"a3",	--4710
		x"40",	--4711
		x"2e",	--4712
		x"12",	--4713
		x"be",	--4714
		x"41",	--4715
		x"00",	--4716
		x"4e",	--4717
		x"00",	--4718
		x"4f",	--4719
		x"00",	--4720
		x"43",	--4721
		x"43",	--4722
		x"40",	--4723
		x"a9",	--4724
		x"40",	--4725
		x"0f",	--4726
		x"40",	--4727
		x"3f",	--4728
		x"12",	--4729
		x"bd",	--4730
		x"4e",	--4731
		x"4f",	--4732
		x"f0",	--4733
		x"ff",	--4734
		x"f3",	--4735
		x"90",	--4736
		x"0f",	--4737
		x"20",	--4738
		x"90",	--4739
		x"3f",	--4740
		x"24",	--4741
		x"40",	--4742
		x"44",	--4743
		x"40",	--4744
		x"37",	--4745
		x"48",	--4746
		x"49",	--4747
		x"12",	--4748
		x"bd",	--4749
		x"4e",	--4750
		x"4f",	--4751
		x"41",	--4752
		x"00",	--4753
		x"4c",	--4754
		x"00",	--4755
		x"4d",	--4756
		x"00",	--4757
		x"48",	--4758
		x"49",	--4759
		x"12",	--4760
		x"be",	--4761
		x"40",	--4762
		x"44",	--4763
		x"40",	--4764
		x"37",	--4765
		x"3c",	--4766
		x"40",	--4767
		x"44",	--4768
		x"40",	--4769
		x"37",	--4770
		x"12",	--4771
		x"bd",	--4772
		x"4e",	--4773
		x"4f",	--4774
		x"40",	--4775
		x"a3",	--4776
		x"40",	--4777
		x"2e",	--4778
		x"12",	--4779
		x"bd",	--4780
		x"4e",	--4781
		x"4f",	--4782
		x"41",	--4783
		x"00",	--4784
		x"4c",	--4785
		x"00",	--4786
		x"4d",	--4787
		x"00",	--4788
		x"4a",	--4789
		x"4b",	--4790
		x"12",	--4791
		x"be",	--4792
		x"40",	--4793
		x"a3",	--4794
		x"40",	--4795
		x"2e",	--4796
		x"12",	--4797
		x"bd",	--4798
		x"41",	--4799
		x"00",	--4800
		x"4e",	--4801
		x"00",	--4802
		x"4f",	--4803
		x"00",	--4804
		x"43",	--4805
		x"43",	--4806
		x"40",	--4807
		x"a9",	--4808
		x"90",	--4809
		x"43",	--4810
		x"38",	--4811
		x"90",	--4812
		x"43",	--4813
		x"38",	--4814
		x"40",	--4815
		x"a8",	--4816
		x"90",	--4817
		x"0f",	--4818
		x"28",	--4819
		x"40",	--4820
		x"a8",	--4821
		x"4e",	--4822
		x"4f",	--4823
		x"f0",	--4824
		x"7f",	--4825
		x"40",	--4826
		x"f9",	--4827
		x"40",	--4828
		x"3f",	--4829
		x"48",	--4830
		x"49",	--4831
		x"12",	--4832
		x"be",	--4833
		x"43",	--4834
		x"40",	--4835
		x"3f",	--4836
		x"12",	--4837
		x"bd",	--4838
		x"12",	--4839
		x"c4",	--4840
		x"4e",	--4841
		x"4f",	--4842
		x"12",	--4843
		x"c3",	--4844
		x"4e",	--4845
		x"00",	--4846
		x"4f",	--4847
		x"00",	--4848
		x"40",	--4849
		x"0f",	--4850
		x"40",	--4851
		x"3f",	--4852
		x"12",	--4853
		x"be",	--4854
		x"4e",	--4855
		x"4f",	--4856
		x"48",	--4857
		x"49",	--4858
		x"12",	--4859
		x"be",	--4860
		x"4e",	--4861
		x"4f",	--4862
		x"40",	--4863
		x"44",	--4864
		x"40",	--4865
		x"37",	--4866
		x"41",	--4867
		x"00",	--4868
		x"41",	--4869
		x"00",	--4870
		x"12",	--4871
		x"be",	--4872
		x"4e",	--4873
		x"00",	--4874
		x"4f",	--4875
		x"00",	--4876
		x"93",	--4877
		x"38",	--4878
		x"93",	--4879
		x"34",	--4880
		x"90",	--4881
		x"00",	--4882
		x"2c",	--4883
		x"4a",	--4884
		x"4b",	--4885
		x"f0",	--4886
		x"ff",	--4887
		x"f3",	--4888
		x"46",	--4889
		x"53",	--4890
		x"5f",	--4891
		x"5f",	--4892
		x"50",	--4893
		x"d8",	--4894
		x"9f",	--4895
		x"20",	--4896
		x"9f",	--4897
		x"00",	--4898
		x"24",	--4899
		x"41",	--4900
		x"00",	--4901
		x"41",	--4902
		x"00",	--4903
		x"40",	--4904
		x"a8",	--4905
		x"41",	--4906
		x"00",	--4907
		x"41",	--4908
		x"00",	--4909
		x"44",	--4910
		x"45",	--4911
		x"12",	--4912
		x"be",	--4913
		x"4e",	--4914
		x"4f",	--4915
		x"41",	--4916
		x"00",	--4917
		x"48",	--4918
		x"00",	--4919
		x"49",	--4920
		x"00",	--4921
		x"4b",	--4922
		x"00",	--4923
		x"4b",	--4924
		x"10",	--4925
		x"11",	--4926
		x"10",	--4927
		x"11",	--4928
		x"4d",	--4929
		x"00",	--4930
		x"40",	--4931
		x"00",	--4932
		x"4f",	--4933
		x"41",	--4934
		x"00",	--4935
		x"41",	--4936
		x"00",	--4937
		x"11",	--4938
		x"10",	--4939
		x"53",	--4940
		x"23",	--4941
		x"4e",	--4942
		x"00",	--4943
		x"4f",	--4944
		x"00",	--4945
		x"4c",	--4946
		x"43",	--4947
		x"40",	--4948
		x"00",	--4949
		x"c3",	--4950
		x"10",	--4951
		x"10",	--4952
		x"53",	--4953
		x"23",	--4954
		x"f0",	--4955
		x"00",	--4956
		x"f3",	--4957
		x"41",	--4958
		x"00",	--4959
		x"41",	--4960
		x"00",	--4961
		x"8a",	--4962
		x"7b",	--4963
		x"93",	--4964
		x"38",	--4965
		x"20",	--4966
		x"90",	--4967
		x"00",	--4968
		x"28",	--4969
		x"40",	--4970
		x"44",	--4971
		x"40",	--4972
		x"37",	--4973
		x"41",	--4974
		x"00",	--4975
		x"41",	--4976
		x"00",	--4977
		x"12",	--4978
		x"be",	--4979
		x"4e",	--4980
		x"4f",	--4981
		x"4e",	--4982
		x"4f",	--4983
		x"44",	--4984
		x"45",	--4985
		x"12",	--4986
		x"be",	--4987
		x"4e",	--4988
		x"00",	--4989
		x"4f",	--4990
		x"00",	--4991
		x"4e",	--4992
		x"4f",	--4993
		x"44",	--4994
		x"45",	--4995
		x"12",	--4996
		x"be",	--4997
		x"48",	--4998
		x"49",	--4999
		x"12",	--5000
		x"be",	--5001
		x"4e",	--5002
		x"4f",	--5003
		x"40",	--5004
		x"a3",	--5005
		x"40",	--5006
		x"2e",	--5007
		x"41",	--5008
		x"00",	--5009
		x"41",	--5010
		x"00",	--5011
		x"12",	--5012
		x"be",	--5013
		x"48",	--5014
		x"49",	--5015
		x"12",	--5016
		x"be",	--5017
		x"4e",	--5018
		x"00",	--5019
		x"4f",	--5020
		x"00",	--5021
		x"4e",	--5022
		x"4f",	--5023
		x"41",	--5024
		x"00",	--5025
		x"41",	--5026
		x"00",	--5027
		x"12",	--5028
		x"be",	--5029
		x"4e",	--5030
		x"4f",	--5031
		x"41",	--5032
		x"00",	--5033
		x"4a",	--5034
		x"00",	--5035
		x"4b",	--5036
		x"00",	--5037
		x"4f",	--5038
		x"43",	--5039
		x"40",	--5040
		x"00",	--5041
		x"c3",	--5042
		x"10",	--5043
		x"10",	--5044
		x"53",	--5045
		x"23",	--5046
		x"f0",	--5047
		x"00",	--5048
		x"f3",	--5049
		x"41",	--5050
		x"00",	--5051
		x"41",	--5052
		x"00",	--5053
		x"8a",	--5054
		x"7b",	--5055
		x"4d",	--5056
		x"4e",	--5057
		x"93",	--5058
		x"38",	--5059
		x"20",	--5060
		x"90",	--5061
		x"00",	--5062
		x"28",	--5063
		x"40",	--5064
		x"a3",	--5065
		x"40",	--5066
		x"2e",	--5067
		x"41",	--5068
		x"00",	--5069
		x"41",	--5070
		x"00",	--5071
		x"12",	--5072
		x"be",	--5073
		x"4e",	--5074
		x"4f",	--5075
		x"4e",	--5076
		x"4f",	--5077
		x"41",	--5078
		x"00",	--5079
		x"41",	--5080
		x"00",	--5081
		x"12",	--5082
		x"be",	--5083
		x"4e",	--5084
		x"4f",	--5085
		x"4e",	--5086
		x"4f",	--5087
		x"41",	--5088
		x"00",	--5089
		x"41",	--5090
		x"00",	--5091
		x"12",	--5092
		x"be",	--5093
		x"4a",	--5094
		x"4b",	--5095
		x"12",	--5096
		x"be",	--5097
		x"4e",	--5098
		x"4f",	--5099
		x"40",	--5100
		x"31",	--5101
		x"40",	--5102
		x"24",	--5103
		x"41",	--5104
		x"00",	--5105
		x"41",	--5106
		x"00",	--5107
		x"12",	--5108
		x"be",	--5109
		x"4a",	--5110
		x"4b",	--5111
		x"12",	--5112
		x"be",	--5113
		x"4e",	--5114
		x"00",	--5115
		x"4f",	--5116
		x"00",	--5117
		x"4e",	--5118
		x"4f",	--5119
		x"44",	--5120
		x"45",	--5121
		x"12",	--5122
		x"be",	--5123
		x"41",	--5124
		x"00",	--5125
		x"4e",	--5126
		x"00",	--5127
		x"4f",	--5128
		x"00",	--5129
		x"3c",	--5130
		x"41",	--5131
		x"00",	--5132
		x"41",	--5133
		x"00",	--5134
		x"41",	--5135
		x"00",	--5136
		x"4e",	--5137
		x"4e",	--5138
		x"00",	--5139
		x"48",	--5140
		x"49",	--5141
		x"44",	--5142
		x"45",	--5143
		x"12",	--5144
		x"be",	--5145
		x"41",	--5146
		x"00",	--5147
		x"41",	--5148
		x"00",	--5149
		x"12",	--5150
		x"be",	--5151
		x"4e",	--5152
		x"4f",	--5153
		x"41",	--5154
		x"00",	--5155
		x"4a",	--5156
		x"00",	--5157
		x"4b",	--5158
		x"00",	--5159
		x"93",	--5160
		x"00",	--5161
		x"34",	--5162
		x"48",	--5163
		x"49",	--5164
		x"e0",	--5165
		x"80",	--5166
		x"4d",	--5167
		x"00",	--5168
		x"4e",	--5169
		x"00",	--5170
		x"4a",	--5171
		x"4b",	--5172
		x"e0",	--5173
		x"80",	--5174
		x"4d",	--5175
		x"00",	--5176
		x"4e",	--5177
		x"00",	--5178
		x"3c",	--5179
		x"90",	--5180
		x"7f",	--5181
		x"38",	--5182
		x"4e",	--5183
		x"4f",	--5184
		x"12",	--5185
		x"be",	--5186
		x"41",	--5187
		x"00",	--5188
		x"4e",	--5189
		x"00",	--5190
		x"4f",	--5191
		x"00",	--5192
		x"4e",	--5193
		x"00",	--5194
		x"4f",	--5195
		x"00",	--5196
		x"43",	--5197
		x"43",	--5198
		x"3c",	--5199
		x"4b",	--5200
		x"4b",	--5201
		x"10",	--5202
		x"11",	--5203
		x"10",	--5204
		x"11",	--5205
		x"40",	--5206
		x"00",	--5207
		x"11",	--5208
		x"10",	--5209
		x"53",	--5210
		x"23",	--5211
		x"4c",	--5212
		x"50",	--5213
		x"ff",	--5214
		x"43",	--5215
		x"43",	--5216
		x"49",	--5217
		x"40",	--5218
		x"00",	--5219
		x"5c",	--5220
		x"6d",	--5221
		x"53",	--5222
		x"23",	--5223
		x"8c",	--5224
		x"7d",	--5225
		x"4a",	--5226
		x"4b",	--5227
		x"12",	--5228
		x"c4",	--5229
		x"12",	--5230
		x"c3",	--5231
		x"4e",	--5232
		x"4f",	--5233
		x"4e",	--5234
		x"00",	--5235
		x"4f",	--5236
		x"00",	--5237
		x"4a",	--5238
		x"4b",	--5239
		x"12",	--5240
		x"be",	--5241
		x"43",	--5242
		x"40",	--5243
		x"43",	--5244
		x"12",	--5245
		x"be",	--5246
		x"4e",	--5247
		x"4f",	--5248
		x"12",	--5249
		x"c4",	--5250
		x"12",	--5251
		x"c3",	--5252
		x"4e",	--5253
		x"4f",	--5254
		x"4e",	--5255
		x"00",	--5256
		x"4f",	--5257
		x"00",	--5258
		x"4a",	--5259
		x"4b",	--5260
		x"12",	--5261
		x"be",	--5262
		x"43",	--5263
		x"40",	--5264
		x"43",	--5265
		x"12",	--5266
		x"be",	--5267
		x"4e",	--5268
		x"00",	--5269
		x"4f",	--5270
		x"00",	--5271
		x"41",	--5272
		x"52",	--5273
		x"40",	--5274
		x"00",	--5275
		x"3c",	--5276
		x"53",	--5277
		x"82",	--5278
		x"43",	--5279
		x"43",	--5280
		x"48",	--5281
		x"00",	--5282
		x"48",	--5283
		x"00",	--5284
		x"12",	--5285
		x"c1",	--5286
		x"93",	--5287
		x"27",	--5288
		x"12",	--5289
		x"d8",	--5290
		x"12",	--5291
		x"4a",	--5292
		x"49",	--5293
		x"41",	--5294
		x"00",	--5295
		x"41",	--5296
		x"52",	--5297
		x"12",	--5298
		x"a9",	--5299
		x"52",	--5300
		x"4f",	--5301
		x"10",	--5302
		x"11",	--5303
		x"10",	--5304
		x"11",	--5305
		x"4f",	--5306
		x"93",	--5307
		x"00",	--5308
		x"34",	--5309
		x"41",	--5310
		x"00",	--5311
		x"e0",	--5312
		x"80",	--5313
		x"00",	--5314
		x"e0",	--5315
		x"80",	--5316
		x"00",	--5317
		x"e3",	--5318
		x"e3",	--5319
		x"53",	--5320
		x"63",	--5321
		x"46",	--5322
		x"47",	--5323
		x"50",	--5324
		x"00",	--5325
		x"41",	--5326
		x"41",	--5327
		x"41",	--5328
		x"41",	--5329
		x"41",	--5330
		x"41",	--5331
		x"41",	--5332
		x"41",	--5333
		x"41",	--5334
		x"12",	--5335
		x"12",	--5336
		x"12",	--5337
		x"12",	--5338
		x"12",	--5339
		x"12",	--5340
		x"12",	--5341
		x"12",	--5342
		x"50",	--5343
		x"fe",	--5344
		x"4f",	--5345
		x"01",	--5346
		x"4e",	--5347
		x"01",	--5348
		x"4c",	--5349
		x"01",	--5350
		x"41",	--5351
		x"01",	--5352
		x"5a",	--5353
		x"43",	--5354
		x"01",	--5355
		x"43",	--5356
		x"01",	--5357
		x"4a",	--5358
		x"dc",	--5359
		x"01",	--5360
		x"41",	--5361
		x"01",	--5362
		x"10",	--5363
		x"11",	--5364
		x"10",	--5365
		x"11",	--5366
		x"4a",	--5367
		x"01",	--5368
		x"4c",	--5369
		x"53",	--5370
		x"4a",	--5371
		x"01",	--5372
		x"10",	--5373
		x"11",	--5374
		x"10",	--5375
		x"11",	--5376
		x"4a",	--5377
		x"01",	--5378
		x"4d",	--5379
		x"50",	--5380
		x"ff",	--5381
		x"93",	--5382
		x"34",	--5383
		x"50",	--5384
		x"00",	--5385
		x"11",	--5386
		x"11",	--5387
		x"11",	--5388
		x"4a",	--5389
		x"10",	--5390
		x"11",	--5391
		x"10",	--5392
		x"11",	--5393
		x"4a",	--5394
		x"01",	--5395
		x"48",	--5396
		x"01",	--5397
		x"34",	--5398
		x"43",	--5399
		x"01",	--5400
		x"43",	--5401
		x"01",	--5402
		x"4d",	--5403
		x"10",	--5404
		x"11",	--5405
		x"10",	--5406
		x"11",	--5407
		x"4d",	--5408
		x"41",	--5409
		x"01",	--5410
		x"41",	--5411
		x"01",	--5412
		x"e3",	--5413
		x"e3",	--5414
		x"5a",	--5415
		x"6b",	--5416
		x"5a",	--5417
		x"6b",	--5418
		x"5a",	--5419
		x"6b",	--5420
		x"48",	--5421
		x"49",	--5422
		x"5a",	--5423
		x"6b",	--5424
		x"4d",	--5425
		x"01",	--5426
		x"4e",	--5427
		x"01",	--5428
		x"41",	--5429
		x"01",	--5430
		x"41",	--5431
		x"01",	--5432
		x"81",	--5433
		x"01",	--5434
		x"71",	--5435
		x"01",	--5436
		x"48",	--5437
		x"01",	--5438
		x"49",	--5439
		x"01",	--5440
		x"41",	--5441
		x"01",	--5442
		x"41",	--5443
		x"01",	--5444
		x"51",	--5445
		x"01",	--5446
		x"61",	--5447
		x"01",	--5448
		x"43",	--5449
		x"43",	--5450
		x"43",	--5451
		x"3c",	--5452
		x"41",	--5453
		x"01",	--5454
		x"41",	--5455
		x"01",	--5456
		x"56",	--5457
		x"67",	--5458
		x"93",	--5459
		x"38",	--5460
		x"41",	--5461
		x"01",	--5462
		x"5f",	--5463
		x"5f",	--5464
		x"51",	--5465
		x"01",	--5466
		x"59",	--5467
		x"4f",	--5468
		x"4f",	--5469
		x"00",	--5470
		x"12",	--5471
		x"c3",	--5472
		x"3c",	--5473
		x"43",	--5474
		x"43",	--5475
		x"40",	--5476
		x"00",	--5477
		x"51",	--5478
		x"59",	--5479
		x"4e",	--5480
		x"00",	--5481
		x"4f",	--5482
		x"00",	--5483
		x"53",	--5484
		x"63",	--5485
		x"52",	--5486
		x"97",	--5487
		x"38",	--5488
		x"95",	--5489
		x"3b",	--5490
		x"96",	--5491
		x"2f",	--5492
		x"43",	--5493
		x"01",	--5494
		x"43",	--5495
		x"01",	--5496
		x"41",	--5497
		x"3c",	--5498
		x"41",	--5499
		x"01",	--5500
		x"53",	--5501
		x"5f",	--5502
		x"5f",	--5503
		x"50",	--5504
		x"00",	--5505
		x"54",	--5506
		x"55",	--5507
		x"4f",	--5508
		x"4f",	--5509
		x"00",	--5510
		x"47",	--5511
		x"47",	--5512
		x"12",	--5513
		x"be",	--5514
		x"4e",	--5515
		x"4f",	--5516
		x"4a",	--5517
		x"4b",	--5518
		x"12",	--5519
		x"bd",	--5520
		x"4e",	--5521
		x"4f",	--5522
		x"53",	--5523
		x"63",	--5524
		x"82",	--5525
		x"99",	--5526
		x"01",	--5527
		x"38",	--5528
		x"91",	--5529
		x"01",	--5530
		x"3b",	--5531
		x"98",	--5532
		x"01",	--5533
		x"2f",	--5534
		x"4a",	--5535
		x"00",	--5536
		x"4b",	--5537
		x"00",	--5538
		x"53",	--5539
		x"01",	--5540
		x"63",	--5541
		x"01",	--5542
		x"52",	--5543
		x"91",	--5544
		x"01",	--5545
		x"01",	--5546
		x"38",	--5547
		x"91",	--5548
		x"01",	--5549
		x"01",	--5550
		x"38",	--5551
		x"91",	--5552
		x"01",	--5553
		x"01",	--5554
		x"2c",	--5555
		x"41",	--5556
		x"01",	--5557
		x"01",	--5558
		x"41",	--5559
		x"01",	--5560
		x"01",	--5561
		x"41",	--5562
		x"01",	--5563
		x"41",	--5564
		x"01",	--5565
		x"53",	--5566
		x"63",	--5567
		x"49",	--5568
		x"01",	--5569
		x"4a",	--5570
		x"01",	--5571
		x"3c",	--5572
		x"41",	--5573
		x"01",	--5574
		x"43",	--5575
		x"43",	--5576
		x"43",	--5577
		x"43",	--5578
		x"43",	--5579
		x"3f",	--5580
		x"41",	--5581
		x"01",	--5582
		x"5f",	--5583
		x"5f",	--5584
		x"51",	--5585
		x"4f",	--5586
		x"4f",	--5587
		x"00",	--5588
		x"41",	--5589
		x"50",	--5590
		x"00",	--5591
		x"4a",	--5592
		x"01",	--5593
		x"41",	--5594
		x"01",	--5595
		x"41",	--5596
		x"01",	--5597
		x"43",	--5598
		x"01",	--5599
		x"46",	--5600
		x"47",	--5601
		x"53",	--5602
		x"63",	--5603
		x"44",	--5604
		x"01",	--5605
		x"45",	--5606
		x"01",	--5607
		x"4a",	--5608
		x"3c",	--5609
		x"43",	--5610
		x"40",	--5611
		x"3b",	--5612
		x"48",	--5613
		x"49",	--5614
		x"12",	--5615
		x"be",	--5616
		x"12",	--5617
		x"c4",	--5618
		x"12",	--5619
		x"c3",	--5620
		x"4e",	--5621
		x"4f",	--5622
		x"43",	--5623
		x"40",	--5624
		x"43",	--5625
		x"12",	--5626
		x"be",	--5627
		x"4e",	--5628
		x"4f",	--5629
		x"48",	--5630
		x"49",	--5631
		x"12",	--5632
		x"be",	--5633
		x"12",	--5634
		x"c4",	--5635
		x"4e",	--5636
		x"00",	--5637
		x"4f",	--5638
		x"00",	--5639
		x"41",	--5640
		x"01",	--5641
		x"5f",	--5642
		x"5f",	--5643
		x"51",	--5644
		x"51",	--5645
		x"01",	--5646
		x"4f",	--5647
		x"00",	--5648
		x"4f",	--5649
		x"00",	--5650
		x"4a",	--5651
		x"4b",	--5652
		x"12",	--5653
		x"bd",	--5654
		x"4e",	--5655
		x"4f",	--5656
		x"53",	--5657
		x"63",	--5658
		x"52",	--5659
		x"82",	--5660
		x"01",	--5661
		x"93",	--5662
		x"38",	--5663
		x"93",	--5664
		x"37",	--5665
		x"93",	--5666
		x"2f",	--5667
		x"41",	--5668
		x"01",	--5669
		x"01",	--5670
		x"41",	--5671
		x"01",	--5672
		x"48",	--5673
		x"49",	--5674
		x"12",	--5675
		x"b8",	--5676
		x"4e",	--5677
		x"4f",	--5678
		x"43",	--5679
		x"40",	--5680
		x"3e",	--5681
		x"12",	--5682
		x"be",	--5683
		x"12",	--5684
		x"b9",	--5685
		x"43",	--5686
		x"40",	--5687
		x"41",	--5688
		x"12",	--5689
		x"be",	--5690
		x"4e",	--5691
		x"4f",	--5692
		x"4a",	--5693
		x"4b",	--5694
		x"12",	--5695
		x"be",	--5696
		x"4e",	--5697
		x"4f",	--5698
		x"12",	--5699
		x"c4",	--5700
		x"4e",	--5701
		x"01",	--5702
		x"4f",	--5703
		x"01",	--5704
		x"12",	--5705
		x"c3",	--5706
		x"4e",	--5707
		x"4f",	--5708
		x"4a",	--5709
		x"4b",	--5710
		x"12",	--5711
		x"be",	--5712
		x"4e",	--5713
		x"01",	--5714
		x"4f",	--5715
		x"01",	--5716
		x"93",	--5717
		x"01",	--5718
		x"38",	--5719
		x"20",	--5720
		x"93",	--5721
		x"01",	--5722
		x"28",	--5723
		x"41",	--5724
		x"01",	--5725
		x"41",	--5726
		x"01",	--5727
		x"53",	--5728
		x"63",	--5729
		x"4c",	--5730
		x"5b",	--5731
		x"5b",	--5732
		x"51",	--5733
		x"4b",	--5734
		x"00",	--5735
		x"4b",	--5736
		x"00",	--5737
		x"41",	--5738
		x"01",	--5739
		x"42",	--5740
		x"8e",	--5741
		x"46",	--5742
		x"47",	--5743
		x"49",	--5744
		x"f0",	--5745
		x"00",	--5746
		x"93",	--5747
		x"24",	--5748
		x"11",	--5749
		x"10",	--5750
		x"53",	--5751
		x"3f",	--5752
		x"5a",	--5753
		x"01",	--5754
		x"6b",	--5755
		x"01",	--5756
		x"f0",	--5757
		x"00",	--5758
		x"93",	--5759
		x"24",	--5760
		x"5a",	--5761
		x"6b",	--5762
		x"53",	--5763
		x"3f",	--5764
		x"46",	--5765
		x"47",	--5766
		x"8a",	--5767
		x"7b",	--5768
		x"4c",	--5769
		x"5f",	--5770
		x"5f",	--5771
		x"51",	--5772
		x"48",	--5773
		x"00",	--5774
		x"49",	--5775
		x"00",	--5776
		x"48",	--5777
		x"49",	--5778
		x"40",	--5779
		x"00",	--5780
		x"8e",	--5781
		x"f0",	--5782
		x"00",	--5783
		x"93",	--5784
		x"24",	--5785
		x"11",	--5786
		x"10",	--5787
		x"53",	--5788
		x"3f",	--5789
		x"93",	--5790
		x"01",	--5791
		x"20",	--5792
		x"93",	--5793
		x"01",	--5794
		x"20",	--5795
		x"41",	--5796
		x"01",	--5797
		x"53",	--5798
		x"5f",	--5799
		x"5f",	--5800
		x"51",	--5801
		x"4f",	--5802
		x"00",	--5803
		x"4f",	--5804
		x"00",	--5805
		x"10",	--5806
		x"10",	--5807
		x"e7",	--5808
		x"e7",	--5809
		x"11",	--5810
		x"3c",	--5811
		x"43",	--5812
		x"40",	--5813
		x"3f",	--5814
		x"41",	--5815
		x"01",	--5816
		x"41",	--5817
		x"01",	--5818
		x"12",	--5819
		x"c2",	--5820
		x"93",	--5821
		x"34",	--5822
		x"43",	--5823
		x"43",	--5824
		x"3c",	--5825
		x"93",	--5826
		x"38",	--5827
		x"20",	--5828
		x"93",	--5829
		x"28",	--5830
		x"3c",	--5831
		x"43",	--5832
		x"43",	--5833
		x"53",	--5834
		x"01",	--5835
		x"63",	--5836
		x"01",	--5837
		x"43",	--5838
		x"43",	--5839
		x"43",	--5840
		x"43",	--5841
		x"41",	--5842
		x"01",	--5843
		x"3c",	--5844
		x"4b",	--5845
		x"4b",	--5846
		x"00",	--5847
		x"93",	--5848
		x"20",	--5849
		x"93",	--5850
		x"20",	--5851
		x"93",	--5852
		x"20",	--5853
		x"93",	--5854
		x"24",	--5855
		x"40",	--5856
		x"01",	--5857
		x"43",	--5858
		x"4e",	--5859
		x"4f",	--5860
		x"8c",	--5861
		x"7d",	--5862
		x"49",	--5863
		x"00",	--5864
		x"4a",	--5865
		x"00",	--5866
		x"3c",	--5867
		x"40",	--5868
		x"00",	--5869
		x"43",	--5870
		x"4e",	--5871
		x"4f",	--5872
		x"8c",	--5873
		x"7d",	--5874
		x"48",	--5875
		x"00",	--5876
		x"49",	--5877
		x"00",	--5878
		x"43",	--5879
		x"43",	--5880
		x"53",	--5881
		x"63",	--5882
		x"52",	--5883
		x"91",	--5884
		x"01",	--5885
		x"3b",	--5886
		x"20",	--5887
		x"91",	--5888
		x"01",	--5889
		x"2b",	--5890
		x"93",	--5891
		x"01",	--5892
		x"38",	--5893
		x"20",	--5894
		x"93",	--5895
		x"01",	--5896
		x"28",	--5897
		x"93",	--5898
		x"01",	--5899
		x"20",	--5900
		x"93",	--5901
		x"01",	--5902
		x"24",	--5903
		x"93",	--5904
		x"01",	--5905
		x"20",	--5906
		x"93",	--5907
		x"01",	--5908
		x"24",	--5909
		x"3c",	--5910
		x"41",	--5911
		x"01",	--5912
		x"53",	--5913
		x"5f",	--5914
		x"5f",	--5915
		x"51",	--5916
		x"f0",	--5917
		x"00",	--5918
		x"00",	--5919
		x"f3",	--5920
		x"00",	--5921
		x"3c",	--5922
		x"41",	--5923
		x"01",	--5924
		x"53",	--5925
		x"5f",	--5926
		x"5f",	--5927
		x"51",	--5928
		x"f0",	--5929
		x"00",	--5930
		x"00",	--5931
		x"f3",	--5932
		x"00",	--5933
		x"93",	--5934
		x"20",	--5935
		x"93",	--5936
		x"20",	--5937
		x"41",	--5938
		x"01",	--5939
		x"41",	--5940
		x"01",	--5941
		x"43",	--5942
		x"40",	--5943
		x"3f",	--5944
		x"12",	--5945
		x"be",	--5946
		x"4e",	--5947
		x"01",	--5948
		x"4f",	--5949
		x"01",	--5950
		x"93",	--5951
		x"20",	--5952
		x"93",	--5953
		x"24",	--5954
		x"41",	--5955
		x"01",	--5956
		x"43",	--5957
		x"40",	--5958
		x"3f",	--5959
		x"12",	--5960
		x"b8",	--5961
		x"4e",	--5962
		x"4f",	--5963
		x"41",	--5964
		x"01",	--5965
		x"41",	--5966
		x"01",	--5967
		x"12",	--5968
		x"be",	--5969
		x"4e",	--5970
		x"01",	--5971
		x"4f",	--5972
		x"01",	--5973
		x"43",	--5974
		x"43",	--5975
		x"41",	--5976
		x"01",	--5977
		x"41",	--5978
		x"01",	--5979
		x"12",	--5980
		x"c1",	--5981
		x"93",	--5982
		x"20",	--5983
		x"41",	--5984
		x"01",	--5985
		x"41",	--5986
		x"01",	--5987
		x"53",	--5988
		x"63",	--5989
		x"41",	--5990
		x"01",	--5991
		x"41",	--5992
		x"01",	--5993
		x"43",	--5994
		x"43",	--5995
		x"01",	--5996
		x"43",	--5997
		x"01",	--5998
		x"3c",	--5999
		x"4a",	--6000
		x"5f",	--6001
		x"5f",	--6002
		x"40",	--6003
		x"00",	--6004
		x"51",	--6005
		x"5e",	--6006
		x"59",	--6007
		x"df",	--6008
		x"00",	--6009
		x"01",	--6010
		x"df",	--6011
		x"00",	--6012
		x"01",	--6013
		x"53",	--6014
		x"63",	--6015
		x"82",	--6016
		x"91",	--6017
		x"01",	--6018
		x"38",	--6019
		x"9d",	--6020
		x"01",	--6021
		x"3b",	--6022
		x"91",	--6023
		x"01",	--6024
		x"2f",	--6025
		x"93",	--6026
		x"01",	--6027
		x"20",	--6028
		x"93",	--6029
		x"01",	--6030
		x"24",	--6031
		x"3c",	--6032
		x"53",	--6033
		x"01",	--6034
		x"63",	--6035
		x"01",	--6036
		x"3c",	--6037
		x"43",	--6038
		x"43",	--6039
		x"01",	--6040
		x"43",	--6041
		x"01",	--6042
		x"82",	--6043
		x"41",	--6044
		x"01",	--6045
		x"5f",	--6046
		x"5f",	--6047
		x"40",	--6048
		x"00",	--6049
		x"51",	--6050
		x"58",	--6051
		x"5e",	--6052
		x"93",	--6053
		x"00",	--6054
		x"20",	--6055
		x"93",	--6056
		x"00",	--6057
		x"27",	--6058
		x"41",	--6059
		x"01",	--6060
		x"41",	--6061
		x"01",	--6062
		x"53",	--6063
		x"63",	--6064
		x"49",	--6065
		x"01",	--6066
		x"4a",	--6067
		x"01",	--6068
		x"43",	--6069
		x"01",	--6070
		x"43",	--6071
		x"49",	--6072
		x"01",	--6073
		x"41",	--6074
		x"01",	--6075
		x"41",	--6076
		x"01",	--6077
		x"59",	--6078
		x"6a",	--6079
		x"4d",	--6080
		x"01",	--6081
		x"4e",	--6082
		x"01",	--6083
		x"49",	--6084
		x"51",	--6085
		x"01",	--6086
		x"48",	--6087
		x"01",	--6088
		x"44",	--6089
		x"3c",	--6090
		x"52",	--6091
		x"01",	--6092
		x"41",	--6093
		x"01",	--6094
		x"5f",	--6095
		x"5f",	--6096
		x"41",	--6097
		x"50",	--6098
		x"00",	--6099
		x"5f",	--6100
		x"41",	--6101
		x"01",	--6102
		x"54",	--6103
		x"41",	--6104
		x"01",	--6105
		x"5f",	--6106
		x"5f",	--6107
		x"51",	--6108
		x"01",	--6109
		x"56",	--6110
		x"4f",	--6111
		x"4f",	--6112
		x"00",	--6113
		x"12",	--6114
		x"c3",	--6115
		x"4e",	--6116
		x"ff",	--6117
		x"4f",	--6118
		x"ff",	--6119
		x"41",	--6120
		x"01",	--6121
		x"41",	--6122
		x"01",	--6123
		x"41",	--6124
		x"01",	--6125
		x"43",	--6126
		x"43",	--6127
		x"43",	--6128
		x"56",	--6129
		x"3c",	--6130
		x"44",	--6131
		x"55",	--6132
		x"4f",	--6133
		x"4f",	--6134
		x"00",	--6135
		x"47",	--6136
		x"47",	--6137
		x"12",	--6138
		x"be",	--6139
		x"4e",	--6140
		x"4f",	--6141
		x"48",	--6142
		x"49",	--6143
		x"12",	--6144
		x"bd",	--6145
		x"4e",	--6146
		x"4f",	--6147
		x"53",	--6148
		x"63",	--6149
		x"82",	--6150
		x"9b",	--6151
		x"01",	--6152
		x"38",	--6153
		x"91",	--6154
		x"01",	--6155
		x"3b",	--6156
		x"9a",	--6157
		x"01",	--6158
		x"2f",	--6159
		x"41",	--6160
		x"01",	--6161
		x"5f",	--6162
		x"5f",	--6163
		x"51",	--6164
		x"51",	--6165
		x"01",	--6166
		x"48",	--6167
		x"ff",	--6168
		x"49",	--6169
		x"ff",	--6170
		x"53",	--6171
		x"01",	--6172
		x"63",	--6173
		x"01",	--6174
		x"52",	--6175
		x"41",	--6176
		x"01",	--6177
		x"41",	--6178
		x"01",	--6179
		x"51",	--6180
		x"01",	--6181
		x"61",	--6182
		x"01",	--6183
		x"91",	--6184
		x"01",	--6185
		x"38",	--6186
		x"9f",	--6187
		x"01",	--6188
		x"3b",	--6189
		x"91",	--6190
		x"01",	--6191
		x"2f",	--6192
		x"4e",	--6193
		x"01",	--6194
		x"4f",	--6195
		x"01",	--6196
		x"40",	--6197
		x"ab",	--6198
		x"46",	--6199
		x"01",	--6200
		x"47",	--6201
		x"01",	--6202
		x"41",	--6203
		x"01",	--6204
		x"e3",	--6205
		x"47",	--6206
		x"53",	--6207
		x"41",	--6208
		x"01",	--6209
		x"41",	--6210
		x"01",	--6211
		x"12",	--6212
		x"b8",	--6213
		x"4e",	--6214
		x"4f",	--6215
		x"43",	--6216
		x"40",	--6217
		x"43",	--6218
		x"12",	--6219
		x"c2",	--6220
		x"93",	--6221
		x"34",	--6222
		x"3c",	--6223
		x"46",	--6224
		x"01",	--6225
		x"47",	--6226
		x"01",	--6227
		x"41",	--6228
		x"01",	--6229
		x"41",	--6230
		x"01",	--6231
		x"53",	--6232
		x"63",	--6233
		x"82",	--6234
		x"01",	--6235
		x"73",	--6236
		x"01",	--6237
		x"46",	--6238
		x"01",	--6239
		x"47",	--6240
		x"01",	--6241
		x"43",	--6242
		x"3c",	--6243
		x"53",	--6244
		x"01",	--6245
		x"63",	--6246
		x"01",	--6247
		x"82",	--6248
		x"01",	--6249
		x"73",	--6250
		x"01",	--6251
		x"82",	--6252
		x"46",	--6253
		x"5f",	--6254
		x"5f",	--6255
		x"40",	--6256
		x"00",	--6257
		x"51",	--6258
		x"59",	--6259
		x"5d",	--6260
		x"93",	--6261
		x"00",	--6262
		x"20",	--6263
		x"93",	--6264
		x"00",	--6265
		x"27",	--6266
		x"3c",	--6267
		x"43",	--6268
		x"40",	--6269
		x"3b",	--6270
		x"46",	--6271
		x"47",	--6272
		x"12",	--6273
		x"be",	--6274
		x"12",	--6275
		x"c4",	--6276
		x"12",	--6277
		x"c3",	--6278
		x"4e",	--6279
		x"4f",	--6280
		x"41",	--6281
		x"01",	--6282
		x"5c",	--6283
		x"5c",	--6284
		x"41",	--6285
		x"5c",	--6286
		x"50",	--6287
		x"00",	--6288
		x"43",	--6289
		x"40",	--6290
		x"43",	--6291
		x"12",	--6292
		x"be",	--6293
		x"4e",	--6294
		x"4f",	--6295
		x"46",	--6296
		x"47",	--6297
		x"12",	--6298
		x"be",	--6299
		x"12",	--6300
		x"c4",	--6301
		x"4e",	--6302
		x"00",	--6303
		x"4f",	--6304
		x"00",	--6305
		x"53",	--6306
		x"01",	--6307
		x"63",	--6308
		x"01",	--6309
		x"52",	--6310
		x"01",	--6311
		x"63",	--6312
		x"01",	--6313
		x"41",	--6314
		x"01",	--6315
		x"5c",	--6316
		x"5c",	--6317
		x"41",	--6318
		x"5c",	--6319
		x"50",	--6320
		x"00",	--6321
		x"44",	--6322
		x"45",	--6323
		x"12",	--6324
		x"c4",	--6325
		x"4e",	--6326
		x"00",	--6327
		x"4f",	--6328
		x"00",	--6329
		x"3c",	--6330
		x"41",	--6331
		x"01",	--6332
		x"5c",	--6333
		x"5c",	--6334
		x"41",	--6335
		x"5c",	--6336
		x"50",	--6337
		x"00",	--6338
		x"46",	--6339
		x"47",	--6340
		x"12",	--6341
		x"c4",	--6342
		x"4e",	--6343
		x"00",	--6344
		x"4f",	--6345
		x"00",	--6346
		x"41",	--6347
		x"01",	--6348
		x"43",	--6349
		x"40",	--6350
		x"3f",	--6351
		x"12",	--6352
		x"b8",	--6353
		x"4e",	--6354
		x"4f",	--6355
		x"41",	--6356
		x"01",	--6357
		x"41",	--6358
		x"01",	--6359
		x"43",	--6360
		x"93",	--6361
		x"38",	--6362
		x"41",	--6363
		x"01",	--6364
		x"5f",	--6365
		x"5f",	--6366
		x"41",	--6367
		x"5f",	--6368
		x"5b",	--6369
		x"40",	--6370
		x"00",	--6371
		x"51",	--6372
		x"5d",	--6373
		x"5b",	--6374
		x"4f",	--6375
		x"4f",	--6376
		x"00",	--6377
		x"12",	--6378
		x"c3",	--6379
		x"4e",	--6380
		x"4f",	--6381
		x"46",	--6382
		x"47",	--6383
		x"12",	--6384
		x"be",	--6385
		x"4e",	--6386
		x"00",	--6387
		x"4f",	--6388
		x"00",	--6389
		x"43",	--6390
		x"40",	--6391
		x"3b",	--6392
		x"46",	--6393
		x"47",	--6394
		x"12",	--6395
		x"be",	--6396
		x"4e",	--6397
		x"4f",	--6398
		x"53",	--6399
		x"63",	--6400
		x"82",	--6401
		x"3f",	--6402
		x"41",	--6403
		x"01",	--6404
		x"01",	--6405
		x"41",	--6406
		x"01",	--6407
		x"01",	--6408
		x"43",	--6409
		x"43",	--6410
		x"43",	--6411
		x"3c",	--6412
		x"41",	--6413
		x"01",	--6414
		x"5f",	--6415
		x"5f",	--6416
		x"51",	--6417
		x"87",	--6418
		x"56",	--6419
		x"4f",	--6420
		x"4f",	--6421
		x"00",	--6422
		x"46",	--6423
		x"dc",	--6424
		x"46",	--6425
		x"dc",	--6426
		x"12",	--6427
		x"be",	--6428
		x"4e",	--6429
		x"4f",	--6430
		x"48",	--6431
		x"49",	--6432
		x"12",	--6433
		x"bd",	--6434
		x"4e",	--6435
		x"4f",	--6436
		x"53",	--6437
		x"63",	--6438
		x"52",	--6439
		x"9b",	--6440
		x"01",	--6441
		x"38",	--6442
		x"20",	--6443
		x"9a",	--6444
		x"01",	--6445
		x"28",	--6446
		x"9b",	--6447
		x"38",	--6448
		x"95",	--6449
		x"3b",	--6450
		x"9a",	--6451
		x"2f",	--6452
		x"40",	--6453
		x"00",	--6454
		x"51",	--6455
		x"57",	--6456
		x"48",	--6457
		x"00",	--6458
		x"49",	--6459
		x"00",	--6460
		x"53",	--6461
		x"01",	--6462
		x"63",	--6463
		x"01",	--6464
		x"52",	--6465
		x"53",	--6466
		x"63",	--6467
		x"93",	--6468
		x"01",	--6469
		x"38",	--6470
		x"43",	--6471
		x"43",	--6472
		x"43",	--6473
		x"43",	--6474
		x"43",	--6475
		x"3f",	--6476
		x"90",	--6477
		x"00",	--6478
		x"01",	--6479
		x"34",	--6480
		x"93",	--6481
		x"01",	--6482
		x"34",	--6483
		x"93",	--6484
		x"01",	--6485
		x"24",	--6486
		x"40",	--6487
		x"b6",	--6488
		x"90",	--6489
		x"00",	--6490
		x"01",	--6491
		x"24",	--6492
		x"40",	--6493
		x"b6",	--6494
		x"3c",	--6495
		x"41",	--6496
		x"01",	--6497
		x"41",	--6498
		x"01",	--6499
		x"43",	--6500
		x"43",	--6501
		x"43",	--6502
		x"93",	--6503
		x"38",	--6504
		x"41",	--6505
		x"01",	--6506
		x"5f",	--6507
		x"5f",	--6508
		x"40",	--6509
		x"00",	--6510
		x"51",	--6511
		x"5e",	--6512
		x"55",	--6513
		x"4f",	--6514
		x"4f",	--6515
		x"00",	--6516
		x"4a",	--6517
		x"4b",	--6518
		x"12",	--6519
		x"bd",	--6520
		x"4e",	--6521
		x"4f",	--6522
		x"53",	--6523
		x"63",	--6524
		x"82",	--6525
		x"3f",	--6526
		x"93",	--6527
		x"01",	--6528
		x"20",	--6529
		x"93",	--6530
		x"01",	--6531
		x"24",	--6532
		x"e0",	--6533
		x"80",	--6534
		x"41",	--6535
		x"01",	--6536
		x"4a",	--6537
		x"00",	--6538
		x"4b",	--6539
		x"00",	--6540
		x"40",	--6541
		x"b6",	--6542
		x"41",	--6543
		x"01",	--6544
		x"41",	--6545
		x"01",	--6546
		x"43",	--6547
		x"43",	--6548
		x"43",	--6549
		x"93",	--6550
		x"38",	--6551
		x"41",	--6552
		x"01",	--6553
		x"5f",	--6554
		x"5f",	--6555
		x"40",	--6556
		x"00",	--6557
		x"51",	--6558
		x"59",	--6559
		x"55",	--6560
		x"4f",	--6561
		x"4f",	--6562
		x"00",	--6563
		x"4a",	--6564
		x"4b",	--6565
		x"12",	--6566
		x"bd",	--6567
		x"4e",	--6568
		x"4f",	--6569
		x"53",	--6570
		x"63",	--6571
		x"82",	--6572
		x"3f",	--6573
		x"4a",	--6574
		x"4b",	--6575
		x"93",	--6576
		x"01",	--6577
		x"20",	--6578
		x"93",	--6579
		x"01",	--6580
		x"24",	--6581
		x"e0",	--6582
		x"80",	--6583
		x"41",	--6584
		x"01",	--6585
		x"4a",	--6586
		x"00",	--6587
		x"4b",	--6588
		x"00",	--6589
		x"41",	--6590
		x"00",	--6591
		x"41",	--6592
		x"00",	--6593
		x"12",	--6594
		x"be",	--6595
		x"41",	--6596
		x"50",	--6597
		x"00",	--6598
		x"43",	--6599
		x"43",	--6600
		x"3c",	--6601
		x"45",	--6602
		x"45",	--6603
		x"12",	--6604
		x"bd",	--6605
		x"53",	--6606
		x"63",	--6607
		x"97",	--6608
		x"01",	--6609
		x"38",	--6610
		x"91",	--6611
		x"01",	--6612
		x"3b",	--6613
		x"96",	--6614
		x"01",	--6615
		x"2f",	--6616
		x"4e",	--6617
		x"4f",	--6618
		x"93",	--6619
		x"01",	--6620
		x"20",	--6621
		x"93",	--6622
		x"01",	--6623
		x"24",	--6624
		x"e0",	--6625
		x"80",	--6626
		x"41",	--6627
		x"01",	--6628
		x"4a",	--6629
		x"00",	--6630
		x"4b",	--6631
		x"00",	--6632
		x"40",	--6633
		x"b6",	--6634
		x"41",	--6635
		x"01",	--6636
		x"5f",	--6637
		x"5f",	--6638
		x"40",	--6639
		x"00",	--6640
		x"51",	--6641
		x"5f",	--6642
		x"51",	--6643
		x"01",	--6644
		x"4a",	--6645
		x"01",	--6646
		x"4a",	--6647
		x"00",	--6648
		x"4a",	--6649
		x"00",	--6650
		x"41",	--6651
		x"01",	--6652
		x"5f",	--6653
		x"5f",	--6654
		x"40",	--6655
		x"00",	--6656
		x"51",	--6657
		x"5f",	--6658
		x"51",	--6659
		x"01",	--6660
		x"49",	--6661
		x"01",	--6662
		x"49",	--6663
		x"49",	--6664
		x"00",	--6665
		x"48",	--6666
		x"49",	--6667
		x"46",	--6668
		x"47",	--6669
		x"12",	--6670
		x"bd",	--6671
		x"4e",	--6672
		x"4f",	--6673
		x"4e",	--6674
		x"4f",	--6675
		x"46",	--6676
		x"47",	--6677
		x"12",	--6678
		x"be",	--6679
		x"4e",	--6680
		x"4f",	--6681
		x"48",	--6682
		x"49",	--6683
		x"12",	--6684
		x"bd",	--6685
		x"41",	--6686
		x"01",	--6687
		x"4e",	--6688
		x"00",	--6689
		x"4f",	--6690
		x"00",	--6691
		x"41",	--6692
		x"01",	--6693
		x"4a",	--6694
		x"00",	--6695
		x"4b",	--6696
		x"00",	--6697
		x"53",	--6698
		x"63",	--6699
		x"82",	--6700
		x"01",	--6701
		x"3c",	--6702
		x"41",	--6703
		x"01",	--6704
		x"41",	--6705
		x"01",	--6706
		x"43",	--6707
		x"01",	--6708
		x"43",	--6709
		x"01",	--6710
		x"4c",	--6711
		x"4d",	--6712
		x"53",	--6713
		x"63",	--6714
		x"48",	--6715
		x"01",	--6716
		x"49",	--6717
		x"01",	--6718
		x"4c",	--6719
		x"4d",	--6720
		x"82",	--6721
		x"01",	--6722
		x"93",	--6723
		x"38",	--6724
		x"93",	--6725
		x"37",	--6726
		x"93",	--6727
		x"2f",	--6728
		x"41",	--6729
		x"01",	--6730
		x"41",	--6731
		x"01",	--6732
		x"43",	--6733
		x"01",	--6734
		x"43",	--6735
		x"01",	--6736
		x"4c",	--6737
		x"4d",	--6738
		x"53",	--6739
		x"63",	--6740
		x"49",	--6741
		x"01",	--6742
		x"4a",	--6743
		x"01",	--6744
		x"4c",	--6745
		x"4d",	--6746
		x"3c",	--6747
		x"41",	--6748
		x"01",	--6749
		x"5f",	--6750
		x"5f",	--6751
		x"40",	--6752
		x"00",	--6753
		x"51",	--6754
		x"5f",	--6755
		x"51",	--6756
		x"01",	--6757
		x"4a",	--6758
		x"01",	--6759
		x"4a",	--6760
		x"00",	--6761
		x"4a",	--6762
		x"00",	--6763
		x"41",	--6764
		x"01",	--6765
		x"5f",	--6766
		x"5f",	--6767
		x"40",	--6768
		x"00",	--6769
		x"51",	--6770
		x"5f",	--6771
		x"51",	--6772
		x"01",	--6773
		x"49",	--6774
		x"01",	--6775
		x"49",	--6776
		x"49",	--6777
		x"00",	--6778
		x"48",	--6779
		x"49",	--6780
		x"46",	--6781
		x"47",	--6782
		x"12",	--6783
		x"bd",	--6784
		x"4e",	--6785
		x"4f",	--6786
		x"4e",	--6787
		x"4f",	--6788
		x"46",	--6789
		x"47",	--6790
		x"12",	--6791
		x"be",	--6792
		x"4e",	--6793
		x"4f",	--6794
		x"48",	--6795
		x"49",	--6796
		x"12",	--6797
		x"bd",	--6798
		x"41",	--6799
		x"01",	--6800
		x"4e",	--6801
		x"00",	--6802
		x"4f",	--6803
		x"00",	--6804
		x"41",	--6805
		x"01",	--6806
		x"4a",	--6807
		x"00",	--6808
		x"4b",	--6809
		x"00",	--6810
		x"53",	--6811
		x"63",	--6812
		x"82",	--6813
		x"01",	--6814
		x"82",	--6815
		x"01",	--6816
		x"93",	--6817
		x"38",	--6818
		x"93",	--6819
		x"37",	--6820
		x"93",	--6821
		x"2f",	--6822
		x"41",	--6823
		x"01",	--6824
		x"41",	--6825
		x"01",	--6826
		x"43",	--6827
		x"43",	--6828
		x"43",	--6829
		x"3c",	--6830
		x"41",	--6831
		x"01",	--6832
		x"5f",	--6833
		x"5f",	--6834
		x"40",	--6835
		x"00",	--6836
		x"51",	--6837
		x"5d",	--6838
		x"55",	--6839
		x"4f",	--6840
		x"4f",	--6841
		x"00",	--6842
		x"4a",	--6843
		x"4b",	--6844
		x"12",	--6845
		x"bd",	--6846
		x"4e",	--6847
		x"4f",	--6848
		x"53",	--6849
		x"63",	--6850
		x"82",	--6851
		x"93",	--6852
		x"38",	--6853
		x"93",	--6854
		x"37",	--6855
		x"93",	--6856
		x"2f",	--6857
		x"93",	--6858
		x"01",	--6859
		x"20",	--6860
		x"93",	--6861
		x"01",	--6862
		x"20",	--6863
		x"41",	--6864
		x"01",	--6865
		x"41",	--6866
		x"00",	--6867
		x"00",	--6868
		x"41",	--6869
		x"00",	--6870
		x"00",	--6871
		x"41",	--6872
		x"00",	--6873
		x"00",	--6874
		x"41",	--6875
		x"00",	--6876
		x"00",	--6877
		x"4a",	--6878
		x"00",	--6879
		x"4b",	--6880
		x"00",	--6881
		x"3c",	--6882
		x"41",	--6883
		x"00",	--6884
		x"41",	--6885
		x"00",	--6886
		x"e0",	--6887
		x"80",	--6888
		x"41",	--6889
		x"01",	--6890
		x"4d",	--6891
		x"00",	--6892
		x"4e",	--6893
		x"00",	--6894
		x"41",	--6895
		x"00",	--6896
		x"41",	--6897
		x"00",	--6898
		x"e0",	--6899
		x"80",	--6900
		x"4d",	--6901
		x"00",	--6902
		x"4e",	--6903
		x"00",	--6904
		x"4a",	--6905
		x"4b",	--6906
		x"e0",	--6907
		x"80",	--6908
		x"4d",	--6909
		x"00",	--6910
		x"4e",	--6911
		x"00",	--6912
		x"41",	--6913
		x"01",	--6914
		x"f0",	--6915
		x"00",	--6916
		x"50",	--6917
		x"01",	--6918
		x"41",	--6919
		x"41",	--6920
		x"41",	--6921
		x"41",	--6922
		x"41",	--6923
		x"41",	--6924
		x"41",	--6925
		x"41",	--6926
		x"41",	--6927
		x"12",	--6928
		x"12",	--6929
		x"82",	--6930
		x"4e",	--6931
		x"4f",	--6932
		x"f3",	--6933
		x"f0",	--6934
		x"7f",	--6935
		x"90",	--6936
		x"3f",	--6937
		x"38",	--6938
		x"90",	--6939
		x"3f",	--6940
		x"34",	--6941
		x"90",	--6942
		x"0f",	--6943
		x"2c",	--6944
		x"43",	--6945
		x"43",	--6946
		x"3c",	--6947
		x"90",	--6948
		x"7f",	--6949
		x"38",	--6950
		x"4e",	--6951
		x"4f",	--6952
		x"12",	--6953
		x"be",	--6954
		x"3c",	--6955
		x"41",	--6956
		x"12",	--6957
		x"a3",	--6958
		x"4e",	--6959
		x"4f",	--6960
		x"f0",	--6961
		x"00",	--6962
		x"f3",	--6963
		x"41",	--6964
		x"00",	--6965
		x"41",	--6966
		x"00",	--6967
		x"41",	--6968
		x"41",	--6969
		x"00",	--6970
		x"93",	--6971
		x"20",	--6972
		x"93",	--6973
		x"24",	--6974
		x"93",	--6975
		x"20",	--6976
		x"93",	--6977
		x"24",	--6978
		x"41",	--6979
		x"41",	--6980
		x"00",	--6981
		x"93",	--6982
		x"20",	--6983
		x"93",	--6984
		x"20",	--6985
		x"12",	--6986
		x"a1",	--6987
		x"3c",	--6988
		x"12",	--6989
		x"12",	--6990
		x"b6",	--6991
		x"53",	--6992
		x"3c",	--6993
		x"12",	--6994
		x"a1",	--6995
		x"e0",	--6996
		x"80",	--6997
		x"3c",	--6998
		x"12",	--6999
		x"12",	--7000
		x"b6",	--7001
		x"53",	--7002
		x"52",	--7003
		x"41",	--7004
		x"41",	--7005
		x"41",	--7006
		x"12",	--7007
		x"b6",	--7008
		x"41",	--7009
		x"12",	--7010
		x"12",	--7011
		x"12",	--7012
		x"12",	--7013
		x"12",	--7014
		x"12",	--7015
		x"12",	--7016
		x"12",	--7017
		x"82",	--7018
		x"4e",	--7019
		x"4f",	--7020
		x"4c",	--7021
		x"00",	--7022
		x"4d",	--7023
		x"00",	--7024
		x"4e",	--7025
		x"4f",	--7026
		x"f3",	--7027
		x"f0",	--7028
		x"7f",	--7029
		x"90",	--7030
		x"32",	--7031
		x"34",	--7032
		x"12",	--7033
		x"c4",	--7034
		x"93",	--7035
		x"24",	--7036
		x"48",	--7037
		x"49",	--7038
		x"48",	--7039
		x"49",	--7040
		x"12",	--7041
		x"be",	--7042
		x"4e",	--7043
		x"4f",	--7044
		x"48",	--7045
		x"49",	--7046
		x"12",	--7047
		x"be",	--7048
		x"4e",	--7049
		x"4f",	--7050
		x"40",	--7051
		x"c9",	--7052
		x"40",	--7053
		x"2f",	--7054
		x"4a",	--7055
		x"4b",	--7056
		x"12",	--7057
		x"be",	--7058
		x"40",	--7059
		x"2f",	--7060
		x"40",	--7061
		x"32",	--7062
		x"12",	--7063
		x"be",	--7064
		x"4e",	--7065
		x"4f",	--7066
		x"4a",	--7067
		x"4b",	--7068
		x"12",	--7069
		x"be",	--7070
		x"40",	--7071
		x"ef",	--7072
		x"40",	--7073
		x"36",	--7074
		x"12",	--7075
		x"bd",	--7076
		x"4e",	--7077
		x"4f",	--7078
		x"4a",	--7079
		x"4b",	--7080
		x"12",	--7081
		x"be",	--7082
		x"40",	--7083
		x"0d",	--7084
		x"40",	--7085
		x"39",	--7086
		x"12",	--7087
		x"be",	--7088
		x"4e",	--7089
		x"4f",	--7090
		x"4a",	--7091
		x"4b",	--7092
		x"12",	--7093
		x"be",	--7094
		x"40",	--7095
		x"88",	--7096
		x"40",	--7097
		x"3c",	--7098
		x"12",	--7099
		x"bd",	--7100
		x"4e",	--7101
		x"4f",	--7102
		x"93",	--7103
		x"00",	--7104
		x"20",	--7105
		x"4e",	--7106
		x"4f",	--7107
		x"4a",	--7108
		x"4b",	--7109
		x"12",	--7110
		x"be",	--7111
		x"40",	--7112
		x"aa",	--7113
		x"40",	--7114
		x"3e",	--7115
		x"12",	--7116
		x"be",	--7117
		x"4e",	--7118
		x"4f",	--7119
		x"46",	--7120
		x"47",	--7121
		x"12",	--7122
		x"be",	--7123
		x"4e",	--7124
		x"4f",	--7125
		x"48",	--7126
		x"49",	--7127
		x"12",	--7128
		x"bd",	--7129
		x"3c",	--7130
		x"43",	--7131
		x"40",	--7132
		x"3f",	--7133
		x"41",	--7134
		x"41",	--7135
		x"00",	--7136
		x"12",	--7137
		x"be",	--7138
		x"4e",	--7139
		x"00",	--7140
		x"4f",	--7141
		x"00",	--7142
		x"44",	--7143
		x"45",	--7144
		x"46",	--7145
		x"47",	--7146
		x"12",	--7147
		x"be",	--7148
		x"4e",	--7149
		x"4f",	--7150
		x"41",	--7151
		x"00",	--7152
		x"41",	--7153
		x"00",	--7154
		x"12",	--7155
		x"be",	--7156
		x"4e",	--7157
		x"4f",	--7158
		x"4a",	--7159
		x"4b",	--7160
		x"12",	--7161
		x"be",	--7162
		x"41",	--7163
		x"41",	--7164
		x"00",	--7165
		x"12",	--7166
		x"be",	--7167
		x"4e",	--7168
		x"4f",	--7169
		x"40",	--7170
		x"aa",	--7171
		x"40",	--7172
		x"3e",	--7173
		x"46",	--7174
		x"47",	--7175
		x"12",	--7176
		x"be",	--7177
		x"4e",	--7178
		x"4f",	--7179
		x"4a",	--7180
		x"4b",	--7181
		x"12",	--7182
		x"bd",	--7183
		x"4e",	--7184
		x"4f",	--7185
		x"48",	--7186
		x"49",	--7187
		x"12",	--7188
		x"be",	--7189
		x"4e",	--7190
		x"4f",	--7191
		x"48",	--7192
		x"49",	--7193
		x"52",	--7194
		x"41",	--7195
		x"41",	--7196
		x"41",	--7197
		x"41",	--7198
		x"41",	--7199
		x"41",	--7200
		x"41",	--7201
		x"41",	--7202
		x"41",	--7203
		x"12",	--7204
		x"12",	--7205
		x"12",	--7206
		x"12",	--7207
		x"12",	--7208
		x"4d",	--7209
		x"4e",	--7210
		x"4f",	--7211
		x"48",	--7212
		x"49",	--7213
		x"f3",	--7214
		x"f0",	--7215
		x"7f",	--7216
		x"93",	--7217
		x"20",	--7218
		x"93",	--7219
		x"24",	--7220
		x"90",	--7221
		x"7f",	--7222
		x"28",	--7223
		x"4e",	--7224
		x"4f",	--7225
		x"12",	--7226
		x"bd",	--7227
		x"3c",	--7228
		x"90",	--7229
		x"00",	--7230
		x"28",	--7231
		x"4d",	--7232
		x"43",	--7233
		x"40",	--7234
		x"00",	--7235
		x"c3",	--7236
		x"10",	--7237
		x"10",	--7238
		x"53",	--7239
		x"23",	--7240
		x"3c",	--7241
		x"43",	--7242
		x"40",	--7243
		x"4c",	--7244
		x"12",	--7245
		x"be",	--7246
		x"4e",	--7247
		x"4f",	--7248
		x"48",	--7249
		x"49",	--7250
		x"f3",	--7251
		x"f0",	--7252
		x"7f",	--7253
		x"4b",	--7254
		x"4b",	--7255
		x"10",	--7256
		x"11",	--7257
		x"10",	--7258
		x"11",	--7259
		x"40",	--7260
		x"00",	--7261
		x"11",	--7262
		x"10",	--7263
		x"53",	--7264
		x"23",	--7265
		x"50",	--7266
		x"ff",	--7267
		x"63",	--7268
		x"47",	--7269
		x"47",	--7270
		x"10",	--7271
		x"11",	--7272
		x"10",	--7273
		x"11",	--7274
		x"4e",	--7275
		x"5a",	--7276
		x"6b",	--7277
		x"93",	--7278
		x"38",	--7279
		x"20",	--7280
		x"90",	--7281
		x"00",	--7282
		x"28",	--7283
		x"40",	--7284
		x"f2",	--7285
		x"40",	--7286
		x"71",	--7287
		x"93",	--7288
		x"34",	--7289
		x"40",	--7290
		x"f2",	--7291
		x"40",	--7292
		x"f1",	--7293
		x"40",	--7294
		x"f2",	--7295
		x"40",	--7296
		x"71",	--7297
		x"4a",	--7298
		x"4b",	--7299
		x"3c",	--7300
		x"93",	--7301
		x"38",	--7302
		x"20",	--7303
		x"93",	--7304
		x"28",	--7305
		x"43",	--7306
		x"43",	--7307
		x"4c",	--7308
		x"40",	--7309
		x"00",	--7310
		x"5a",	--7311
		x"6b",	--7312
		x"53",	--7313
		x"23",	--7314
		x"f3",	--7315
		x"f0",	--7316
		x"80",	--7317
		x"da",	--7318
		x"db",	--7319
		x"48",	--7320
		x"49",	--7321
		x"3c",	--7322
		x"93",	--7323
		x"38",	--7324
		x"93",	--7325
		x"34",	--7326
		x"90",	--7327
		x"ff",	--7328
		x"2c",	--7329
		x"4f",	--7330
		x"f0",	--7331
		x"80",	--7332
		x"90",	--7333
		x"75",	--7334
		x"38",	--7335
		x"40",	--7336
		x"f2",	--7337
		x"40",	--7338
		x"71",	--7339
		x"93",	--7340
		x"24",	--7341
		x"40",	--7342
		x"f2",	--7343
		x"40",	--7344
		x"f1",	--7345
		x"40",	--7346
		x"f2",	--7347
		x"40",	--7348
		x"71",	--7349
		x"3c",	--7350
		x"40",	--7351
		x"42",	--7352
		x"40",	--7353
		x"0d",	--7354
		x"93",	--7355
		x"24",	--7356
		x"40",	--7357
		x"42",	--7358
		x"40",	--7359
		x"8d",	--7360
		x"40",	--7361
		x"42",	--7362
		x"40",	--7363
		x"0d",	--7364
		x"3c",	--7365
		x"43",	--7366
		x"43",	--7367
		x"4c",	--7368
		x"50",	--7369
		x"00",	--7370
		x"40",	--7371
		x"00",	--7372
		x"5a",	--7373
		x"6b",	--7374
		x"53",	--7375
		x"23",	--7376
		x"48",	--7377
		x"49",	--7378
		x"f3",	--7379
		x"f0",	--7380
		x"80",	--7381
		x"da",	--7382
		x"db",	--7383
		x"43",	--7384
		x"40",	--7385
		x"33",	--7386
		x"12",	--7387
		x"be",	--7388
		x"41",	--7389
		x"41",	--7390
		x"41",	--7391
		x"41",	--7392
		x"41",	--7393
		x"41",	--7394
		x"12",	--7395
		x"b8",	--7396
		x"41",	--7397
		x"12",	--7398
		x"12",	--7399
		x"12",	--7400
		x"12",	--7401
		x"12",	--7402
		x"12",	--7403
		x"12",	--7404
		x"12",	--7405
		x"83",	--7406
		x"4e",	--7407
		x"4f",	--7408
		x"4e",	--7409
		x"4f",	--7410
		x"f3",	--7411
		x"f0",	--7412
		x"7f",	--7413
		x"49",	--7414
		x"43",	--7415
		x"40",	--7416
		x"00",	--7417
		x"c3",	--7418
		x"10",	--7419
		x"10",	--7420
		x"53",	--7421
		x"23",	--7422
		x"50",	--7423
		x"ff",	--7424
		x"63",	--7425
		x"93",	--7426
		x"38",	--7427
		x"93",	--7428
		x"34",	--7429
		x"90",	--7430
		x"00",	--7431
		x"2c",	--7432
		x"46",	--7433
		x"47",	--7434
		x"93",	--7435
		x"38",	--7436
		x"4c",	--7437
		x"00",	--7438
		x"43",	--7439
		x"40",	--7440
		x"00",	--7441
		x"41",	--7442
		x"f0",	--7443
		x"00",	--7444
		x"3c",	--7445
		x"40",	--7446
		x"f2",	--7447
		x"40",	--7448
		x"71",	--7449
		x"12",	--7450
		x"bd",	--7451
		x"43",	--7452
		x"43",	--7453
		x"12",	--7454
		x"c2",	--7455
		x"93",	--7456
		x"24",	--7457
		x"38",	--7458
		x"93",	--7459
		x"38",	--7460
		x"43",	--7461
		x"43",	--7462
		x"3c",	--7463
		x"93",	--7464
		x"20",	--7465
		x"93",	--7466
		x"24",	--7467
		x"43",	--7468
		x"40",	--7469
		x"bf",	--7470
		x"3c",	--7471
		x"11",	--7472
		x"10",	--7473
		x"53",	--7474
		x"93",	--7475
		x"23",	--7476
		x"48",	--7477
		x"49",	--7478
		x"f6",	--7479
		x"f7",	--7480
		x"93",	--7481
		x"20",	--7482
		x"93",	--7483
		x"24",	--7484
		x"40",	--7485
		x"f2",	--7486
		x"40",	--7487
		x"71",	--7488
		x"12",	--7489
		x"bd",	--7490
		x"43",	--7491
		x"43",	--7492
		x"12",	--7493
		x"c2",	--7494
		x"93",	--7495
		x"24",	--7496
		x"38",	--7497
		x"93",	--7498
		x"34",	--7499
		x"43",	--7500
		x"40",	--7501
		x"00",	--7502
		x"41",	--7503
		x"f0",	--7504
		x"00",	--7505
		x"93",	--7506
		x"24",	--7507
		x"11",	--7508
		x"10",	--7509
		x"53",	--7510
		x"3f",	--7511
		x"56",	--7512
		x"67",	--7513
		x"c8",	--7514
		x"c9",	--7515
		x"3c",	--7516
		x"90",	--7517
		x"7f",	--7518
		x"28",	--7519
		x"4e",	--7520
		x"4f",	--7521
		x"12",	--7522
		x"bd",	--7523
		x"3c",	--7524
		x"4a",	--7525
		x"4b",	--7526
		x"53",	--7527
		x"41",	--7528
		x"41",	--7529
		x"41",	--7530
		x"41",	--7531
		x"41",	--7532
		x"41",	--7533
		x"41",	--7534
		x"41",	--7535
		x"41",	--7536
		x"12",	--7537
		x"b9",	--7538
		x"41",	--7539
		x"12",	--7540
		x"12",	--7541
		x"4e",	--7542
		x"4f",	--7543
		x"43",	--7544
		x"40",	--7545
		x"4f",	--7546
		x"12",	--7547
		x"c2",	--7548
		x"93",	--7549
		x"34",	--7550
		x"4a",	--7551
		x"4b",	--7552
		x"12",	--7553
		x"c4",	--7554
		x"41",	--7555
		x"41",	--7556
		x"41",	--7557
		x"43",	--7558
		x"40",	--7559
		x"4f",	--7560
		x"4a",	--7561
		x"4b",	--7562
		x"12",	--7563
		x"be",	--7564
		x"12",	--7565
		x"c4",	--7566
		x"53",	--7567
		x"60",	--7568
		x"80",	--7569
		x"41",	--7570
		x"41",	--7571
		x"41",	--7572
		x"12",	--7573
		x"12",	--7574
		x"12",	--7575
		x"12",	--7576
		x"12",	--7577
		x"12",	--7578
		x"12",	--7579
		x"12",	--7580
		x"50",	--7581
		x"ff",	--7582
		x"4d",	--7583
		x"4f",	--7584
		x"93",	--7585
		x"28",	--7586
		x"4e",	--7587
		x"93",	--7588
		x"28",	--7589
		x"92",	--7590
		x"20",	--7591
		x"40",	--7592
		x"bd",	--7593
		x"92",	--7594
		x"24",	--7595
		x"93",	--7596
		x"24",	--7597
		x"93",	--7598
		x"24",	--7599
		x"4f",	--7600
		x"00",	--7601
		x"00",	--7602
		x"4e",	--7603
		x"00",	--7604
		x"4f",	--7605
		x"00",	--7606
		x"4f",	--7607
		x"00",	--7608
		x"4e",	--7609
		x"00",	--7610
		x"4e",	--7611
		x"00",	--7612
		x"41",	--7613
		x"8b",	--7614
		x"4c",	--7615
		x"93",	--7616
		x"38",	--7617
		x"90",	--7618
		x"00",	--7619
		x"34",	--7620
		x"93",	--7621
		x"38",	--7622
		x"46",	--7623
		x"00",	--7624
		x"47",	--7625
		x"00",	--7626
		x"49",	--7627
		x"f0",	--7628
		x"00",	--7629
		x"24",	--7630
		x"46",	--7631
		x"47",	--7632
		x"c3",	--7633
		x"10",	--7634
		x"10",	--7635
		x"53",	--7636
		x"23",	--7637
		x"4a",	--7638
		x"00",	--7639
		x"4b",	--7640
		x"00",	--7641
		x"43",	--7642
		x"43",	--7643
		x"f0",	--7644
		x"00",	--7645
		x"24",	--7646
		x"5c",	--7647
		x"6d",	--7648
		x"53",	--7649
		x"23",	--7650
		x"53",	--7651
		x"63",	--7652
		x"f6",	--7653
		x"f7",	--7654
		x"43",	--7655
		x"43",	--7656
		x"93",	--7657
		x"20",	--7658
		x"93",	--7659
		x"24",	--7660
		x"41",	--7661
		x"00",	--7662
		x"41",	--7663
		x"00",	--7664
		x"da",	--7665
		x"db",	--7666
		x"4f",	--7667
		x"00",	--7668
		x"9e",	--7669
		x"00",	--7670
		x"20",	--7671
		x"4f",	--7672
		x"00",	--7673
		x"41",	--7674
		x"00",	--7675
		x"46",	--7676
		x"47",	--7677
		x"54",	--7678
		x"65",	--7679
		x"4e",	--7680
		x"00",	--7681
		x"4f",	--7682
		x"00",	--7683
		x"40",	--7684
		x"00",	--7685
		x"00",	--7686
		x"93",	--7687
		x"38",	--7688
		x"48",	--7689
		x"50",	--7690
		x"00",	--7691
		x"41",	--7692
		x"41",	--7693
		x"41",	--7694
		x"41",	--7695
		x"41",	--7696
		x"41",	--7697
		x"41",	--7698
		x"41",	--7699
		x"41",	--7700
		x"91",	--7701
		x"38",	--7702
		x"4b",	--7703
		x"00",	--7704
		x"43",	--7705
		x"43",	--7706
		x"4f",	--7707
		x"00",	--7708
		x"9e",	--7709
		x"00",	--7710
		x"27",	--7711
		x"93",	--7712
		x"24",	--7713
		x"46",	--7714
		x"47",	--7715
		x"84",	--7716
		x"75",	--7717
		x"93",	--7718
		x"38",	--7719
		x"43",	--7720
		x"00",	--7721
		x"41",	--7722
		x"00",	--7723
		x"4e",	--7724
		x"00",	--7725
		x"4f",	--7726
		x"00",	--7727
		x"4e",	--7728
		x"4f",	--7729
		x"53",	--7730
		x"63",	--7731
		x"90",	--7732
		x"3f",	--7733
		x"28",	--7734
		x"90",	--7735
		x"40",	--7736
		x"2c",	--7737
		x"93",	--7738
		x"2c",	--7739
		x"48",	--7740
		x"00",	--7741
		x"53",	--7742
		x"5e",	--7743
		x"6f",	--7744
		x"4b",	--7745
		x"53",	--7746
		x"4e",	--7747
		x"4f",	--7748
		x"53",	--7749
		x"63",	--7750
		x"90",	--7751
		x"3f",	--7752
		x"2b",	--7753
		x"24",	--7754
		x"4e",	--7755
		x"00",	--7756
		x"4f",	--7757
		x"00",	--7758
		x"4a",	--7759
		x"00",	--7760
		x"40",	--7761
		x"00",	--7762
		x"00",	--7763
		x"93",	--7764
		x"37",	--7765
		x"4e",	--7766
		x"4f",	--7767
		x"f3",	--7768
		x"f3",	--7769
		x"c3",	--7770
		x"10",	--7771
		x"10",	--7772
		x"4c",	--7773
		x"4d",	--7774
		x"de",	--7775
		x"df",	--7776
		x"4a",	--7777
		x"00",	--7778
		x"4b",	--7779
		x"00",	--7780
		x"53",	--7781
		x"00",	--7782
		x"48",	--7783
		x"3f",	--7784
		x"93",	--7785
		x"23",	--7786
		x"4f",	--7787
		x"00",	--7788
		x"4f",	--7789
		x"00",	--7790
		x"00",	--7791
		x"4f",	--7792
		x"00",	--7793
		x"00",	--7794
		x"4f",	--7795
		x"00",	--7796
		x"00",	--7797
		x"4e",	--7798
		x"00",	--7799
		x"ff",	--7800
		x"00",	--7801
		x"4e",	--7802
		x"00",	--7803
		x"4d",	--7804
		x"3f",	--7805
		x"43",	--7806
		x"43",	--7807
		x"3f",	--7808
		x"e3",	--7809
		x"53",	--7810
		x"90",	--7811
		x"00",	--7812
		x"37",	--7813
		x"3f",	--7814
		x"93",	--7815
		x"2b",	--7816
		x"3f",	--7817
		x"44",	--7818
		x"45",	--7819
		x"86",	--7820
		x"77",	--7821
		x"3f",	--7822
		x"4e",	--7823
		x"3f",	--7824
		x"43",	--7825
		x"00",	--7826
		x"41",	--7827
		x"00",	--7828
		x"e3",	--7829
		x"e3",	--7830
		x"53",	--7831
		x"63",	--7832
		x"4e",	--7833
		x"00",	--7834
		x"4f",	--7835
		x"00",	--7836
		x"3f",	--7837
		x"93",	--7838
		x"27",	--7839
		x"59",	--7840
		x"00",	--7841
		x"44",	--7842
		x"00",	--7843
		x"45",	--7844
		x"00",	--7845
		x"49",	--7846
		x"f0",	--7847
		x"00",	--7848
		x"24",	--7849
		x"4d",	--7850
		x"44",	--7851
		x"45",	--7852
		x"c3",	--7853
		x"10",	--7854
		x"10",	--7855
		x"53",	--7856
		x"23",	--7857
		x"4c",	--7858
		x"00",	--7859
		x"4d",	--7860
		x"00",	--7861
		x"43",	--7862
		x"43",	--7863
		x"f0",	--7864
		x"00",	--7865
		x"24",	--7866
		x"5c",	--7867
		x"6d",	--7868
		x"53",	--7869
		x"23",	--7870
		x"53",	--7871
		x"63",	--7872
		x"f4",	--7873
		x"f5",	--7874
		x"43",	--7875
		x"43",	--7876
		x"93",	--7877
		x"20",	--7878
		x"93",	--7879
		x"20",	--7880
		x"43",	--7881
		x"43",	--7882
		x"41",	--7883
		x"00",	--7884
		x"41",	--7885
		x"00",	--7886
		x"da",	--7887
		x"db",	--7888
		x"3f",	--7889
		x"43",	--7890
		x"43",	--7891
		x"3f",	--7892
		x"92",	--7893
		x"23",	--7894
		x"9e",	--7895
		x"00",	--7896
		x"00",	--7897
		x"27",	--7898
		x"40",	--7899
		x"dc",	--7900
		x"3f",	--7901
		x"50",	--7902
		x"ff",	--7903
		x"4e",	--7904
		x"00",	--7905
		x"4f",	--7906
		x"00",	--7907
		x"4c",	--7908
		x"00",	--7909
		x"4d",	--7910
		x"00",	--7911
		x"41",	--7912
		x"50",	--7913
		x"00",	--7914
		x"41",	--7915
		x"52",	--7916
		x"12",	--7917
		x"c7",	--7918
		x"41",	--7919
		x"50",	--7920
		x"00",	--7921
		x"41",	--7922
		x"12",	--7923
		x"c7",	--7924
		x"41",	--7925
		x"52",	--7926
		x"41",	--7927
		x"50",	--7928
		x"00",	--7929
		x"41",	--7930
		x"50",	--7931
		x"00",	--7932
		x"12",	--7933
		x"bb",	--7934
		x"12",	--7935
		x"c5",	--7936
		x"50",	--7937
		x"00",	--7938
		x"41",	--7939
		x"50",	--7940
		x"ff",	--7941
		x"4e",	--7942
		x"00",	--7943
		x"4f",	--7944
		x"00",	--7945
		x"4c",	--7946
		x"00",	--7947
		x"4d",	--7948
		x"00",	--7949
		x"41",	--7950
		x"50",	--7951
		x"00",	--7952
		x"41",	--7953
		x"52",	--7954
		x"12",	--7955
		x"c7",	--7956
		x"41",	--7957
		x"50",	--7958
		x"00",	--7959
		x"41",	--7960
		x"12",	--7961
		x"c7",	--7962
		x"e3",	--7963
		x"00",	--7964
		x"41",	--7965
		x"52",	--7966
		x"41",	--7967
		x"50",	--7968
		x"00",	--7969
		x"41",	--7970
		x"50",	--7971
		x"00",	--7972
		x"12",	--7973
		x"bb",	--7974
		x"12",	--7975
		x"c5",	--7976
		x"50",	--7977
		x"00",	--7978
		x"41",	--7979
		x"12",	--7980
		x"12",	--7981
		x"12",	--7982
		x"12",	--7983
		x"12",	--7984
		x"12",	--7985
		x"12",	--7986
		x"12",	--7987
		x"50",	--7988
		x"ff",	--7989
		x"4e",	--7990
		x"00",	--7991
		x"4f",	--7992
		x"00",	--7993
		x"4c",	--7994
		x"00",	--7995
		x"4d",	--7996
		x"00",	--7997
		x"41",	--7998
		x"50",	--7999
		x"00",	--8000
		x"41",	--8001
		x"52",	--8002
		x"12",	--8003
		x"c7",	--8004
		x"41",	--8005
		x"50",	--8006
		x"00",	--8007
		x"41",	--8008
		x"12",	--8009
		x"c7",	--8010
		x"41",	--8011
		x"00",	--8012
		x"93",	--8013
		x"28",	--8014
		x"41",	--8015
		x"00",	--8016
		x"93",	--8017
		x"28",	--8018
		x"92",	--8019
		x"24",	--8020
		x"92",	--8021
		x"24",	--8022
		x"93",	--8023
		x"24",	--8024
		x"93",	--8025
		x"24",	--8026
		x"41",	--8027
		x"00",	--8028
		x"41",	--8029
		x"00",	--8030
		x"41",	--8031
		x"00",	--8032
		x"41",	--8033
		x"00",	--8034
		x"40",	--8035
		x"00",	--8036
		x"43",	--8037
		x"43",	--8038
		x"43",	--8039
		x"43",	--8040
		x"43",	--8041
		x"00",	--8042
		x"43",	--8043
		x"00",	--8044
		x"43",	--8045
		x"43",	--8046
		x"4c",	--8047
		x"00",	--8048
		x"3c",	--8049
		x"58",	--8050
		x"69",	--8051
		x"c3",	--8052
		x"10",	--8053
		x"10",	--8054
		x"53",	--8055
		x"00",	--8056
		x"24",	--8057
		x"b3",	--8058
		x"24",	--8059
		x"58",	--8060
		x"69",	--8061
		x"56",	--8062
		x"67",	--8063
		x"43",	--8064
		x"43",	--8065
		x"99",	--8066
		x"28",	--8067
		x"24",	--8068
		x"43",	--8069
		x"43",	--8070
		x"5c",	--8071
		x"6d",	--8072
		x"56",	--8073
		x"67",	--8074
		x"93",	--8075
		x"37",	--8076
		x"d3",	--8077
		x"d3",	--8078
		x"3f",	--8079
		x"98",	--8080
		x"2b",	--8081
		x"3f",	--8082
		x"4a",	--8083
		x"00",	--8084
		x"4b",	--8085
		x"00",	--8086
		x"4f",	--8087
		x"41",	--8088
		x"00",	--8089
		x"51",	--8090
		x"00",	--8091
		x"4a",	--8092
		x"53",	--8093
		x"46",	--8094
		x"00",	--8095
		x"43",	--8096
		x"91",	--8097
		x"00",	--8098
		x"00",	--8099
		x"24",	--8100
		x"4d",	--8101
		x"00",	--8102
		x"93",	--8103
		x"38",	--8104
		x"90",	--8105
		x"40",	--8106
		x"2c",	--8107
		x"41",	--8108
		x"00",	--8109
		x"53",	--8110
		x"41",	--8111
		x"00",	--8112
		x"41",	--8113
		x"00",	--8114
		x"4d",	--8115
		x"5e",	--8116
		x"6f",	--8117
		x"93",	--8118
		x"38",	--8119
		x"5a",	--8120
		x"6b",	--8121
		x"53",	--8122
		x"90",	--8123
		x"40",	--8124
		x"2b",	--8125
		x"4a",	--8126
		x"00",	--8127
		x"4b",	--8128
		x"00",	--8129
		x"4c",	--8130
		x"00",	--8131
		x"4e",	--8132
		x"4f",	--8133
		x"f0",	--8134
		x"00",	--8135
		x"f3",	--8136
		x"90",	--8137
		x"00",	--8138
		x"24",	--8139
		x"4e",	--8140
		x"00",	--8141
		x"4f",	--8142
		x"00",	--8143
		x"40",	--8144
		x"00",	--8145
		x"00",	--8146
		x"41",	--8147
		x"52",	--8148
		x"12",	--8149
		x"c5",	--8150
		x"50",	--8151
		x"00",	--8152
		x"41",	--8153
		x"41",	--8154
		x"41",	--8155
		x"41",	--8156
		x"41",	--8157
		x"41",	--8158
		x"41",	--8159
		x"41",	--8160
		x"41",	--8161
		x"d3",	--8162
		x"d3",	--8163
		x"3f",	--8164
		x"50",	--8165
		x"00",	--8166
		x"4a",	--8167
		x"b3",	--8168
		x"24",	--8169
		x"41",	--8170
		x"00",	--8171
		x"41",	--8172
		x"00",	--8173
		x"c3",	--8174
		x"10",	--8175
		x"10",	--8176
		x"4c",	--8177
		x"4d",	--8178
		x"d3",	--8179
		x"d0",	--8180
		x"80",	--8181
		x"46",	--8182
		x"00",	--8183
		x"47",	--8184
		x"00",	--8185
		x"c3",	--8186
		x"10",	--8187
		x"10",	--8188
		x"53",	--8189
		x"93",	--8190
		x"3b",	--8191
		x"48",	--8192
		x"00",	--8193
		x"3f",	--8194
		x"93",	--8195
		x"24",	--8196
		x"43",	--8197
		x"91",	--8198
		x"00",	--8199
		x"00",	--8200
		x"24",	--8201
		x"4f",	--8202
		x"00",	--8203
		x"41",	--8204
		x"50",	--8205
		x"00",	--8206
		x"3f",	--8207
		x"93",	--8208
		x"23",	--8209
		x"4e",	--8210
		x"4f",	--8211
		x"f0",	--8212
		x"00",	--8213
		x"f3",	--8214
		x"93",	--8215
		x"23",	--8216
		x"93",	--8217
		x"23",	--8218
		x"93",	--8219
		x"00",	--8220
		x"20",	--8221
		x"93",	--8222
		x"00",	--8223
		x"27",	--8224
		x"50",	--8225
		x"00",	--8226
		x"63",	--8227
		x"f0",	--8228
		x"ff",	--8229
		x"f3",	--8230
		x"3f",	--8231
		x"43",	--8232
		x"3f",	--8233
		x"43",	--8234
		x"3f",	--8235
		x"43",	--8236
		x"91",	--8237
		x"00",	--8238
		x"00",	--8239
		x"24",	--8240
		x"4f",	--8241
		x"00",	--8242
		x"41",	--8243
		x"50",	--8244
		x"00",	--8245
		x"3f",	--8246
		x"43",	--8247
		x"3f",	--8248
		x"93",	--8249
		x"23",	--8250
		x"40",	--8251
		x"dc",	--8252
		x"3f",	--8253
		x"12",	--8254
		x"12",	--8255
		x"12",	--8256
		x"12",	--8257
		x"12",	--8258
		x"50",	--8259
		x"ff",	--8260
		x"4e",	--8261
		x"00",	--8262
		x"4f",	--8263
		x"00",	--8264
		x"4c",	--8265
		x"00",	--8266
		x"4d",	--8267
		x"00",	--8268
		x"41",	--8269
		x"50",	--8270
		x"00",	--8271
		x"41",	--8272
		x"52",	--8273
		x"12",	--8274
		x"c7",	--8275
		x"41",	--8276
		x"52",	--8277
		x"41",	--8278
		x"12",	--8279
		x"c7",	--8280
		x"41",	--8281
		x"00",	--8282
		x"93",	--8283
		x"28",	--8284
		x"41",	--8285
		x"00",	--8286
		x"93",	--8287
		x"28",	--8288
		x"e1",	--8289
		x"00",	--8290
		x"00",	--8291
		x"92",	--8292
		x"24",	--8293
		x"93",	--8294
		x"24",	--8295
		x"92",	--8296
		x"24",	--8297
		x"93",	--8298
		x"24",	--8299
		x"41",	--8300
		x"00",	--8301
		x"81",	--8302
		x"00",	--8303
		x"4d",	--8304
		x"00",	--8305
		x"41",	--8306
		x"00",	--8307
		x"41",	--8308
		x"00",	--8309
		x"41",	--8310
		x"00",	--8311
		x"41",	--8312
		x"00",	--8313
		x"99",	--8314
		x"2c",	--8315
		x"5e",	--8316
		x"6f",	--8317
		x"53",	--8318
		x"4d",	--8319
		x"00",	--8320
		x"40",	--8321
		x"00",	--8322
		x"43",	--8323
		x"40",	--8324
		x"40",	--8325
		x"43",	--8326
		x"43",	--8327
		x"3c",	--8328
		x"dc",	--8329
		x"dd",	--8330
		x"88",	--8331
		x"79",	--8332
		x"c3",	--8333
		x"10",	--8334
		x"10",	--8335
		x"5e",	--8336
		x"6f",	--8337
		x"53",	--8338
		x"24",	--8339
		x"99",	--8340
		x"2b",	--8341
		x"23",	--8342
		x"98",	--8343
		x"2b",	--8344
		x"3f",	--8345
		x"9f",	--8346
		x"2b",	--8347
		x"98",	--8348
		x"2f",	--8349
		x"3f",	--8350
		x"4a",	--8351
		x"4b",	--8352
		x"f0",	--8353
		x"00",	--8354
		x"f3",	--8355
		x"90",	--8356
		x"00",	--8357
		x"24",	--8358
		x"4a",	--8359
		x"00",	--8360
		x"4b",	--8361
		x"00",	--8362
		x"41",	--8363
		x"50",	--8364
		x"00",	--8365
		x"12",	--8366
		x"c5",	--8367
		x"50",	--8368
		x"00",	--8369
		x"41",	--8370
		x"41",	--8371
		x"41",	--8372
		x"41",	--8373
		x"41",	--8374
		x"41",	--8375
		x"42",	--8376
		x"00",	--8377
		x"41",	--8378
		x"50",	--8379
		x"00",	--8380
		x"3f",	--8381
		x"9e",	--8382
		x"23",	--8383
		x"40",	--8384
		x"dc",	--8385
		x"3f",	--8386
		x"93",	--8387
		x"23",	--8388
		x"4a",	--8389
		x"4b",	--8390
		x"f0",	--8391
		x"00",	--8392
		x"f3",	--8393
		x"93",	--8394
		x"23",	--8395
		x"93",	--8396
		x"23",	--8397
		x"93",	--8398
		x"20",	--8399
		x"93",	--8400
		x"27",	--8401
		x"50",	--8402
		x"00",	--8403
		x"63",	--8404
		x"f0",	--8405
		x"ff",	--8406
		x"f3",	--8407
		x"3f",	--8408
		x"43",	--8409
		x"00",	--8410
		x"43",	--8411
		x"00",	--8412
		x"43",	--8413
		x"00",	--8414
		x"41",	--8415
		x"50",	--8416
		x"00",	--8417
		x"3f",	--8418
		x"41",	--8419
		x"52",	--8420
		x"3f",	--8421
		x"50",	--8422
		x"ff",	--8423
		x"4e",	--8424
		x"00",	--8425
		x"4f",	--8426
		x"00",	--8427
		x"4c",	--8428
		x"00",	--8429
		x"4d",	--8430
		x"00",	--8431
		x"41",	--8432
		x"50",	--8433
		x"00",	--8434
		x"41",	--8435
		x"52",	--8436
		x"12",	--8437
		x"c7",	--8438
		x"41",	--8439
		x"52",	--8440
		x"41",	--8441
		x"12",	--8442
		x"c7",	--8443
		x"93",	--8444
		x"00",	--8445
		x"28",	--8446
		x"93",	--8447
		x"00",	--8448
		x"28",	--8449
		x"41",	--8450
		x"52",	--8451
		x"41",	--8452
		x"50",	--8453
		x"00",	--8454
		x"12",	--8455
		x"c8",	--8456
		x"50",	--8457
		x"00",	--8458
		x"41",	--8459
		x"43",	--8460
		x"3f",	--8461
		x"50",	--8462
		x"ff",	--8463
		x"4e",	--8464
		x"00",	--8465
		x"4f",	--8466
		x"00",	--8467
		x"4c",	--8468
		x"00",	--8469
		x"4d",	--8470
		x"00",	--8471
		x"41",	--8472
		x"50",	--8473
		x"00",	--8474
		x"41",	--8475
		x"52",	--8476
		x"12",	--8477
		x"c7",	--8478
		x"41",	--8479
		x"52",	--8480
		x"41",	--8481
		x"12",	--8482
		x"c7",	--8483
		x"93",	--8484
		x"00",	--8485
		x"28",	--8486
		x"93",	--8487
		x"00",	--8488
		x"28",	--8489
		x"41",	--8490
		x"52",	--8491
		x"41",	--8492
		x"50",	--8493
		x"00",	--8494
		x"12",	--8495
		x"c8",	--8496
		x"50",	--8497
		x"00",	--8498
		x"41",	--8499
		x"43",	--8500
		x"3f",	--8501
		x"50",	--8502
		x"ff",	--8503
		x"4e",	--8504
		x"00",	--8505
		x"4f",	--8506
		x"00",	--8507
		x"4c",	--8508
		x"00",	--8509
		x"4d",	--8510
		x"00",	--8511
		x"41",	--8512
		x"50",	--8513
		x"00",	--8514
		x"41",	--8515
		x"52",	--8516
		x"12",	--8517
		x"c7",	--8518
		x"41",	--8519
		x"52",	--8520
		x"41",	--8521
		x"12",	--8522
		x"c7",	--8523
		x"93",	--8524
		x"00",	--8525
		x"28",	--8526
		x"93",	--8527
		x"00",	--8528
		x"28",	--8529
		x"41",	--8530
		x"52",	--8531
		x"41",	--8532
		x"50",	--8533
		x"00",	--8534
		x"12",	--8535
		x"c8",	--8536
		x"50",	--8537
		x"00",	--8538
		x"41",	--8539
		x"43",	--8540
		x"3f",	--8541
		x"50",	--8542
		x"ff",	--8543
		x"4e",	--8544
		x"00",	--8545
		x"4f",	--8546
		x"00",	--8547
		x"4c",	--8548
		x"00",	--8549
		x"4d",	--8550
		x"00",	--8551
		x"41",	--8552
		x"50",	--8553
		x"00",	--8554
		x"41",	--8555
		x"52",	--8556
		x"12",	--8557
		x"c7",	--8558
		x"41",	--8559
		x"52",	--8560
		x"41",	--8561
		x"12",	--8562
		x"c7",	--8563
		x"93",	--8564
		x"00",	--8565
		x"28",	--8566
		x"93",	--8567
		x"00",	--8568
		x"28",	--8569
		x"41",	--8570
		x"52",	--8571
		x"41",	--8572
		x"50",	--8573
		x"00",	--8574
		x"12",	--8575
		x"c8",	--8576
		x"50",	--8577
		x"00",	--8578
		x"41",	--8579
		x"43",	--8580
		x"3f",	--8581
		x"50",	--8582
		x"ff",	--8583
		x"4e",	--8584
		x"00",	--8585
		x"4f",	--8586
		x"00",	--8587
		x"4c",	--8588
		x"00",	--8589
		x"4d",	--8590
		x"00",	--8591
		x"41",	--8592
		x"50",	--8593
		x"00",	--8594
		x"41",	--8595
		x"52",	--8596
		x"12",	--8597
		x"c7",	--8598
		x"41",	--8599
		x"52",	--8600
		x"41",	--8601
		x"12",	--8602
		x"c7",	--8603
		x"93",	--8604
		x"00",	--8605
		x"28",	--8606
		x"93",	--8607
		x"00",	--8608
		x"28",	--8609
		x"41",	--8610
		x"52",	--8611
		x"41",	--8612
		x"50",	--8613
		x"00",	--8614
		x"12",	--8615
		x"c8",	--8616
		x"50",	--8617
		x"00",	--8618
		x"41",	--8619
		x"43",	--8620
		x"3f",	--8621
		x"12",	--8622
		x"12",	--8623
		x"82",	--8624
		x"40",	--8625
		x"00",	--8626
		x"00",	--8627
		x"4f",	--8628
		x"5d",	--8629
		x"43",	--8630
		x"6d",	--8631
		x"4d",	--8632
		x"4d",	--8633
		x"00",	--8634
		x"93",	--8635
		x"20",	--8636
		x"93",	--8637
		x"20",	--8638
		x"43",	--8639
		x"00",	--8640
		x"41",	--8641
		x"12",	--8642
		x"c5",	--8643
		x"52",	--8644
		x"41",	--8645
		x"41",	--8646
		x"41",	--8647
		x"40",	--8648
		x"00",	--8649
		x"00",	--8650
		x"93",	--8651
		x"20",	--8652
		x"4e",	--8653
		x"4f",	--8654
		x"4a",	--8655
		x"00",	--8656
		x"4b",	--8657
		x"00",	--8658
		x"4a",	--8659
		x"4b",	--8660
		x"12",	--8661
		x"c5",	--8662
		x"53",	--8663
		x"93",	--8664
		x"3b",	--8665
		x"4a",	--8666
		x"00",	--8667
		x"4b",	--8668
		x"00",	--8669
		x"4f",	--8670
		x"f0",	--8671
		x"00",	--8672
		x"20",	--8673
		x"40",	--8674
		x"00",	--8675
		x"8f",	--8676
		x"4e",	--8677
		x"00",	--8678
		x"3f",	--8679
		x"93",	--8680
		x"24",	--8681
		x"4e",	--8682
		x"4f",	--8683
		x"e3",	--8684
		x"e3",	--8685
		x"53",	--8686
		x"63",	--8687
		x"3f",	--8688
		x"51",	--8689
		x"00",	--8690
		x"00",	--8691
		x"61",	--8692
		x"00",	--8693
		x"00",	--8694
		x"53",	--8695
		x"23",	--8696
		x"3f",	--8697
		x"90",	--8698
		x"80",	--8699
		x"23",	--8700
		x"43",	--8701
		x"40",	--8702
		x"cf",	--8703
		x"3f",	--8704
		x"50",	--8705
		x"ff",	--8706
		x"4e",	--8707
		x"00",	--8708
		x"4f",	--8709
		x"00",	--8710
		x"41",	--8711
		x"52",	--8712
		x"41",	--8713
		x"12",	--8714
		x"c7",	--8715
		x"41",	--8716
		x"00",	--8717
		x"93",	--8718
		x"24",	--8719
		x"28",	--8720
		x"92",	--8721
		x"24",	--8722
		x"41",	--8723
		x"00",	--8724
		x"93",	--8725
		x"38",	--8726
		x"90",	--8727
		x"00",	--8728
		x"38",	--8729
		x"93",	--8730
		x"00",	--8731
		x"20",	--8732
		x"43",	--8733
		x"40",	--8734
		x"7f",	--8735
		x"50",	--8736
		x"00",	--8737
		x"41",	--8738
		x"41",	--8739
		x"00",	--8740
		x"41",	--8741
		x"00",	--8742
		x"40",	--8743
		x"00",	--8744
		x"8d",	--8745
		x"4c",	--8746
		x"f0",	--8747
		x"00",	--8748
		x"20",	--8749
		x"93",	--8750
		x"00",	--8751
		x"27",	--8752
		x"e3",	--8753
		x"e3",	--8754
		x"53",	--8755
		x"63",	--8756
		x"50",	--8757
		x"00",	--8758
		x"41",	--8759
		x"43",	--8760
		x"43",	--8761
		x"50",	--8762
		x"00",	--8763
		x"41",	--8764
		x"c3",	--8765
		x"10",	--8766
		x"10",	--8767
		x"53",	--8768
		x"23",	--8769
		x"3f",	--8770
		x"43",	--8771
		x"40",	--8772
		x"80",	--8773
		x"50",	--8774
		x"00",	--8775
		x"41",	--8776
		x"12",	--8777
		x"12",	--8778
		x"12",	--8779
		x"12",	--8780
		x"82",	--8781
		x"4e",	--8782
		x"4f",	--8783
		x"43",	--8784
		x"00",	--8785
		x"93",	--8786
		x"20",	--8787
		x"93",	--8788
		x"20",	--8789
		x"43",	--8790
		x"00",	--8791
		x"41",	--8792
		x"12",	--8793
		x"c5",	--8794
		x"52",	--8795
		x"41",	--8796
		x"41",	--8797
		x"41",	--8798
		x"41",	--8799
		x"41",	--8800
		x"40",	--8801
		x"00",	--8802
		x"00",	--8803
		x"40",	--8804
		x"00",	--8805
		x"00",	--8806
		x"4a",	--8807
		x"00",	--8808
		x"4b",	--8809
		x"00",	--8810
		x"4a",	--8811
		x"4b",	--8812
		x"12",	--8813
		x"c5",	--8814
		x"53",	--8815
		x"93",	--8816
		x"38",	--8817
		x"27",	--8818
		x"4a",	--8819
		x"00",	--8820
		x"4b",	--8821
		x"00",	--8822
		x"4f",	--8823
		x"f0",	--8824
		x"00",	--8825
		x"20",	--8826
		x"40",	--8827
		x"00",	--8828
		x"8f",	--8829
		x"4e",	--8830
		x"00",	--8831
		x"3f",	--8832
		x"51",	--8833
		x"00",	--8834
		x"00",	--8835
		x"61",	--8836
		x"00",	--8837
		x"00",	--8838
		x"53",	--8839
		x"23",	--8840
		x"3f",	--8841
		x"4f",	--8842
		x"e3",	--8843
		x"53",	--8844
		x"43",	--8845
		x"43",	--8846
		x"4e",	--8847
		x"f0",	--8848
		x"00",	--8849
		x"24",	--8850
		x"5c",	--8851
		x"6d",	--8852
		x"53",	--8853
		x"23",	--8854
		x"53",	--8855
		x"63",	--8856
		x"fa",	--8857
		x"fb",	--8858
		x"43",	--8859
		x"43",	--8860
		x"93",	--8861
		x"20",	--8862
		x"93",	--8863
		x"20",	--8864
		x"43",	--8865
		x"43",	--8866
		x"f0",	--8867
		x"00",	--8868
		x"20",	--8869
		x"48",	--8870
		x"49",	--8871
		x"da",	--8872
		x"db",	--8873
		x"4d",	--8874
		x"00",	--8875
		x"4e",	--8876
		x"00",	--8877
		x"40",	--8878
		x"00",	--8879
		x"8f",	--8880
		x"4e",	--8881
		x"00",	--8882
		x"3f",	--8883
		x"c3",	--8884
		x"10",	--8885
		x"10",	--8886
		x"53",	--8887
		x"23",	--8888
		x"3f",	--8889
		x"12",	--8890
		x"12",	--8891
		x"12",	--8892
		x"93",	--8893
		x"2c",	--8894
		x"90",	--8895
		x"01",	--8896
		x"28",	--8897
		x"40",	--8898
		x"00",	--8899
		x"43",	--8900
		x"42",	--8901
		x"4e",	--8902
		x"4f",	--8903
		x"49",	--8904
		x"93",	--8905
		x"20",	--8906
		x"50",	--8907
		x"dc",	--8908
		x"4c",	--8909
		x"43",	--8910
		x"8e",	--8911
		x"7f",	--8912
		x"4a",	--8913
		x"41",	--8914
		x"41",	--8915
		x"41",	--8916
		x"41",	--8917
		x"90",	--8918
		x"01",	--8919
		x"28",	--8920
		x"42",	--8921
		x"43",	--8922
		x"40",	--8923
		x"00",	--8924
		x"4e",	--8925
		x"4f",	--8926
		x"49",	--8927
		x"93",	--8928
		x"27",	--8929
		x"c3",	--8930
		x"10",	--8931
		x"10",	--8932
		x"53",	--8933
		x"23",	--8934
		x"3f",	--8935
		x"40",	--8936
		x"00",	--8937
		x"43",	--8938
		x"40",	--8939
		x"00",	--8940
		x"3f",	--8941
		x"40",	--8942
		x"00",	--8943
		x"43",	--8944
		x"43",	--8945
		x"3f",	--8946
		x"12",	--8947
		x"12",	--8948
		x"12",	--8949
		x"12",	--8950
		x"12",	--8951
		x"4f",	--8952
		x"4f",	--8953
		x"00",	--8954
		x"4f",	--8955
		x"00",	--8956
		x"4d",	--8957
		x"00",	--8958
		x"4d",	--8959
		x"93",	--8960
		x"28",	--8961
		x"92",	--8962
		x"24",	--8963
		x"93",	--8964
		x"24",	--8965
		x"93",	--8966
		x"24",	--8967
		x"4d",	--8968
		x"00",	--8969
		x"90",	--8970
		x"ff",	--8971
		x"38",	--8972
		x"90",	--8973
		x"00",	--8974
		x"34",	--8975
		x"4e",	--8976
		x"4f",	--8977
		x"f0",	--8978
		x"00",	--8979
		x"f3",	--8980
		x"90",	--8981
		x"00",	--8982
		x"24",	--8983
		x"50",	--8984
		x"00",	--8985
		x"63",	--8986
		x"93",	--8987
		x"38",	--8988
		x"4b",	--8989
		x"50",	--8990
		x"00",	--8991
		x"c3",	--8992
		x"10",	--8993
		x"10",	--8994
		x"c3",	--8995
		x"10",	--8996
		x"10",	--8997
		x"c3",	--8998
		x"10",	--8999
		x"10",	--9000
		x"c3",	--9001
		x"10",	--9002
		x"10",	--9003
		x"c3",	--9004
		x"10",	--9005
		x"10",	--9006
		x"c3",	--9007
		x"10",	--9008
		x"10",	--9009
		x"c3",	--9010
		x"10",	--9011
		x"10",	--9012
		x"f3",	--9013
		x"f0",	--9014
		x"00",	--9015
		x"4d",	--9016
		x"3c",	--9017
		x"93",	--9018
		x"23",	--9019
		x"43",	--9020
		x"43",	--9021
		x"43",	--9022
		x"4d",	--9023
		x"5d",	--9024
		x"5d",	--9025
		x"5d",	--9026
		x"5d",	--9027
		x"5d",	--9028
		x"5d",	--9029
		x"5d",	--9030
		x"4f",	--9031
		x"f0",	--9032
		x"00",	--9033
		x"dd",	--9034
		x"4a",	--9035
		x"11",	--9036
		x"43",	--9037
		x"10",	--9038
		x"4c",	--9039
		x"df",	--9040
		x"4d",	--9041
		x"41",	--9042
		x"41",	--9043
		x"41",	--9044
		x"41",	--9045
		x"41",	--9046
		x"41",	--9047
		x"93",	--9048
		x"23",	--9049
		x"4e",	--9050
		x"4f",	--9051
		x"f0",	--9052
		x"00",	--9053
		x"f3",	--9054
		x"93",	--9055
		x"20",	--9056
		x"93",	--9057
		x"27",	--9058
		x"50",	--9059
		x"00",	--9060
		x"63",	--9061
		x"3f",	--9062
		x"c3",	--9063
		x"10",	--9064
		x"10",	--9065
		x"4b",	--9066
		x"50",	--9067
		x"00",	--9068
		x"3f",	--9069
		x"43",	--9070
		x"43",	--9071
		x"43",	--9072
		x"3f",	--9073
		x"d3",	--9074
		x"d0",	--9075
		x"00",	--9076
		x"f3",	--9077
		x"f0",	--9078
		x"00",	--9079
		x"43",	--9080
		x"3f",	--9081
		x"40",	--9082
		x"ff",	--9083
		x"8b",	--9084
		x"90",	--9085
		x"00",	--9086
		x"34",	--9087
		x"4e",	--9088
		x"4f",	--9089
		x"47",	--9090
		x"f0",	--9091
		x"00",	--9092
		x"24",	--9093
		x"c3",	--9094
		x"10",	--9095
		x"10",	--9096
		x"53",	--9097
		x"23",	--9098
		x"43",	--9099
		x"43",	--9100
		x"f0",	--9101
		x"00",	--9102
		x"24",	--9103
		x"58",	--9104
		x"69",	--9105
		x"53",	--9106
		x"23",	--9107
		x"53",	--9108
		x"63",	--9109
		x"fe",	--9110
		x"ff",	--9111
		x"43",	--9112
		x"43",	--9113
		x"93",	--9114
		x"20",	--9115
		x"93",	--9116
		x"20",	--9117
		x"43",	--9118
		x"43",	--9119
		x"4e",	--9120
		x"4f",	--9121
		x"dc",	--9122
		x"dd",	--9123
		x"48",	--9124
		x"49",	--9125
		x"f0",	--9126
		x"00",	--9127
		x"f3",	--9128
		x"90",	--9129
		x"00",	--9130
		x"24",	--9131
		x"50",	--9132
		x"00",	--9133
		x"63",	--9134
		x"48",	--9135
		x"49",	--9136
		x"c3",	--9137
		x"10",	--9138
		x"10",	--9139
		x"c3",	--9140
		x"10",	--9141
		x"10",	--9142
		x"c3",	--9143
		x"10",	--9144
		x"10",	--9145
		x"c3",	--9146
		x"10",	--9147
		x"10",	--9148
		x"c3",	--9149
		x"10",	--9150
		x"10",	--9151
		x"c3",	--9152
		x"10",	--9153
		x"10",	--9154
		x"c3",	--9155
		x"10",	--9156
		x"10",	--9157
		x"f3",	--9158
		x"f0",	--9159
		x"00",	--9160
		x"43",	--9161
		x"90",	--9162
		x"40",	--9163
		x"2f",	--9164
		x"43",	--9165
		x"3f",	--9166
		x"43",	--9167
		x"43",	--9168
		x"3f",	--9169
		x"93",	--9170
		x"23",	--9171
		x"48",	--9172
		x"49",	--9173
		x"f0",	--9174
		x"00",	--9175
		x"f3",	--9176
		x"93",	--9177
		x"24",	--9178
		x"50",	--9179
		x"00",	--9180
		x"63",	--9181
		x"3f",	--9182
		x"93",	--9183
		x"27",	--9184
		x"3f",	--9185
		x"12",	--9186
		x"12",	--9187
		x"4f",	--9188
		x"4f",	--9189
		x"00",	--9190
		x"f0",	--9191
		x"00",	--9192
		x"4f",	--9193
		x"00",	--9194
		x"c3",	--9195
		x"10",	--9196
		x"c3",	--9197
		x"10",	--9198
		x"c3",	--9199
		x"10",	--9200
		x"c3",	--9201
		x"10",	--9202
		x"c3",	--9203
		x"10",	--9204
		x"c3",	--9205
		x"10",	--9206
		x"c3",	--9207
		x"10",	--9208
		x"4d",	--9209
		x"4f",	--9210
		x"00",	--9211
		x"b0",	--9212
		x"00",	--9213
		x"43",	--9214
		x"6f",	--9215
		x"4f",	--9216
		x"00",	--9217
		x"93",	--9218
		x"20",	--9219
		x"93",	--9220
		x"24",	--9221
		x"40",	--9222
		x"ff",	--9223
		x"00",	--9224
		x"4a",	--9225
		x"4b",	--9226
		x"5c",	--9227
		x"6d",	--9228
		x"5c",	--9229
		x"6d",	--9230
		x"5c",	--9231
		x"6d",	--9232
		x"5c",	--9233
		x"6d",	--9234
		x"5c",	--9235
		x"6d",	--9236
		x"5c",	--9237
		x"6d",	--9238
		x"5c",	--9239
		x"6d",	--9240
		x"40",	--9241
		x"00",	--9242
		x"00",	--9243
		x"90",	--9244
		x"40",	--9245
		x"2c",	--9246
		x"40",	--9247
		x"ff",	--9248
		x"5c",	--9249
		x"6d",	--9250
		x"4f",	--9251
		x"53",	--9252
		x"90",	--9253
		x"40",	--9254
		x"2b",	--9255
		x"4a",	--9256
		x"00",	--9257
		x"4c",	--9258
		x"00",	--9259
		x"4d",	--9260
		x"00",	--9261
		x"41",	--9262
		x"41",	--9263
		x"41",	--9264
		x"90",	--9265
		x"00",	--9266
		x"24",	--9267
		x"50",	--9268
		x"ff",	--9269
		x"4d",	--9270
		x"00",	--9271
		x"40",	--9272
		x"00",	--9273
		x"00",	--9274
		x"4a",	--9275
		x"4b",	--9276
		x"5c",	--9277
		x"6d",	--9278
		x"5c",	--9279
		x"6d",	--9280
		x"5c",	--9281
		x"6d",	--9282
		x"5c",	--9283
		x"6d",	--9284
		x"5c",	--9285
		x"6d",	--9286
		x"5c",	--9287
		x"6d",	--9288
		x"5c",	--9289
		x"6d",	--9290
		x"4c",	--9291
		x"4d",	--9292
		x"d3",	--9293
		x"d0",	--9294
		x"40",	--9295
		x"4a",	--9296
		x"00",	--9297
		x"4b",	--9298
		x"00",	--9299
		x"41",	--9300
		x"41",	--9301
		x"41",	--9302
		x"93",	--9303
		x"23",	--9304
		x"43",	--9305
		x"00",	--9306
		x"41",	--9307
		x"41",	--9308
		x"41",	--9309
		x"93",	--9310
		x"24",	--9311
		x"4a",	--9312
		x"4b",	--9313
		x"f3",	--9314
		x"f0",	--9315
		x"00",	--9316
		x"93",	--9317
		x"20",	--9318
		x"93",	--9319
		x"24",	--9320
		x"43",	--9321
		x"00",	--9322
		x"3f",	--9323
		x"93",	--9324
		x"23",	--9325
		x"42",	--9326
		x"00",	--9327
		x"3f",	--9328
		x"43",	--9329
		x"00",	--9330
		x"3f",	--9331
		x"12",	--9332
		x"4f",	--9333
		x"93",	--9334
		x"28",	--9335
		x"4e",	--9336
		x"93",	--9337
		x"28",	--9338
		x"92",	--9339
		x"24",	--9340
		x"92",	--9341
		x"24",	--9342
		x"93",	--9343
		x"24",	--9344
		x"93",	--9345
		x"24",	--9346
		x"4f",	--9347
		x"00",	--9348
		x"9e",	--9349
		x"00",	--9350
		x"24",	--9351
		x"93",	--9352
		x"20",	--9353
		x"43",	--9354
		x"4e",	--9355
		x"41",	--9356
		x"41",	--9357
		x"93",	--9358
		x"24",	--9359
		x"93",	--9360
		x"00",	--9361
		x"23",	--9362
		x"43",	--9363
		x"4e",	--9364
		x"41",	--9365
		x"41",	--9366
		x"93",	--9367
		x"00",	--9368
		x"27",	--9369
		x"43",	--9370
		x"3f",	--9371
		x"4f",	--9372
		x"00",	--9373
		x"4e",	--9374
		x"00",	--9375
		x"9b",	--9376
		x"3b",	--9377
		x"9c",	--9378
		x"38",	--9379
		x"4f",	--9380
		x"00",	--9381
		x"4f",	--9382
		x"00",	--9383
		x"4e",	--9384
		x"00",	--9385
		x"4e",	--9386
		x"00",	--9387
		x"9f",	--9388
		x"2b",	--9389
		x"9e",	--9390
		x"28",	--9391
		x"9b",	--9392
		x"2b",	--9393
		x"9e",	--9394
		x"28",	--9395
		x"9f",	--9396
		x"28",	--9397
		x"9c",	--9398
		x"28",	--9399
		x"43",	--9400
		x"3f",	--9401
		x"93",	--9402
		x"23",	--9403
		x"43",	--9404
		x"3f",	--9405
		x"92",	--9406
		x"23",	--9407
		x"4e",	--9408
		x"00",	--9409
		x"4f",	--9410
		x"00",	--9411
		x"8f",	--9412
		x"3f",	--9413
		x"42",	--9414
		x"02",	--9415
		x"93",	--9416
		x"38",	--9417
		x"42",	--9418
		x"02",	--9419
		x"4f",	--9420
		x"00",	--9421
		x"53",	--9422
		x"4d",	--9423
		x"02",	--9424
		x"53",	--9425
		x"4e",	--9426
		x"02",	--9427
		x"41",	--9428
		x"43",	--9429
		x"41",	--9430
		x"12",	--9431
		x"12",	--9432
		x"83",	--9433
		x"4e",	--9434
		x"00",	--9435
		x"42",	--9436
		x"02",	--9437
		x"42",	--9438
		x"02",	--9439
		x"4e",	--9440
		x"4f",	--9441
		x"40",	--9442
		x"c9",	--9443
		x"12",	--9444
		x"cb",	--9445
		x"9b",	--9446
		x"38",	--9447
		x"4a",	--9448
		x"5b",	--9449
		x"43",	--9450
		x"ff",	--9451
		x"3c",	--9452
		x"42",	--9453
		x"02",	--9454
		x"43",	--9455
		x"00",	--9456
		x"53",	--9457
		x"41",	--9458
		x"41",	--9459
		x"41",	--9460
		x"41",	--9461
		x"00",	--9462
		x"02",	--9463
		x"40",	--9464
		x"7f",	--9465
		x"02",	--9466
		x"41",	--9467
		x"50",	--9468
		x"00",	--9469
		x"41",	--9470
		x"00",	--9471
		x"12",	--9472
		x"c9",	--9473
		x"41",	--9474
		x"41",	--9475
		x"00",	--9476
		x"02",	--9477
		x"41",	--9478
		x"00",	--9479
		x"02",	--9480
		x"41",	--9481
		x"52",	--9482
		x"41",	--9483
		x"00",	--9484
		x"12",	--9485
		x"c9",	--9486
		x"41",	--9487
		x"4e",	--9488
		x"4f",	--9489
		x"02",	--9490
		x"40",	--9491
		x"7f",	--9492
		x"02",	--9493
		x"4d",	--9494
		x"4c",	--9495
		x"12",	--9496
		x"c9",	--9497
		x"41",	--9498
		x"4f",	--9499
		x"02",	--9500
		x"4e",	--9501
		x"02",	--9502
		x"4c",	--9503
		x"4d",	--9504
		x"12",	--9505
		x"c9",	--9506
		x"41",	--9507
		x"12",	--9508
		x"12",	--9509
		x"12",	--9510
		x"12",	--9511
		x"12",	--9512
		x"12",	--9513
		x"12",	--9514
		x"12",	--9515
		x"82",	--9516
		x"4f",	--9517
		x"4e",	--9518
		x"00",	--9519
		x"4d",	--9520
		x"41",	--9521
		x"00",	--9522
		x"41",	--9523
		x"00",	--9524
		x"4d",	--9525
		x"4d",	--9526
		x"10",	--9527
		x"44",	--9528
		x"4f",	--9529
		x"b0",	--9530
		x"00",	--9531
		x"24",	--9532
		x"40",	--9533
		x"00",	--9534
		x"00",	--9535
		x"4f",	--9536
		x"10",	--9537
		x"f3",	--9538
		x"24",	--9539
		x"40",	--9540
		x"00",	--9541
		x"3c",	--9542
		x"40",	--9543
		x"00",	--9544
		x"4e",	--9545
		x"00",	--9546
		x"41",	--9547
		x"53",	--9548
		x"3c",	--9549
		x"f0",	--9550
		x"00",	--9551
		x"24",	--9552
		x"40",	--9553
		x"00",	--9554
		x"00",	--9555
		x"3c",	--9556
		x"93",	--9557
		x"24",	--9558
		x"4d",	--9559
		x"00",	--9560
		x"41",	--9561
		x"53",	--9562
		x"3c",	--9563
		x"41",	--9564
		x"4c",	--9565
		x"10",	--9566
		x"11",	--9567
		x"10",	--9568
		x"11",	--9569
		x"4c",	--9570
		x"41",	--9571
		x"41",	--9572
		x"10",	--9573
		x"11",	--9574
		x"10",	--9575
		x"11",	--9576
		x"4c",	--9577
		x"86",	--9578
		x"77",	--9579
		x"4f",	--9580
		x"10",	--9581
		x"4e",	--9582
		x"00",	--9583
		x"f2",	--9584
		x"24",	--9585
		x"45",	--9586
		x"3c",	--9587
		x"43",	--9588
		x"4f",	--9589
		x"b0",	--9590
		x"00",	--9591
		x"20",	--9592
		x"41",	--9593
		x"00",	--9594
		x"53",	--9595
		x"53",	--9596
		x"93",	--9597
		x"00",	--9598
		x"23",	--9599
		x"81",	--9600
		x"00",	--9601
		x"9a",	--9602
		x"28",	--9603
		x"8a",	--9604
		x"3c",	--9605
		x"43",	--9606
		x"b3",	--9607
		x"00",	--9608
		x"24",	--9609
		x"95",	--9610
		x"28",	--9611
		x"85",	--9612
		x"3c",	--9613
		x"43",	--9614
		x"4d",	--9615
		x"9d",	--9616
		x"2c",	--9617
		x"47",	--9618
		x"93",	--9619
		x"38",	--9620
		x"40",	--9621
		x"00",	--9622
		x"00",	--9623
		x"43",	--9624
		x"43",	--9625
		x"3c",	--9626
		x"41",	--9627
		x"56",	--9628
		x"4f",	--9629
		x"11",	--9630
		x"53",	--9631
		x"12",	--9632
		x"3c",	--9633
		x"43",	--9634
		x"9a",	--9635
		x"3b",	--9636
		x"4a",	--9637
		x"40",	--9638
		x"00",	--9639
		x"00",	--9640
		x"8b",	--9641
		x"3c",	--9642
		x"41",	--9643
		x"00",	--9644
		x"11",	--9645
		x"12",	--9646
		x"53",	--9647
		x"45",	--9648
		x"5b",	--9649
		x"99",	--9650
		x"2b",	--9651
		x"3c",	--9652
		x"43",	--9653
		x"43",	--9654
		x"3c",	--9655
		x"53",	--9656
		x"41",	--9657
		x"56",	--9658
		x"4f",	--9659
		x"11",	--9660
		x"53",	--9661
		x"12",	--9662
		x"9a",	--9663
		x"3b",	--9664
		x"b3",	--9665
		x"00",	--9666
		x"24",	--9667
		x"44",	--9668
		x"3c",	--9669
		x"41",	--9670
		x"00",	--9671
		x"8b",	--9672
		x"3c",	--9673
		x"40",	--9674
		x"00",	--9675
		x"12",	--9676
		x"53",	--9677
		x"93",	--9678
		x"23",	--9679
		x"44",	--9680
		x"54",	--9681
		x"3f",	--9682
		x"53",	--9683
		x"11",	--9684
		x"12",	--9685
		x"53",	--9686
		x"4a",	--9687
		x"5b",	--9688
		x"4f",	--9689
		x"93",	--9690
		x"24",	--9691
		x"93",	--9692
		x"23",	--9693
		x"3c",	--9694
		x"40",	--9695
		x"00",	--9696
		x"12",	--9697
		x"53",	--9698
		x"99",	--9699
		x"2b",	--9700
		x"4b",	--9701
		x"52",	--9702
		x"41",	--9703
		x"41",	--9704
		x"41",	--9705
		x"41",	--9706
		x"41",	--9707
		x"41",	--9708
		x"41",	--9709
		x"41",	--9710
		x"41",	--9711
		x"12",	--9712
		x"12",	--9713
		x"12",	--9714
		x"12",	--9715
		x"12",	--9716
		x"12",	--9717
		x"12",	--9718
		x"12",	--9719
		x"50",	--9720
		x"ff",	--9721
		x"4f",	--9722
		x"00",	--9723
		x"4e",	--9724
		x"4d",	--9725
		x"4e",	--9726
		x"00",	--9727
		x"43",	--9728
		x"00",	--9729
		x"43",	--9730
		x"00",	--9731
		x"43",	--9732
		x"00",	--9733
		x"43",	--9734
		x"00",	--9735
		x"43",	--9736
		x"00",	--9737
		x"43",	--9738
		x"00",	--9739
		x"43",	--9740
		x"43",	--9741
		x"00",	--9742
		x"41",	--9743
		x"50",	--9744
		x"00",	--9745
		x"4e",	--9746
		x"00",	--9747
		x"40",	--9748
		x"d2",	--9749
		x"46",	--9750
		x"53",	--9751
		x"4f",	--9752
		x"00",	--9753
		x"93",	--9754
		x"20",	--9755
		x"90",	--9756
		x"00",	--9757
		x"20",	--9758
		x"43",	--9759
		x"00",	--9760
		x"43",	--9761
		x"00",	--9762
		x"46",	--9763
		x"00",	--9764
		x"43",	--9765
		x"00",	--9766
		x"43",	--9767
		x"00",	--9768
		x"43",	--9769
		x"00",	--9770
		x"43",	--9771
		x"00",	--9772
		x"43",	--9773
		x"00",	--9774
		x"40",	--9775
		x"d2",	--9776
		x"47",	--9777
		x"11",	--9778
		x"4e",	--9779
		x"12",	--9780
		x"00",	--9781
		x"53",	--9782
		x"00",	--9783
		x"40",	--9784
		x"d2",	--9785
		x"90",	--9786
		x"00",	--9787
		x"24",	--9788
		x"90",	--9789
		x"00",	--9790
		x"34",	--9791
		x"90",	--9792
		x"00",	--9793
		x"24",	--9794
		x"90",	--9795
		x"00",	--9796
		x"34",	--9797
		x"90",	--9798
		x"00",	--9799
		x"24",	--9800
		x"90",	--9801
		x"00",	--9802
		x"34",	--9803
		x"90",	--9804
		x"00",	--9805
		x"24",	--9806
		x"90",	--9807
		x"00",	--9808
		x"27",	--9809
		x"90",	--9810
		x"00",	--9811
		x"20",	--9812
		x"3c",	--9813
		x"90",	--9814
		x"00",	--9815
		x"24",	--9816
		x"90",	--9817
		x"00",	--9818
		x"24",	--9819
		x"90",	--9820
		x"00",	--9821
		x"20",	--9822
		x"3c",	--9823
		x"90",	--9824
		x"00",	--9825
		x"38",	--9826
		x"90",	--9827
		x"00",	--9828
		x"20",	--9829
		x"3c",	--9830
		x"90",	--9831
		x"00",	--9832
		x"24",	--9833
		x"90",	--9834
		x"00",	--9835
		x"34",	--9836
		x"90",	--9837
		x"00",	--9838
		x"24",	--9839
		x"90",	--9840
		x"00",	--9841
		x"24",	--9842
		x"90",	--9843
		x"00",	--9844
		x"20",	--9845
		x"3c",	--9846
		x"90",	--9847
		x"00",	--9848
		x"24",	--9849
		x"90",	--9850
		x"00",	--9851
		x"34",	--9852
		x"90",	--9853
		x"00",	--9854
		x"20",	--9855
		x"3c",	--9856
		x"90",	--9857
		x"00",	--9858
		x"24",	--9859
		x"90",	--9860
		x"00",	--9861
		x"24",	--9862
		x"41",	--9863
		x"00",	--9864
		x"41",	--9865
		x"00",	--9866
		x"89",	--9867
		x"40",	--9868
		x"d2",	--9869
		x"42",	--9870
		x"00",	--9871
		x"3c",	--9872
		x"d2",	--9873
		x"00",	--9874
		x"40",	--9875
		x"d2",	--9876
		x"41",	--9877
		x"f3",	--9878
		x"41",	--9879
		x"24",	--9880
		x"f0",	--9881
		x"ff",	--9882
		x"d3",	--9883
		x"3c",	--9884
		x"d3",	--9885
		x"4e",	--9886
		x"00",	--9887
		x"40",	--9888
		x"d2",	--9889
		x"d0",	--9890
		x"00",	--9891
		x"00",	--9892
		x"40",	--9893
		x"d2",	--9894
		x"40",	--9895
		x"00",	--9896
		x"00",	--9897
		x"40",	--9898
		x"d2",	--9899
		x"90",	--9900
		x"00",	--9901
		x"00",	--9902
		x"20",	--9903
		x"40",	--9904
		x"d2",	--9905
		x"40",	--9906
		x"00",	--9907
		x"00",	--9908
		x"40",	--9909
		x"d2",	--9910
		x"93",	--9911
		x"00",	--9912
		x"24",	--9913
		x"40",	--9914
		x"d2",	--9915
		x"43",	--9916
		x"00",	--9917
		x"40",	--9918
		x"d2",	--9919
		x"45",	--9920
		x"53",	--9921
		x"45",	--9922
		x"93",	--9923
		x"38",	--9924
		x"4a",	--9925
		x"00",	--9926
		x"3c",	--9927
		x"93",	--9928
		x"00",	--9929
		x"24",	--9930
		x"40",	--9931
		x"d2",	--9932
		x"d0",	--9933
		x"00",	--9934
		x"00",	--9935
		x"e3",	--9936
		x"4a",	--9937
		x"00",	--9938
		x"53",	--9939
		x"00",	--9940
		x"4e",	--9941
		x"3c",	--9942
		x"93",	--9943
		x"00",	--9944
		x"20",	--9945
		x"93",	--9946
		x"00",	--9947
		x"20",	--9948
		x"41",	--9949
		x"f0",	--9950
		x"00",	--9951
		x"43",	--9952
		x"24",	--9953
		x"43",	--9954
		x"4e",	--9955
		x"11",	--9956
		x"43",	--9957
		x"10",	--9958
		x"41",	--9959
		x"f0",	--9960
		x"00",	--9961
		x"de",	--9962
		x"4a",	--9963
		x"00",	--9964
		x"40",	--9965
		x"d2",	--9966
		x"41",	--9967
		x"00",	--9968
		x"5a",	--9969
		x"4a",	--9970
		x"5c",	--9971
		x"5c",	--9972
		x"5c",	--9973
		x"4a",	--9974
		x"00",	--9975
		x"50",	--9976
		x"ff",	--9977
		x"00",	--9978
		x"11",	--9979
		x"5e",	--9980
		x"00",	--9981
		x"43",	--9982
		x"00",	--9983
		x"40",	--9984
		x"d2",	--9985
		x"45",	--9986
		x"53",	--9987
		x"45",	--9988
		x"93",	--9989
		x"00",	--9990
		x"20",	--9991
		x"93",	--9992
		x"00",	--9993
		x"27",	--9994
		x"4e",	--9995
		x"00",	--9996
		x"43",	--9997
		x"00",	--9998
		x"41",	--9999
		x"52",	--10000
		x"3c",	--10001
		x"45",	--10002
		x"53",	--10003
		x"45",	--10004
		x"93",	--10005
		x"00",	--10006
		x"24",	--10007
		x"d2",	--10008
		x"00",	--10009
		x"41",	--10010
		x"00",	--10011
		x"4f",	--10012
		x"00",	--10013
		x"3c",	--10014
		x"93",	--10015
		x"00",	--10016
		x"24",	--10017
		x"41",	--10018
		x"00",	--10019
		x"00",	--10020
		x"93",	--10021
		x"20",	--10022
		x"40",	--10023
		x"dd",	--10024
		x"12",	--10025
		x"00",	--10026
		x"12",	--10027
		x"00",	--10028
		x"41",	--10029
		x"00",	--10030
		x"41",	--10031
		x"00",	--10032
		x"12",	--10033
		x"ca",	--10034
		x"52",	--10035
		x"5f",	--10036
		x"00",	--10037
		x"47",	--10038
		x"40",	--10039
		x"d2",	--10040
		x"45",	--10041
		x"53",	--10042
		x"45",	--10043
		x"49",	--10044
		x"00",	--10045
		x"43",	--10046
		x"93",	--10047
		x"20",	--10048
		x"43",	--10049
		x"5e",	--10050
		x"5e",	--10051
		x"5e",	--10052
		x"41",	--10053
		x"f0",	--10054
		x"ff",	--10055
		x"de",	--10056
		x"4a",	--10057
		x"00",	--10058
		x"47",	--10059
		x"40",	--10060
		x"00",	--10061
		x"00",	--10062
		x"3c",	--10063
		x"d3",	--10064
		x"00",	--10065
		x"3c",	--10066
		x"d2",	--10067
		x"00",	--10068
		x"40",	--10069
		x"00",	--10070
		x"00",	--10071
		x"3c",	--10072
		x"40",	--10073
		x"00",	--10074
		x"00",	--10075
		x"41",	--10076
		x"b3",	--10077
		x"24",	--10078
		x"45",	--10079
		x"52",	--10080
		x"45",	--10081
		x"45",	--10082
		x"00",	--10083
		x"45",	--10084
		x"00",	--10085
		x"45",	--10086
		x"00",	--10087
		x"48",	--10088
		x"00",	--10089
		x"47",	--10090
		x"00",	--10091
		x"46",	--10092
		x"00",	--10093
		x"4b",	--10094
		x"00",	--10095
		x"43",	--10096
		x"00",	--10097
		x"93",	--10098
		x"20",	--10099
		x"93",	--10100
		x"20",	--10101
		x"93",	--10102
		x"20",	--10103
		x"93",	--10104
		x"24",	--10105
		x"43",	--10106
		x"00",	--10107
		x"5b",	--10108
		x"43",	--10109
		x"6b",	--10110
		x"4b",	--10111
		x"00",	--10112
		x"4c",	--10113
		x"3c",	--10114
		x"f3",	--10115
		x"45",	--10116
		x"24",	--10117
		x"52",	--10118
		x"45",	--10119
		x"45",	--10120
		x"00",	--10121
		x"48",	--10122
		x"00",	--10123
		x"4b",	--10124
		x"00",	--10125
		x"43",	--10126
		x"00",	--10127
		x"93",	--10128
		x"20",	--10129
		x"3c",	--10130
		x"53",	--10131
		x"45",	--10132
		x"4b",	--10133
		x"00",	--10134
		x"43",	--10135
		x"00",	--10136
		x"93",	--10137
		x"24",	--10138
		x"43",	--10139
		x"00",	--10140
		x"5b",	--10141
		x"43",	--10142
		x"6b",	--10143
		x"4b",	--10144
		x"00",	--10145
		x"47",	--10146
		x"b2",	--10147
		x"00",	--10148
		x"24",	--10149
		x"93",	--10150
		x"00",	--10151
		x"20",	--10152
		x"41",	--10153
		x"90",	--10154
		x"00",	--10155
		x"00",	--10156
		x"20",	--10157
		x"d0",	--10158
		x"00",	--10159
		x"3c",	--10160
		x"92",	--10161
		x"00",	--10162
		x"20",	--10163
		x"d0",	--10164
		x"00",	--10165
		x"48",	--10166
		x"00",	--10167
		x"41",	--10168
		x"b2",	--10169
		x"24",	--10170
		x"93",	--10171
		x"00",	--10172
		x"24",	--10173
		x"40",	--10174
		x"00",	--10175
		x"00",	--10176
		x"b3",	--10177
		x"24",	--10178
		x"e3",	--10179
		x"00",	--10180
		x"e3",	--10181
		x"00",	--10182
		x"e3",	--10183
		x"00",	--10184
		x"e3",	--10185
		x"00",	--10186
		x"53",	--10187
		x"00",	--10188
		x"63",	--10189
		x"00",	--10190
		x"63",	--10191
		x"00",	--10192
		x"63",	--10193
		x"00",	--10194
		x"3c",	--10195
		x"b3",	--10196
		x"24",	--10197
		x"41",	--10198
		x"00",	--10199
		x"41",	--10200
		x"00",	--10201
		x"e3",	--10202
		x"e3",	--10203
		x"4a",	--10204
		x"4b",	--10205
		x"53",	--10206
		x"63",	--10207
		x"4e",	--10208
		x"00",	--10209
		x"4f",	--10210
		x"00",	--10211
		x"3c",	--10212
		x"41",	--10213
		x"00",	--10214
		x"e3",	--10215
		x"53",	--10216
		x"4a",	--10217
		x"00",	--10218
		x"43",	--10219
		x"00",	--10220
		x"b3",	--10221
		x"24",	--10222
		x"41",	--10223
		x"00",	--10224
		x"41",	--10225
		x"00",	--10226
		x"00",	--10227
		x"41",	--10228
		x"00",	--10229
		x"41",	--10230
		x"00",	--10231
		x"41",	--10232
		x"50",	--10233
		x"00",	--10234
		x"46",	--10235
		x"41",	--10236
		x"00",	--10237
		x"00",	--10238
		x"41",	--10239
		x"00",	--10240
		x"10",	--10241
		x"11",	--10242
		x"10",	--10243
		x"11",	--10244
		x"4b",	--10245
		x"00",	--10246
		x"4b",	--10247
		x"00",	--10248
		x"4b",	--10249
		x"00",	--10250
		x"12",	--10251
		x"00",	--10252
		x"12",	--10253
		x"00",	--10254
		x"12",	--10255
		x"00",	--10256
		x"12",	--10257
		x"00",	--10258
		x"49",	--10259
		x"41",	--10260
		x"00",	--10261
		x"48",	--10262
		x"44",	--10263
		x"12",	--10264
		x"d3",	--10265
		x"52",	--10266
		x"4c",	--10267
		x"90",	--10268
		x"00",	--10269
		x"34",	--10270
		x"50",	--10271
		x"00",	--10272
		x"4b",	--10273
		x"00",	--10274
		x"3c",	--10275
		x"4c",	--10276
		x"b3",	--10277
		x"00",	--10278
		x"24",	--10279
		x"40",	--10280
		x"00",	--10281
		x"3c",	--10282
		x"40",	--10283
		x"00",	--10284
		x"5b",	--10285
		x"4a",	--10286
		x"00",	--10287
		x"47",	--10288
		x"53",	--10289
		x"12",	--10290
		x"00",	--10291
		x"12",	--10292
		x"00",	--10293
		x"12",	--10294
		x"00",	--10295
		x"12",	--10296
		x"00",	--10297
		x"49",	--10298
		x"41",	--10299
		x"00",	--10300
		x"48",	--10301
		x"44",	--10302
		x"12",	--10303
		x"d3",	--10304
		x"52",	--10305
		x"4c",	--10306
		x"4d",	--10307
		x"00",	--10308
		x"4e",	--10309
		x"4f",	--10310
		x"53",	--10311
		x"93",	--10312
		x"23",	--10313
		x"93",	--10314
		x"23",	--10315
		x"93",	--10316
		x"23",	--10317
		x"93",	--10318
		x"23",	--10319
		x"43",	--10320
		x"00",	--10321
		x"43",	--10322
		x"00",	--10323
		x"43",	--10324
		x"00",	--10325
		x"43",	--10326
		x"00",	--10327
		x"3c",	--10328
		x"b3",	--10329
		x"24",	--10330
		x"41",	--10331
		x"00",	--10332
		x"41",	--10333
		x"00",	--10334
		x"41",	--10335
		x"50",	--10336
		x"00",	--10337
		x"41",	--10338
		x"00",	--10339
		x"10",	--10340
		x"11",	--10341
		x"10",	--10342
		x"11",	--10343
		x"41",	--10344
		x"00",	--10345
		x"49",	--10346
		x"44",	--10347
		x"47",	--10348
		x"12",	--10349
		x"d2",	--10350
		x"4e",	--10351
		x"90",	--10352
		x"00",	--10353
		x"34",	--10354
		x"50",	--10355
		x"00",	--10356
		x"4b",	--10357
		x"00",	--10358
		x"3c",	--10359
		x"4e",	--10360
		x"b3",	--10361
		x"00",	--10362
		x"24",	--10363
		x"40",	--10364
		x"00",	--10365
		x"3c",	--10366
		x"40",	--10367
		x"00",	--10368
		x"5b",	--10369
		x"4a",	--10370
		x"00",	--10371
		x"48",	--10372
		x"53",	--10373
		x"41",	--10374
		x"00",	--10375
		x"49",	--10376
		x"44",	--10377
		x"47",	--10378
		x"12",	--10379
		x"d2",	--10380
		x"4e",	--10381
		x"4f",	--10382
		x"53",	--10383
		x"93",	--10384
		x"23",	--10385
		x"93",	--10386
		x"23",	--10387
		x"43",	--10388
		x"00",	--10389
		x"43",	--10390
		x"00",	--10391
		x"3c",	--10392
		x"41",	--10393
		x"00",	--10394
		x"41",	--10395
		x"50",	--10396
		x"00",	--10397
		x"41",	--10398
		x"00",	--10399
		x"47",	--10400
		x"12",	--10401
		x"d3",	--10402
		x"4f",	--10403
		x"90",	--10404
		x"00",	--10405
		x"34",	--10406
		x"50",	--10407
		x"00",	--10408
		x"4d",	--10409
		x"00",	--10410
		x"3c",	--10411
		x"4f",	--10412
		x"b3",	--10413
		x"00",	--10414
		x"24",	--10415
		x"40",	--10416
		x"00",	--10417
		x"3c",	--10418
		x"40",	--10419
		x"00",	--10420
		x"5d",	--10421
		x"4c",	--10422
		x"00",	--10423
		x"48",	--10424
		x"53",	--10425
		x"41",	--10426
		x"00",	--10427
		x"47",	--10428
		x"12",	--10429
		x"d3",	--10430
		x"4f",	--10431
		x"53",	--10432
		x"93",	--10433
		x"23",	--10434
		x"43",	--10435
		x"00",	--10436
		x"90",	--10437
		x"00",	--10438
		x"00",	--10439
		x"24",	--10440
		x"43",	--10441
		x"00",	--10442
		x"93",	--10443
		x"00",	--10444
		x"24",	--10445
		x"41",	--10446
		x"50",	--10447
		x"00",	--10448
		x"4f",	--10449
		x"00",	--10450
		x"41",	--10451
		x"00",	--10452
		x"10",	--10453
		x"11",	--10454
		x"10",	--10455
		x"11",	--10456
		x"4a",	--10457
		x"00",	--10458
		x"46",	--10459
		x"00",	--10460
		x"46",	--10461
		x"10",	--10462
		x"11",	--10463
		x"10",	--10464
		x"11",	--10465
		x"4a",	--10466
		x"00",	--10467
		x"41",	--10468
		x"00",	--10469
		x"41",	--10470
		x"00",	--10471
		x"81",	--10472
		x"00",	--10473
		x"71",	--10474
		x"00",	--10475
		x"83",	--10476
		x"91",	--10477
		x"00",	--10478
		x"2c",	--10479
		x"d3",	--10480
		x"00",	--10481
		x"41",	--10482
		x"00",	--10483
		x"8c",	--10484
		x"4e",	--10485
		x"00",	--10486
		x"3c",	--10487
		x"93",	--10488
		x"00",	--10489
		x"24",	--10490
		x"41",	--10491
		x"00",	--10492
		x"00",	--10493
		x"12",	--10494
		x"00",	--10495
		x"12",	--10496
		x"00",	--10497
		x"41",	--10498
		x"00",	--10499
		x"46",	--10500
		x"53",	--10501
		x"41",	--10502
		x"00",	--10503
		x"12",	--10504
		x"ca",	--10505
		x"52",	--10506
		x"5f",	--10507
		x"00",	--10508
		x"3c",	--10509
		x"49",	--10510
		x"11",	--10511
		x"12",	--10512
		x"00",	--10513
		x"49",	--10514
		x"58",	--10515
		x"91",	--10516
		x"00",	--10517
		x"2b",	--10518
		x"49",	--10519
		x"00",	--10520
		x"4e",	--10521
		x"00",	--10522
		x"43",	--10523
		x"3c",	--10524
		x"41",	--10525
		x"00",	--10526
		x"00",	--10527
		x"43",	--10528
		x"00",	--10529
		x"43",	--10530
		x"00",	--10531
		x"3c",	--10532
		x"4e",	--10533
		x"43",	--10534
		x"00",	--10535
		x"43",	--10536
		x"00",	--10537
		x"43",	--10538
		x"41",	--10539
		x"00",	--10540
		x"46",	--10541
		x"93",	--10542
		x"24",	--10543
		x"40",	--10544
		x"cc",	--10545
		x"41",	--10546
		x"00",	--10547
		x"50",	--10548
		x"00",	--10549
		x"41",	--10550
		x"41",	--10551
		x"41",	--10552
		x"41",	--10553
		x"41",	--10554
		x"41",	--10555
		x"41",	--10556
		x"41",	--10557
		x"41",	--10558
		x"43",	--10559
		x"93",	--10560
		x"34",	--10561
		x"40",	--10562
		x"00",	--10563
		x"e3",	--10564
		x"53",	--10565
		x"93",	--10566
		x"34",	--10567
		x"e3",	--10568
		x"e3",	--10569
		x"53",	--10570
		x"12",	--10571
		x"12",	--10572
		x"d3",	--10573
		x"41",	--10574
		x"b3",	--10575
		x"24",	--10576
		x"e3",	--10577
		x"53",	--10578
		x"b3",	--10579
		x"24",	--10580
		x"e3",	--10581
		x"53",	--10582
		x"41",	--10583
		x"12",	--10584
		x"d2",	--10585
		x"4e",	--10586
		x"41",	--10587
		x"12",	--10588
		x"12",	--10589
		x"12",	--10590
		x"40",	--10591
		x"00",	--10592
		x"4c",	--10593
		x"4d",	--10594
		x"43",	--10595
		x"43",	--10596
		x"5e",	--10597
		x"6f",	--10598
		x"6c",	--10599
		x"6d",	--10600
		x"9b",	--10601
		x"28",	--10602
		x"20",	--10603
		x"9a",	--10604
		x"28",	--10605
		x"8a",	--10606
		x"7b",	--10607
		x"d3",	--10608
		x"83",	--10609
		x"23",	--10610
		x"41",	--10611
		x"41",	--10612
		x"41",	--10613
		x"41",	--10614
		x"12",	--10615
		x"d2",	--10616
		x"4c",	--10617
		x"4d",	--10618
		x"41",	--10619
		x"12",	--10620
		x"43",	--10621
		x"93",	--10622
		x"34",	--10623
		x"40",	--10624
		x"00",	--10625
		x"e3",	--10626
		x"e3",	--10627
		x"53",	--10628
		x"63",	--10629
		x"93",	--10630
		x"34",	--10631
		x"e3",	--10632
		x"e3",	--10633
		x"e3",	--10634
		x"53",	--10635
		x"63",	--10636
		x"12",	--10637
		x"d2",	--10638
		x"b3",	--10639
		x"24",	--10640
		x"e3",	--10641
		x"e3",	--10642
		x"53",	--10643
		x"63",	--10644
		x"b3",	--10645
		x"24",	--10646
		x"e3",	--10647
		x"e3",	--10648
		x"53",	--10649
		x"63",	--10650
		x"41",	--10651
		x"41",	--10652
		x"12",	--10653
		x"d2",	--10654
		x"4c",	--10655
		x"4d",	--10656
		x"41",	--10657
		x"40",	--10658
		x"00",	--10659
		x"4e",	--10660
		x"43",	--10661
		x"5f",	--10662
		x"6e",	--10663
		x"9d",	--10664
		x"28",	--10665
		x"8d",	--10666
		x"d3",	--10667
		x"83",	--10668
		x"23",	--10669
		x"41",	--10670
		x"12",	--10671
		x"d3",	--10672
		x"4e",	--10673
		x"41",	--10674
		x"12",	--10675
		x"12",	--10676
		x"12",	--10677
		x"12",	--10678
		x"12",	--10679
		x"00",	--10680
		x"48",	--10681
		x"49",	--10682
		x"4a",	--10683
		x"4b",	--10684
		x"43",	--10685
		x"43",	--10686
		x"43",	--10687
		x"43",	--10688
		x"5c",	--10689
		x"6d",	--10690
		x"6e",	--10691
		x"6f",	--10692
		x"68",	--10693
		x"69",	--10694
		x"6a",	--10695
		x"6b",	--10696
		x"97",	--10697
		x"28",	--10698
		x"20",	--10699
		x"96",	--10700
		x"28",	--10701
		x"20",	--10702
		x"95",	--10703
		x"28",	--10704
		x"20",	--10705
		x"94",	--10706
		x"28",	--10707
		x"84",	--10708
		x"75",	--10709
		x"76",	--10710
		x"77",	--10711
		x"d3",	--10712
		x"83",	--10713
		x"00",	--10714
		x"23",	--10715
		x"53",	--10716
		x"41",	--10717
		x"41",	--10718
		x"41",	--10719
		x"41",	--10720
		x"41",	--10721
		x"12",	--10722
		x"12",	--10723
		x"12",	--10724
		x"12",	--10725
		x"41",	--10726
		x"00",	--10727
		x"41",	--10728
		x"00",	--10729
		x"41",	--10730
		x"00",	--10731
		x"41",	--10732
		x"00",	--10733
		x"12",	--10734
		x"d3",	--10735
		x"41",	--10736
		x"41",	--10737
		x"41",	--10738
		x"41",	--10739
		x"41",	--10740
		x"12",	--10741
		x"12",	--10742
		x"12",	--10743
		x"12",	--10744
		x"41",	--10745
		x"00",	--10746
		x"41",	--10747
		x"00",	--10748
		x"41",	--10749
		x"00",	--10750
		x"41",	--10751
		x"00",	--10752
		x"12",	--10753
		x"d3",	--10754
		x"48",	--10755
		x"49",	--10756
		x"4a",	--10757
		x"4b",	--10758
		x"41",	--10759
		x"41",	--10760
		x"41",	--10761
		x"41",	--10762
		x"41",	--10763
		x"12",	--10764
		x"12",	--10765
		x"12",	--10766
		x"12",	--10767
		x"12",	--10768
		x"41",	--10769
		x"00",	--10770
		x"41",	--10771
		x"00",	--10772
		x"41",	--10773
		x"00",	--10774
		x"41",	--10775
		x"00",	--10776
		x"12",	--10777
		x"d3",	--10778
		x"41",	--10779
		x"00",	--10780
		x"48",	--10781
		x"00",	--10782
		x"49",	--10783
		x"00",	--10784
		x"4a",	--10785
		x"00",	--10786
		x"4b",	--10787
		x"00",	--10788
		x"41",	--10789
		x"41",	--10790
		x"41",	--10791
		x"41",	--10792
		x"41",	--10793
		x"41",	--10794
		x"13",	--10795
		x"d0",	--10796
		x"00",	--10797
		x"3f",	--10798
		x"20",	--10799
		x"25",	--10800
		x"20",	--10801
		x"64",	--10802
		x"25",	--10803
		x"00",	--10804
		x"73",	--10805
		x"0a",	--10806
		x"6f",	--10807
		x"00",	--10808
		x"64",	--10809
		x"00",	--10810
		x"0a",	--10811
		x"00",	--10812
		x"85",	--10813
		x"85",	--10814
		x"85",	--10815
		x"85",	--10816
		x"86",	--10817
		x"86",	--10818
		x"85",	--10819
		x"85",	--10820
		x"0a",	--10821
		x"3d",	--10822
		x"3d",	--10823
		x"3d",	--10824
		x"4d",	--10825
		x"72",	--10826
		x"65",	--10827
		x"20",	--10828
		x"43",	--10829
		x"20",	--10830
		x"3d",	--10831
		x"3d",	--10832
		x"3d",	--10833
		x"0a",	--10834
		x"69",	--10835
		x"74",	--10836
		x"72",	--10837
		x"63",	--10838
		x"69",	--10839
		x"65",	--10840
		x"6d",	--10841
		x"64",	--10842
		x"00",	--10843
		x"72",	--10844
		x"74",	--10845
		x"00",	--10846
		x"65",	--10847
		x"64",	--10848
		x"62",	--10849
		x"7a",	--10850
		x"65",	--10851
		x"00",	--10852
		x"77",	--10853
		x"00",	--10854
		x"6e",	--10855
		x"6f",	--10856
		x"65",	--10857
		x"00",	--10858
		x"70",	--10859
		x"65",	--10860
		x"20",	--10861
		x"6f",	--10862
		x"74",	--10863
		x"6f",	--10864
		x"6c",	--10865
		x"72",	--10866
		x"6f",	--10867
		x"6f",	--10868
		x"65",	--10869
		x"72",	--10870
		x"00",	--10871
		x"70",	--10872
		x"65",	--10873
		x"20",	--10874
		x"6f",	--10875
		x"66",	--10876
		x"67",	--10877
		x"72",	--10878
		x"74",	--10879
		x"6f",	--10880
		x"00",	--10881
		x"62",	--10882
		x"74",	--10883
		x"63",	--10884
		x"65",	--10885
		x"61",	--10886
		x"6f",	--10887
		x"64",	--10888
		x"6e",	--10889
		x"65",	--10890
		x"72",	--10891
		x"61",	--10892
		x"00",	--10893
		x"6f",	--10894
		x"74",	--10895
		x"6f",	--10896
		x"64",	--10897
		x"72",	--10898
		x"0d",	--10899
		x"00",	--10900
		x"20",	--10901
		x"00",	--10902
		x"63",	--10903
		x"55",	--10904
		x"0d",	--10905
		x"00",	--10906
		x"4f",	--10907
		x"4e",	--10908
		x"0a",	--10909
		x"52",	--10910
		x"47",	--10911
		x"54",	--10912
		x"0a",	--10913
		x"4c",	--10914
		x"46",	--10915
		x"0d",	--10916
		x"00",	--10917
		x"74",	--10918
		x"70",	--10919
		x"0a",	--10920
		x"63",	--10921
		x"72",	--10922
		x"65",	--10923
		x"74",	--10924
		x"75",	--10925
		x"61",	--10926
		x"65",	--10927
		x"0d",	--10928
		x"00",	--10929
		x"25",	--10930
		x"20",	--10931
		x"6f",	--10932
		x"20",	--10933
		x"45",	--10934
		x"54",	--10935
		x"52",	--10936
		x"47",	--10937
		x"54",	--10938
		x"3c",	--10939
		x"49",	--10940
		x"45",	--10941
		x"55",	--10942
		x"3e",	--10943
		x"0a",	--10944
		x"25",	--10945
		x"20",	--10946
		x"64",	--10947
		x"0a",	--10948
		x"4e",	--10949
		x"74",	--10950
		x"69",	--10951
		x"70",	--10952
		x"65",	--10953
		x"65",	--10954
		x"74",	--10955
		x"64",	--10956
		x"59",	--10957
		x"74",	--10958
		x"0a",	--10959
		x"57",	--10960
		x"69",	--10961
		x"69",	--10962
		x"67",	--10963
		x"66",	--10964
		x"72",	--10965
		x"61",	--10966
		x"6e",	--10967
		x"77",	--10968
		x"2e",	--10969
		x"69",	--10970
		x"20",	--10971
		x"69",	--10972
		x"65",	--10973
		x"0a",	--10974
		x"57",	--10975
		x"20",	--10976
		x"68",	--10977
		x"75",	--10978
		x"64",	--10979
		x"6e",	--10980
		x"74",	--10981
		x"73",	--10982
		x"65",	--10983
		x"74",	--10984
		x"61",	--10985
		x"0d",	--10986
		x"00",	--10987
		x"63",	--10988
		x"69",	--10989
		x"20",	--10990
		x"6f",	--10991
		x"20",	--10992
		x"20",	--10993
		x"75",	--10994
		x"62",	--10995
		x"72",	--10996
		x"0a",	--10997
		x"53",	--10998
		x"6f",	--10999
		x"0d",	--11000
		x"00",	--11001
		x"72",	--11002
		x"6f",	--11003
		x"3a",	--11004
		x"6d",	--11005
		x"73",	--11006
		x"69",	--11007
		x"67",	--11008
		x"61",	--11009
		x"67",	--11010
		x"6d",	--11011
		x"6e",	--11012
		x"0d",	--11013
		x"00",	--11014
		x"6f",	--11015
		x"72",	--11016
		x"63",	--11017
		x"20",	--11018
		x"73",	--11019
		x"67",	--11020
		x"3a",	--11021
		x"0a",	--11022
		x"09",	--11023
		x"73",	--11024
		x"4c",	--11025
		x"46",	--11026
		x"20",	--11027
		x"49",	--11028
		x"48",	--11029
		x"20",	--11030
		x"54",	--11031
		x"4d",	--11032
		x"4f",	--11033
		x"54",	--11034
		x"0d",	--11035
		x"00",	--11036
		x"64",	--11037
		x"25",	--11038
		x"0d",	--11039
		x"00",	--11040
		x"6c",	--11041
		x"20",	--11042
		x"6c",	--11043
		x"00",	--11044
		x"73",	--11045
		x"0a",	--11046
		x"25",	--11047
		x"20",	--11048
		x"64",	--11049
		x"0a",	--11050
		x"00",	--11051
		x"64",	--11052
		x"00",	--11053
		x"0a",	--11054
		x"59",	--11055
		x"20",	--11056
		x"65",	--11057
		x"69",	--11058
		x"64",	--11059
		x"6d",	--11060
		x"0d",	--11061
		x"00",	--11062
		x"6f",	--11063
		x"69",	--11064
		x"20",	--11065
		x"72",	--11066
		x"6e",	--11067
		x"0d",	--11068
		x"00",	--11069
		x"6f",	--11070
		x"6f",	--11071
		x"20",	--11072
		x"68",	--11073
		x"20",	--11074
		x"69",	--11075
		x"68",	--11076
		x"0d",	--11077
		x"00",	--11078
		x"6f",	--11079
		x"6f",	--11080
		x"20",	--11081
		x"68",	--11082
		x"20",	--11083
		x"65",	--11084
		x"74",	--11085
		x"0a",	--11086
		x"25",	--11087
		x"0d",	--11088
		x"00",	--11089
		x"74",	--11090
		x"70",	--11091
		x"0a",	--11092
		x"66",	--11093
		x"6f",	--11094
		x"74",	--11095
		x"72",	--11096
		x"74",	--11097
		x"74",	--11098
		x"6f",	--11099
		x"0d",	--11100
		x"00",	--11101
		x"65",	--11102
		x"74",	--11103
		x"72",	--11104
		x"74",	--11105
		x"74",	--11106
		x"6f",	--11107
		x"0d",	--11108
		x"00",	--11109
		x"69",	--11110
		x"68",	--11111
		x"3a",	--11112
		x"6f",	--11113
		x"61",	--11114
		x"69",	--11115
		x"6e",	--11116
		x"0a",	--11117
		x"52",	--11118
		x"61",	--11119
		x"69",	--11120
		x"67",	--11121
		x"61",	--11122
		x"74",	--11123
		x"76",	--11124
		x"74",	--11125
		x"64",	--11126
		x"0a",	--11127
		x"52",	--11128
		x"61",	--11129
		x"69",	--11130
		x"67",	--11131
		x"64",	--11132
		x"61",	--11133
		x"74",	--11134
		x"76",	--11135
		x"74",	--11136
		x"64",	--11137
		x"0a",	--11138
		x"00",	--11139
		x"01",	--11140
		x"01",	--11141
		x"01",	--11142
		x"01",	--11143
		x"00",	--11144
		x"72",	--11145
		x"74",	--11146
		x"0a",	--11147
		x"00",	--11148
		x"72",	--11149
		x"6f",	--11150
		x"3a",	--11151
		x"6d",	--11152
		x"73",	--11153
		x"69",	--11154
		x"67",	--11155
		x"61",	--11156
		x"67",	--11157
		x"6d",	--11158
		x"6e",	--11159
		x"0d",	--11160
		x"00",	--11161
		x"6f",	--11162
		x"72",	--11163
		x"63",	--11164
		x"20",	--11165
		x"73",	--11166
		x"67",	--11167
		x"3a",	--11168
		x"0a",	--11169
		x"09",	--11170
		x"73",	--11171
		x"52",	--11172
		x"47",	--11173
		x"53",	--11174
		x"45",	--11175
		x"20",	--11176
		x"41",	--11177
		x"55",	--11178
		x"0d",	--11179
		x"00",	--11180
		x"3d",	--11181
		x"64",	--11182
		x"76",	--11183
		x"25",	--11184
		x"0d",	--11185
		x"00",	--11186
		x"25",	--11187
		x"20",	--11188
		x"45",	--11189
		x"49",	--11190
		x"54",	--11191
		x"52",	--11192
		x"0a",	--11193
		x"72",	--11194
		x"61",	--11195
		x"0a",	--11196
		x"00",	--11197
		x"63",	--11198
		x"25",	--11199
		x"0d",	--11200
		x"00",	--11201
		x"63",	--11202
		x"20",	--11203
		x"6f",	--11204
		x"73",	--11205
		x"63",	--11206
		x"20",	--11207
		x"6f",	--11208
		x"6d",	--11209
		x"6e",	--11210
		x"0d",	--11211
		x"00",	--11212
		x"9d",	--11213
		x"9c",	--11214
		x"9c",	--11215
		x"9c",	--11216
		x"9c",	--11217
		x"9c",	--11218
		x"9c",	--11219
		x"9c",	--11220
		x"9c",	--11221
		x"9c",	--11222
		x"9c",	--11223
		x"9c",	--11224
		x"9c",	--11225
		x"9c",	--11226
		x"9c",	--11227
		x"9c",	--11228
		x"9c",	--11229
		x"9c",	--11230
		x"9c",	--11231
		x"9c",	--11232
		x"9c",	--11233
		x"9c",	--11234
		x"9c",	--11235
		x"9c",	--11236
		x"9c",	--11237
		x"9c",	--11238
		x"9c",	--11239
		x"9c",	--11240
		x"9c",	--11241
		x"9d",	--11242
		x"9c",	--11243
		x"9c",	--11244
		x"9c",	--11245
		x"9c",	--11246
		x"9c",	--11247
		x"9c",	--11248
		x"9c",	--11249
		x"9c",	--11250
		x"9c",	--11251
		x"9c",	--11252
		x"9c",	--11253
		x"9c",	--11254
		x"9c",	--11255
		x"9c",	--11256
		x"9c",	--11257
		x"9c",	--11258
		x"9c",	--11259
		x"9c",	--11260
		x"9c",	--11261
		x"9c",	--11262
		x"9c",	--11263
		x"9c",	--11264
		x"9c",	--11265
		x"9c",	--11266
		x"9c",	--11267
		x"9c",	--11268
		x"9c",	--11269
		x"9c",	--11270
		x"9c",	--11271
		x"9c",	--11272
		x"9c",	--11273
		x"9d",	--11274
		x"9c",	--11275
		x"9c",	--11276
		x"9c",	--11277
		x"9c",	--11278
		x"9c",	--11279
		x"9c",	--11280
		x"9c",	--11281
		x"9c",	--11282
		x"9c",	--11283
		x"9c",	--11284
		x"9c",	--11285
		x"9c",	--11286
		x"9c",	--11287
		x"9c",	--11288
		x"9c",	--11289
		x"9c",	--11290
		x"9c",	--11291
		x"9c",	--11292
		x"9c",	--11293
		x"9c",	--11294
		x"9c",	--11295
		x"9c",	--11296
		x"31",	--11297
		x"33",	--11298
		x"35",	--11299
		x"37",	--11300
		x"39",	--11301
		x"62",	--11302
		x"64",	--11303
		x"66",	--11304
		x"00",	--11305
		x"63",	--11306
		x"3e",	--11307
		x"0f",	--11308
		x"3f",	--11309
		x"98",	--11310
		x"3f",	--11311
		x"0f",	--11312
		x"3f",	--11313
		x"37",	--11314
		x"31",	--11315
		x"21",	--11316
		x"33",	--11317
		x"0f",	--11318
		x"33",	--11319
		x"21",	--11320
		x"33",	--11321
		x"0f",	--11322
		x"3f",	--11323
		x"0f",	--11324
		x"40",	--11325
		x"cb",	--11326
		x"40",	--11327
		x"0f",	--11328
		x"40",	--11329
		x"53",	--11330
		x"40",	--11331
		x"cb",	--11332
		x"41",	--11333
		x"ed",	--11334
		x"41",	--11335
		x"0f",	--11336
		x"41",	--11337
		x"31",	--11338
		x"41",	--11339
		x"53",	--11340
		x"41",	--11341
		x"3a",	--11342
		x"41",	--11343
		x"cb",	--11344
		x"41",	--11345
		x"5c",	--11346
		x"41",	--11347
		x"ed",	--11348
		x"41",	--11349
		x"7e",	--11350
		x"41",	--11351
		x"0f",	--11352
		x"41",	--11353
		x"a0",	--11354
		x"41",	--11355
		x"31",	--11356
		x"41",	--11357
		x"c2",	--11358
		x"41",	--11359
		x"53",	--11360
		x"41",	--11361
		x"f2",	--11362
		x"42",	--11363
		x"3a",	--11364
		x"42",	--11365
		x"83",	--11366
		x"42",	--11367
		x"cb",	--11368
		x"42",	--11369
		x"14",	--11370
		x"42",	--11371
		x"5c",	--11372
		x"42",	--11373
		x"a5",	--11374
		x"42",	--11375
		x"ed",	--11376
		x"42",	--11377
		x"36",	--11378
		x"42",	--11379
		x"7e",	--11380
		x"42",	--11381
		x"c7",	--11382
		x"42",	--11383
		x"0f",	--11384
		x"42",	--11385
		x"00",	--11386
		x"00",	--11387
		x"00",	--11388
		x"00",	--11389
		x"00",	--11390
		x"00",	--11391
		x"00",	--11392
		x"00",	--11393
		x"00",	--11394
		x"00",	--11395
		x"00",	--11396
		x"00",	--11397
		x"00",	--11398
		x"00",	--11399
		x"00",	--11400
		x"00",	--11401
		x"00",	--11402
		x"00",	--11403
		x"00",	--11404
		x"00",	--11405
		x"00",	--11406
		x"00",	--11407
		x"00",	--11408
		x"00",	--11409
		x"00",	--11410
		x"00",	--11411
		x"00",	--11412
		x"00",	--11413
		x"00",	--11414
		x"00",	--11415
		x"00",	--11416
		x"00",	--11417
		x"00",	--11418
		x"00",	--11419
		x"00",	--11420
		x"00",	--11421
		x"00",	--11422
		x"00",	--11423
		x"00",	--11424
		x"00",	--11425
		x"00",	--11426
		x"00",	--11427
		x"00",	--11428
		x"00",	--11429
		x"00",	--11430
		x"00",	--11431
		x"00",	--11432
		x"00",	--11433
		x"00",	--11434
		x"00",	--11435
		x"00",	--11436
		x"00",	--11437
		x"00",	--11438
		x"00",	--11439
		x"00",	--11440
		x"00",	--11441
		x"00",	--11442
		x"00",	--11443
		x"00",	--11444
		x"00",	--11445
		x"00",	--11446
		x"00",	--11447
		x"00",	--11448
		x"00",	--11449
		x"00",	--11450
		x"00",	--11451
		x"00",	--11452
		x"00",	--11453
		x"00",	--11454
		x"00",	--11455
		x"00",	--11456
		x"00",	--11457
		x"00",	--11458
		x"00",	--11459
		x"00",	--11460
		x"00",	--11461
		x"00",	--11462
		x"00",	--11463
		x"00",	--11464
		x"00",	--11465
		x"00",	--11466
		x"00",	--11467
		x"00",	--11468
		x"00",	--11469
		x"00",	--11470
		x"00",	--11471
		x"00",	--11472
		x"00",	--11473
		x"00",	--11474
		x"00",	--11475
		x"00",	--11476
		x"00",	--11477
		x"00",	--11478
		x"00",	--11479
		x"00",	--11480
		x"00",	--11481
		x"00",	--11482
		x"00",	--11483
		x"00",	--11484
		x"00",	--11485
		x"00",	--11486
		x"00",	--11487
		x"00",	--11488
		x"00",	--11489
		x"00",	--11490
		x"00",	--11491
		x"00",	--11492
		x"00",	--11493
		x"00",	--11494
		x"00",	--11495
		x"00",	--11496
		x"00",	--11497
		x"00",	--11498
		x"00",	--11499
		x"00",	--11500
		x"00",	--11501
		x"00",	--11502
		x"00",	--11503
		x"00",	--11504
		x"00",	--11505
		x"00",	--11506
		x"00",	--11507
		x"00",	--11508
		x"00",	--11509
		x"00",	--11510
		x"00",	--11511
		x"00",	--11512
		x"00",	--11513
		x"00",	--11514
		x"00",	--11515
		x"00",	--11516
		x"00",	--11517
		x"00",	--11518
		x"00",	--11519
		x"00",	--11520
		x"00",	--11521
		x"00",	--11522
		x"00",	--11523
		x"00",	--11524
		x"00",	--11525
		x"00",	--11526
		x"00",	--11527
		x"00",	--11528
		x"00",	--11529
		x"00",	--11530
		x"00",	--11531
		x"00",	--11532
		x"00",	--11533
		x"00",	--11534
		x"00",	--11535
		x"00",	--11536
		x"00",	--11537
		x"00",	--11538
		x"00",	--11539
		x"00",	--11540
		x"00",	--11541
		x"00",	--11542
		x"00",	--11543
		x"00",	--11544
		x"00",	--11545
		x"00",	--11546
		x"00",	--11547
		x"00",	--11548
		x"00",	--11549
		x"00",	--11550
		x"00",	--11551
		x"00",	--11552
		x"00",	--11553
		x"00",	--11554
		x"00",	--11555
		x"00",	--11556
		x"00",	--11557
		x"00",	--11558
		x"00",	--11559
		x"00",	--11560
		x"00",	--11561
		x"00",	--11562
		x"00",	--11563
		x"00",	--11564
		x"00",	--11565
		x"00",	--11566
		x"00",	--11567
		x"00",	--11568
		x"00",	--11569
		x"00",	--11570
		x"00",	--11571
		x"00",	--11572
		x"00",	--11573
		x"00",	--11574
		x"00",	--11575
		x"00",	--11576
		x"00",	--11577
		x"00",	--11578
		x"00",	--11579
		x"00",	--11580
		x"00",	--11581
		x"00",	--11582
		x"00",	--11583
		x"00",	--11584
		x"00",	--11585
		x"00",	--11586
		x"00",	--11587
		x"00",	--11588
		x"00",	--11589
		x"00",	--11590
		x"00",	--11591
		x"00",	--11592
		x"00",	--11593
		x"00",	--11594
		x"00",	--11595
		x"00",	--11596
		x"00",	--11597
		x"00",	--11598
		x"00",	--11599
		x"00",	--11600
		x"00",	--11601
		x"00",	--11602
		x"00",	--11603
		x"00",	--11604
		x"00",	--11605
		x"00",	--11606
		x"00",	--11607
		x"00",	--11608
		x"00",	--11609
		x"00",	--11610
		x"00",	--11611
		x"00",	--11612
		x"00",	--11613
		x"00",	--11614
		x"00",	--11615
		x"00",	--11616
		x"00",	--11617
		x"00",	--11618
		x"00",	--11619
		x"00",	--11620
		x"00",	--11621
		x"00",	--11622
		x"00",	--11623
		x"00",	--11624
		x"00",	--11625
		x"00",	--11626
		x"00",	--11627
		x"00",	--11628
		x"00",	--11629
		x"00",	--11630
		x"00",	--11631
		x"00",	--11632
		x"00",	--11633
		x"00",	--11634
		x"00",	--11635
		x"00",	--11636
		x"00",	--11637
		x"00",	--11638
		x"00",	--11639
		x"00",	--11640
		x"00",	--11641
		x"00",	--11642
		x"00",	--11643
		x"00",	--11644
		x"00",	--11645
		x"00",	--11646
		x"00",	--11647
		x"00",	--11648
		x"00",	--11649
		x"00",	--11650
		x"00",	--11651
		x"00",	--11652
		x"00",	--11653
		x"00",	--11654
		x"00",	--11655
		x"00",	--11656
		x"00",	--11657
		x"00",	--11658
		x"00",	--11659
		x"00",	--11660
		x"00",	--11661
		x"00",	--11662
		x"00",	--11663
		x"00",	--11664
		x"00",	--11665
		x"00",	--11666
		x"00",	--11667
		x"00",	--11668
		x"00",	--11669
		x"00",	--11670
		x"00",	--11671
		x"00",	--11672
		x"00",	--11673
		x"00",	--11674
		x"00",	--11675
		x"00",	--11676
		x"00",	--11677
		x"00",	--11678
		x"00",	--11679
		x"00",	--11680
		x"00",	--11681
		x"00",	--11682
		x"00",	--11683
		x"00",	--11684
		x"00",	--11685
		x"00",	--11686
		x"00",	--11687
		x"00",	--11688
		x"00",	--11689
		x"00",	--11690
		x"00",	--11691
		x"00",	--11692
		x"00",	--11693
		x"00",	--11694
		x"00",	--11695
		x"00",	--11696
		x"00",	--11697
		x"00",	--11698
		x"00",	--11699
		x"00",	--11700
		x"00",	--11701
		x"00",	--11702
		x"00",	--11703
		x"00",	--11704
		x"00",	--11705
		x"00",	--11706
		x"00",	--11707
		x"00",	--11708
		x"00",	--11709
		x"00",	--11710
		x"00",	--11711
		x"00",	--11712
		x"00",	--11713
		x"00",	--11714
		x"00",	--11715
		x"00",	--11716
		x"00",	--11717
		x"00",	--11718
		x"00",	--11719
		x"00",	--11720
		x"00",	--11721
		x"00",	--11722
		x"00",	--11723
		x"00",	--11724
		x"00",	--11725
		x"00",	--11726
		x"00",	--11727
		x"00",	--11728
		x"00",	--11729
		x"00",	--11730
		x"00",	--11731
		x"00",	--11732
		x"00",	--11733
		x"00",	--11734
		x"00",	--11735
		x"00",	--11736
		x"00",	--11737
		x"00",	--11738
		x"00",	--11739
		x"00",	--11740
		x"00",	--11741
		x"00",	--11742
		x"00",	--11743
		x"00",	--11744
		x"00",	--11745
		x"00",	--11746
		x"00",	--11747
		x"00",	--11748
		x"00",	--11749
		x"00",	--11750
		x"00",	--11751
		x"00",	--11752
		x"00",	--11753
		x"00",	--11754
		x"00",	--11755
		x"00",	--11756
		x"00",	--11757
		x"00",	--11758
		x"00",	--11759
		x"00",	--11760
		x"00",	--11761
		x"00",	--11762
		x"00",	--11763
		x"00",	--11764
		x"00",	--11765
		x"00",	--11766
		x"00",	--11767
		x"00",	--11768
		x"00",	--11769
		x"00",	--11770
		x"00",	--11771
		x"00",	--11772
		x"00",	--11773
		x"00",	--11774
		x"00",	--11775
		x"00",	--11776
		x"00",	--11777
		x"00",	--11778
		x"00",	--11779
		x"00",	--11780
		x"00",	--11781
		x"00",	--11782
		x"00",	--11783
		x"00",	--11784
		x"00",	--11785
		x"3f",	--11786
		x"00",	--11787
		x"39",	--11788
		x"00",	--11789
		x"37",	--11790
		x"00",	--11791
		x"33",	--11792
		x"00",	--11793
		x"2e",	--11794
		x"00",	--11795
		x"2b",	--11796
		x"00",	--11797
		x"27",	--11798
		x"00",	--11799
		x"22",	--11800
		x"00",	--11801
		x"1f",	--11802
		x"00",	--11803
		x"1b",	--11804
		x"00",	--11805
		x"17",	--11806
		x"00",	--11807
		x"00",	--11808
		x"00",	--11809
		x"00",	--11810
		x"01",	--11811
		x"02",	--11812
		x"03",	--11813
		x"03",	--11814
		x"04",	--11815
		x"04",	--11816
		x"04",	--11817
		x"04",	--11818
		x"05",	--11819
		x"05",	--11820
		x"05",	--11821
		x"05",	--11822
		x"05",	--11823
		x"05",	--11824
		x"05",	--11825
		x"05",	--11826
		x"06",	--11827
		x"06",	--11828
		x"06",	--11829
		x"06",	--11830
		x"06",	--11831
		x"06",	--11832
		x"06",	--11833
		x"06",	--11834
		x"06",	--11835
		x"06",	--11836
		x"06",	--11837
		x"06",	--11838
		x"06",	--11839
		x"06",	--11840
		x"06",	--11841
		x"06",	--11842
		x"07",	--11843
		x"07",	--11844
		x"07",	--11845
		x"07",	--11846
		x"07",	--11847
		x"07",	--11848
		x"07",	--11849
		x"07",	--11850
		x"07",	--11851
		x"07",	--11852
		x"07",	--11853
		x"07",	--11854
		x"07",	--11855
		x"07",	--11856
		x"07",	--11857
		x"07",	--11858
		x"07",	--11859
		x"07",	--11860
		x"07",	--11861
		x"07",	--11862
		x"07",	--11863
		x"07",	--11864
		x"07",	--11865
		x"07",	--11866
		x"07",	--11867
		x"07",	--11868
		x"07",	--11869
		x"07",	--11870
		x"07",	--11871
		x"07",	--11872
		x"07",	--11873
		x"07",	--11874
		x"08",	--11875
		x"08",	--11876
		x"08",	--11877
		x"08",	--11878
		x"08",	--11879
		x"08",	--11880
		x"08",	--11881
		x"08",	--11882
		x"08",	--11883
		x"08",	--11884
		x"08",	--11885
		x"08",	--11886
		x"08",	--11887
		x"08",	--11888
		x"08",	--11889
		x"08",	--11890
		x"08",	--11891
		x"08",	--11892
		x"08",	--11893
		x"08",	--11894
		x"08",	--11895
		x"08",	--11896
		x"08",	--11897
		x"08",	--11898
		x"08",	--11899
		x"08",	--11900
		x"08",	--11901
		x"08",	--11902
		x"08",	--11903
		x"08",	--11904
		x"08",	--11905
		x"08",	--11906
		x"08",	--11907
		x"08",	--11908
		x"08",	--11909
		x"08",	--11910
		x"08",	--11911
		x"08",	--11912
		x"08",	--11913
		x"08",	--11914
		x"08",	--11915
		x"08",	--11916
		x"08",	--11917
		x"08",	--11918
		x"08",	--11919
		x"08",	--11920
		x"08",	--11921
		x"08",	--11922
		x"08",	--11923
		x"08",	--11924
		x"08",	--11925
		x"08",	--11926
		x"08",	--11927
		x"08",	--11928
		x"08",	--11929
		x"08",	--11930
		x"08",	--11931
		x"08",	--11932
		x"08",	--11933
		x"08",	--11934
		x"08",	--11935
		x"08",	--11936
		x"08",	--11937
		x"08",	--11938
		x"6e",	--11939
		x"6c",	--11940
		x"29",	--11941
		x"00",	--11942
		x"ff",	--11943
		x"ff",	--11944
		x"ff",	--11945
		x"ff",	--11946
		x"65",	--11947
		x"70",	--11948
		x"00",	--11949
		x"ff",	--11950
		x"ff",	--11951
		x"ff",	--11952
		x"ff",	--11953
		x"ff",	--11954
		x"ff",	--11955
		x"ff",	--11956
		x"ff",	--11957
		x"ff",	--11958
		x"ff",	--11959
		x"ff",	--11960
		x"ff",	--11961
		x"ff",	--11962
		x"ff",	--11963
		x"ff",	--11964
		x"ff",	--11965
		x"ff",	--11966
		x"ff",	--11967
		x"ff",	--11968
		x"ff",	--11969
		x"ff",	--11970
		x"ff",	--11971
		x"ff",	--11972
		x"ff",	--11973
		x"ff",	--11974
		x"ff",	--11975
		x"ff",	--11976
		x"ff",	--11977
		x"ff",	--11978
		x"ff",	--11979
		x"ff",	--11980
		x"ff",	--11981
		x"ff",	--11982
		x"ff",	--11983
		x"ff",	--11984
		x"ff",	--11985
		x"ff",	--11986
		x"ff",	--11987
		x"ff",	--11988
		x"ff",	--11989
		x"ff",	--11990
		x"ff",	--11991
		x"ff",	--11992
		x"ff",	--11993
		x"ff",	--11994
		x"ff",	--11995
		x"ff",	--11996
		x"ff",	--11997
		x"ff",	--11998
		x"ff",	--11999
		x"ff",	--12000
		x"ff",	--12001
		x"ff",	--12002
		x"ff",	--12003
		x"ff",	--12004
		x"ff",	--12005
		x"ff",	--12006
		x"ff",	--12007
		x"ff",	--12008
		x"ff",	--12009
		x"ff",	--12010
		x"ff",	--12011
		x"ff",	--12012
		x"ff",	--12013
		x"ff",	--12014
		x"ff",	--12015
		x"ff",	--12016
		x"ff",	--12017
		x"ff",	--12018
		x"ff",	--12019
		x"ff",	--12020
		x"ff",	--12021
		x"ff",	--12022
		x"ff",	--12023
		x"ff",	--12024
		x"ff",	--12025
		x"ff",	--12026
		x"ff",	--12027
		x"ff",	--12028
		x"ff",	--12029
		x"ff",	--12030
		x"ff",	--12031
		x"ff",	--12032
		x"ff",	--12033
		x"ff",	--12034
		x"ff",	--12035
		x"ff",	--12036
		x"ff",	--12037
		x"ff",	--12038
		x"ff",	--12039
		x"ff",	--12040
		x"ff",	--12041
		x"ff",	--12042
		x"ff",	--12043
		x"ff",	--12044
		x"ff",	--12045
		x"ff",	--12046
		x"ff",	--12047
		x"ff",	--12048
		x"ff",	--12049
		x"ff",	--12050
		x"ff",	--12051
		x"ff",	--12052
		x"ff",	--12053
		x"ff",	--12054
		x"ff",	--12055
		x"ff",	--12056
		x"ff",	--12057
		x"ff",	--12058
		x"ff",	--12059
		x"ff",	--12060
		x"ff",	--12061
		x"ff",	--12062
		x"ff",	--12063
		x"ff",	--12064
		x"ff",	--12065
		x"ff",	--12066
		x"ff",	--12067
		x"ff",	--12068
		x"ff",	--12069
		x"ff",	--12070
		x"ff",	--12071
		x"ff",	--12072
		x"ff",	--12073
		x"ff",	--12074
		x"ff",	--12075
		x"ff",	--12076
		x"ff",	--12077
		x"ff",	--12078
		x"ff",	--12079
		x"ff",	--12080
		x"ff",	--12081
		x"ff",	--12082
		x"ff",	--12083
		x"ff",	--12084
		x"ff",	--12085
		x"ff",	--12086
		x"ff",	--12087
		x"ff",	--12088
		x"ff",	--12089
		x"ff",	--12090
		x"ff",	--12091
		x"ff",	--12092
		x"ff",	--12093
		x"ff",	--12094
		x"ff",	--12095
		x"ff",	--12096
		x"ff",	--12097
		x"ff",	--12098
		x"ff",	--12099
		x"ff",	--12100
		x"ff",	--12101
		x"ff",	--12102
		x"ff",	--12103
		x"ff",	--12104
		x"ff",	--12105
		x"ff",	--12106
		x"ff",	--12107
		x"ff",	--12108
		x"ff",	--12109
		x"ff",	--12110
		x"ff",	--12111
		x"ff",	--12112
		x"ff",	--12113
		x"ff",	--12114
		x"ff",	--12115
		x"ff",	--12116
		x"ff",	--12117
		x"ff",	--12118
		x"ff",	--12119
		x"ff",	--12120
		x"ff",	--12121
		x"ff",	--12122
		x"ff",	--12123
		x"ff",	--12124
		x"ff",	--12125
		x"ff",	--12126
		x"ff",	--12127
		x"ff",	--12128
		x"ff",	--12129
		x"ff",	--12130
		x"ff",	--12131
		x"ff",	--12132
		x"ff",	--12133
		x"ff",	--12134
		x"ff",	--12135
		x"ff",	--12136
		x"ff",	--12137
		x"ff",	--12138
		x"ff",	--12139
		x"ff",	--12140
		x"ff",	--12141
		x"ff",	--12142
		x"ff",	--12143
		x"ff",	--12144
		x"ff",	--12145
		x"ff",	--12146
		x"ff",	--12147
		x"ff",	--12148
		x"ff",	--12149
		x"ff",	--12150
		x"ff",	--12151
		x"ff",	--12152
		x"ff",	--12153
		x"ff",	--12154
		x"ff",	--12155
		x"ff",	--12156
		x"ff",	--12157
		x"ff",	--12158
		x"ff",	--12159
		x"ff",	--12160
		x"ff",	--12161
		x"ff",	--12162
		x"ff",	--12163
		x"ff",	--12164
		x"ff",	--12165
		x"ff",	--12166
		x"ff",	--12167
		x"ff",	--12168
		x"ff",	--12169
		x"ff",	--12170
		x"ff",	--12171
		x"ff",	--12172
		x"ff",	--12173
		x"ff",	--12174
		x"ff",	--12175
		x"ff",	--12176
		x"ff",	--12177
		x"ff",	--12178
		x"ff",	--12179
		x"ff",	--12180
		x"ff",	--12181
		x"ff",	--12182
		x"ff",	--12183
		x"ff",	--12184
		x"ff",	--12185
		x"ff",	--12186
		x"ff",	--12187
		x"ff",	--12188
		x"ff",	--12189
		x"ff",	--12190
		x"ff",	--12191
		x"ff",	--12192
		x"ff",	--12193
		x"ff",	--12194
		x"ff",	--12195
		x"ff",	--12196
		x"ff",	--12197
		x"ff",	--12198
		x"ff",	--12199
		x"ff",	--12200
		x"ff",	--12201
		x"ff",	--12202
		x"ff",	--12203
		x"ff",	--12204
		x"ff",	--12205
		x"ff",	--12206
		x"ff",	--12207
		x"ff",	--12208
		x"ff",	--12209
		x"ff",	--12210
		x"ff",	--12211
		x"ff",	--12212
		x"ff",	--12213
		x"ff",	--12214
		x"ff",	--12215
		x"ff",	--12216
		x"ff",	--12217
		x"ff",	--12218
		x"ff",	--12219
		x"ff",	--12220
		x"ff",	--12221
		x"ff",	--12222
		x"ff",	--12223
		x"ff",	--12224
		x"ff",	--12225
		x"ff",	--12226
		x"ff",	--12227
		x"ff",	--12228
		x"ff",	--12229
		x"ff",	--12230
		x"ff",	--12231
		x"ff",	--12232
		x"ff",	--12233
		x"ff",	--12234
		x"ff",	--12235
		x"ff",	--12236
		x"ff",	--12237
		x"ff",	--12238
		x"ff",	--12239
		x"ff",	--12240
		x"ff",	--12241
		x"ff",	--12242
		x"ff",	--12243
		x"ff",	--12244
		x"ff",	--12245
		x"ff",	--12246
		x"ff",	--12247
		x"ff",	--12248
		x"ff",	--12249
		x"ff",	--12250
		x"ff",	--12251
		x"ff",	--12252
		x"ff",	--12253
		x"ff",	--12254
		x"ff",	--12255
		x"ff",	--12256
		x"ff",	--12257
		x"ff",	--12258
		x"ff",	--12259
		x"ff",	--12260
		x"ff",	--12261
		x"ff",	--12262
		x"ff",	--12263
		x"ff",	--12264
		x"ff",	--12265
		x"ff",	--12266
		x"ff",	--12267
		x"ff",	--12268
		x"ff",	--12269
		x"ff",	--12270
		x"ff",	--12271
		x"ff",	--12272
		x"ff",	--12273
		x"ff",	--12274
		x"ff",	--12275
		x"ff",	--12276
		x"ff",	--12277
		x"ff",	--12278
		x"ff",	--12279
		x"ff",	--12280
		x"ff",	--12281
		x"ff",	--12282
		x"ff",	--12283
		x"ff",	--12284
		x"ff",	--12285
		x"ff",	--12286
		x"ff",	--12287
		x"ff",	--12288
		x"ff",	--12289
		x"ff",	--12290
		x"ff",	--12291
		x"ff",	--12292
		x"ff",	--12293
		x"ff",	--12294
		x"ff",	--12295
		x"ff",	--12296
		x"ff",	--12297
		x"ff",	--12298
		x"ff",	--12299
		x"ff",	--12300
		x"ff",	--12301
		x"ff",	--12302
		x"ff",	--12303
		x"ff",	--12304
		x"ff",	--12305
		x"ff",	--12306
		x"ff",	--12307
		x"ff",	--12308
		x"ff",	--12309
		x"ff",	--12310
		x"ff",	--12311
		x"ff",	--12312
		x"ff",	--12313
		x"ff",	--12314
		x"ff",	--12315
		x"ff",	--12316
		x"ff",	--12317
		x"ff",	--12318
		x"ff",	--12319
		x"ff",	--12320
		x"ff",	--12321
		x"ff",	--12322
		x"ff",	--12323
		x"ff",	--12324
		x"ff",	--12325
		x"ff",	--12326
		x"ff",	--12327
		x"ff",	--12328
		x"ff",	--12329
		x"ff",	--12330
		x"ff",	--12331
		x"ff",	--12332
		x"ff",	--12333
		x"ff",	--12334
		x"ff",	--12335
		x"ff",	--12336
		x"ff",	--12337
		x"ff",	--12338
		x"ff",	--12339
		x"ff",	--12340
		x"ff",	--12341
		x"ff",	--12342
		x"ff",	--12343
		x"ff",	--12344
		x"ff",	--12345
		x"ff",	--12346
		x"ff",	--12347
		x"ff",	--12348
		x"ff",	--12349
		x"ff",	--12350
		x"ff",	--12351
		x"ff",	--12352
		x"ff",	--12353
		x"ff",	--12354
		x"ff",	--12355
		x"ff",	--12356
		x"ff",	--12357
		x"ff",	--12358
		x"ff",	--12359
		x"ff",	--12360
		x"ff",	--12361
		x"ff",	--12362
		x"ff",	--12363
		x"ff",	--12364
		x"ff",	--12365
		x"ff",	--12366
		x"ff",	--12367
		x"ff",	--12368
		x"ff",	--12369
		x"ff",	--12370
		x"ff",	--12371
		x"ff",	--12372
		x"ff",	--12373
		x"ff",	--12374
		x"ff",	--12375
		x"ff",	--12376
		x"ff",	--12377
		x"ff",	--12378
		x"ff",	--12379
		x"ff",	--12380
		x"ff",	--12381
		x"ff",	--12382
		x"ff",	--12383
		x"ff",	--12384
		x"ff",	--12385
		x"ff",	--12386
		x"ff",	--12387
		x"ff",	--12388
		x"ff",	--12389
		x"ff",	--12390
		x"ff",	--12391
		x"ff",	--12392
		x"ff",	--12393
		x"ff",	--12394
		x"ff",	--12395
		x"ff",	--12396
		x"ff",	--12397
		x"ff",	--12398
		x"ff",	--12399
		x"ff",	--12400
		x"ff",	--12401
		x"ff",	--12402
		x"ff",	--12403
		x"ff",	--12404
		x"ff",	--12405
		x"ff",	--12406
		x"ff",	--12407
		x"ff",	--12408
		x"ff",	--12409
		x"ff",	--12410
		x"ff",	--12411
		x"ff",	--12412
		x"ff",	--12413
		x"ff",	--12414
		x"ff",	--12415
		x"ff",	--12416
		x"ff",	--12417
		x"ff",	--12418
		x"ff",	--12419
		x"ff",	--12420
		x"ff",	--12421
		x"ff",	--12422
		x"ff",	--12423
		x"ff",	--12424
		x"ff",	--12425
		x"ff",	--12426
		x"ff",	--12427
		x"ff",	--12428
		x"ff",	--12429
		x"ff",	--12430
		x"ff",	--12431
		x"ff",	--12432
		x"ff",	--12433
		x"ff",	--12434
		x"ff",	--12435
		x"ff",	--12436
		x"ff",	--12437
		x"ff",	--12438
		x"ff",	--12439
		x"ff",	--12440
		x"ff",	--12441
		x"ff",	--12442
		x"ff",	--12443
		x"ff",	--12444
		x"ff",	--12445
		x"ff",	--12446
		x"ff",	--12447
		x"ff",	--12448
		x"ff",	--12449
		x"ff",	--12450
		x"ff",	--12451
		x"ff",	--12452
		x"ff",	--12453
		x"ff",	--12454
		x"ff",	--12455
		x"ff",	--12456
		x"ff",	--12457
		x"ff",	--12458
		x"ff",	--12459
		x"ff",	--12460
		x"ff",	--12461
		x"ff",	--12462
		x"ff",	--12463
		x"ff",	--12464
		x"ff",	--12465
		x"ff",	--12466
		x"ff",	--12467
		x"ff",	--12468
		x"ff",	--12469
		x"ff",	--12470
		x"ff",	--12471
		x"ff",	--12472
		x"ff",	--12473
		x"ff",	--12474
		x"ff",	--12475
		x"ff",	--12476
		x"ff",	--12477
		x"ff",	--12478
		x"ff",	--12479
		x"ff",	--12480
		x"ff",	--12481
		x"ff",	--12482
		x"ff",	--12483
		x"ff",	--12484
		x"ff",	--12485
		x"ff",	--12486
		x"ff",	--12487
		x"ff",	--12488
		x"ff",	--12489
		x"ff",	--12490
		x"ff",	--12491
		x"ff",	--12492
		x"ff",	--12493
		x"ff",	--12494
		x"ff",	--12495
		x"ff",	--12496
		x"ff",	--12497
		x"ff",	--12498
		x"ff",	--12499
		x"ff",	--12500
		x"ff",	--12501
		x"ff",	--12502
		x"ff",	--12503
		x"ff",	--12504
		x"ff",	--12505
		x"ff",	--12506
		x"ff",	--12507
		x"ff",	--12508
		x"ff",	--12509
		x"ff",	--12510
		x"ff",	--12511
		x"ff",	--12512
		x"ff",	--12513
		x"ff",	--12514
		x"ff",	--12515
		x"ff",	--12516
		x"ff",	--12517
		x"ff",	--12518
		x"ff",	--12519
		x"ff",	--12520
		x"ff",	--12521
		x"ff",	--12522
		x"ff",	--12523
		x"ff",	--12524
		x"ff",	--12525
		x"ff",	--12526
		x"ff",	--12527
		x"ff",	--12528
		x"ff",	--12529
		x"ff",	--12530
		x"ff",	--12531
		x"ff",	--12532
		x"ff",	--12533
		x"ff",	--12534
		x"ff",	--12535
		x"ff",	--12536
		x"ff",	--12537
		x"ff",	--12538
		x"ff",	--12539
		x"ff",	--12540
		x"ff",	--12541
		x"ff",	--12542
		x"ff",	--12543
		x"ff",	--12544
		x"ff",	--12545
		x"ff",	--12546
		x"ff",	--12547
		x"ff",	--12548
		x"ff",	--12549
		x"ff",	--12550
		x"ff",	--12551
		x"ff",	--12552
		x"ff",	--12553
		x"ff",	--12554
		x"ff",	--12555
		x"ff",	--12556
		x"ff",	--12557
		x"ff",	--12558
		x"ff",	--12559
		x"ff",	--12560
		x"ff",	--12561
		x"ff",	--12562
		x"ff",	--12563
		x"ff",	--12564
		x"ff",	--12565
		x"ff",	--12566
		x"ff",	--12567
		x"ff",	--12568
		x"ff",	--12569
		x"ff",	--12570
		x"ff",	--12571
		x"ff",	--12572
		x"ff",	--12573
		x"ff",	--12574
		x"ff",	--12575
		x"ff",	--12576
		x"ff",	--12577
		x"ff",	--12578
		x"ff",	--12579
		x"ff",	--12580
		x"ff",	--12581
		x"ff",	--12582
		x"ff",	--12583
		x"ff",	--12584
		x"ff",	--12585
		x"ff",	--12586
		x"ff",	--12587
		x"ff",	--12588
		x"ff",	--12589
		x"ff",	--12590
		x"ff",	--12591
		x"ff",	--12592
		x"ff",	--12593
		x"ff",	--12594
		x"ff",	--12595
		x"ff",	--12596
		x"ff",	--12597
		x"ff",	--12598
		x"ff",	--12599
		x"ff",	--12600
		x"ff",	--12601
		x"ff",	--12602
		x"ff",	--12603
		x"ff",	--12604
		x"ff",	--12605
		x"ff",	--12606
		x"ff",	--12607
		x"ff",	--12608
		x"ff",	--12609
		x"ff",	--12610
		x"ff",	--12611
		x"ff",	--12612
		x"ff",	--12613
		x"ff",	--12614
		x"ff",	--12615
		x"ff",	--12616
		x"ff",	--12617
		x"ff",	--12618
		x"ff",	--12619
		x"ff",	--12620
		x"ff",	--12621
		x"ff",	--12622
		x"ff",	--12623
		x"ff",	--12624
		x"ff",	--12625
		x"ff",	--12626
		x"ff",	--12627
		x"ff",	--12628
		x"ff",	--12629
		x"ff",	--12630
		x"ff",	--12631
		x"ff",	--12632
		x"ff",	--12633
		x"ff",	--12634
		x"ff",	--12635
		x"ff",	--12636
		x"ff",	--12637
		x"ff",	--12638
		x"ff",	--12639
		x"ff",	--12640
		x"ff",	--12641
		x"ff",	--12642
		x"ff",	--12643
		x"ff",	--12644
		x"ff",	--12645
		x"ff",	--12646
		x"ff",	--12647
		x"ff",	--12648
		x"ff",	--12649
		x"ff",	--12650
		x"ff",	--12651
		x"ff",	--12652
		x"ff",	--12653
		x"ff",	--12654
		x"ff",	--12655
		x"ff",	--12656
		x"ff",	--12657
		x"ff",	--12658
		x"ff",	--12659
		x"ff",	--12660
		x"ff",	--12661
		x"ff",	--12662
		x"ff",	--12663
		x"ff",	--12664
		x"ff",	--12665
		x"ff",	--12666
		x"ff",	--12667
		x"ff",	--12668
		x"ff",	--12669
		x"ff",	--12670
		x"ff",	--12671
		x"ff",	--12672
		x"ff",	--12673
		x"ff",	--12674
		x"ff",	--12675
		x"ff",	--12676
		x"ff",	--12677
		x"ff",	--12678
		x"ff",	--12679
		x"ff",	--12680
		x"ff",	--12681
		x"ff",	--12682
		x"ff",	--12683
		x"ff",	--12684
		x"ff",	--12685
		x"ff",	--12686
		x"ff",	--12687
		x"ff",	--12688
		x"ff",	--12689
		x"ff",	--12690
		x"ff",	--12691
		x"ff",	--12692
		x"ff",	--12693
		x"ff",	--12694
		x"ff",	--12695
		x"ff",	--12696
		x"ff",	--12697
		x"ff",	--12698
		x"ff",	--12699
		x"ff",	--12700
		x"ff",	--12701
		x"ff",	--12702
		x"ff",	--12703
		x"ff",	--12704
		x"ff",	--12705
		x"ff",	--12706
		x"ff",	--12707
		x"ff",	--12708
		x"ff",	--12709
		x"ff",	--12710
		x"ff",	--12711
		x"ff",	--12712
		x"ff",	--12713
		x"ff",	--12714
		x"ff",	--12715
		x"ff",	--12716
		x"ff",	--12717
		x"ff",	--12718
		x"ff",	--12719
		x"ff",	--12720
		x"ff",	--12721
		x"ff",	--12722
		x"ff",	--12723
		x"ff",	--12724
		x"ff",	--12725
		x"ff",	--12726
		x"ff",	--12727
		x"ff",	--12728
		x"ff",	--12729
		x"ff",	--12730
		x"ff",	--12731
		x"ff",	--12732
		x"ff",	--12733
		x"ff",	--12734
		x"ff",	--12735
		x"ff",	--12736
		x"ff",	--12737
		x"ff",	--12738
		x"ff",	--12739
		x"ff",	--12740
		x"ff",	--12741
		x"ff",	--12742
		x"ff",	--12743
		x"ff",	--12744
		x"ff",	--12745
		x"ff",	--12746
		x"ff",	--12747
		x"ff",	--12748
		x"ff",	--12749
		x"ff",	--12750
		x"ff",	--12751
		x"ff",	--12752
		x"ff",	--12753
		x"ff",	--12754
		x"ff",	--12755
		x"ff",	--12756
		x"ff",	--12757
		x"ff",	--12758
		x"ff",	--12759
		x"ff",	--12760
		x"ff",	--12761
		x"ff",	--12762
		x"ff",	--12763
		x"ff",	--12764
		x"ff",	--12765
		x"ff",	--12766
		x"ff",	--12767
		x"ff",	--12768
		x"ff",	--12769
		x"ff",	--12770
		x"ff",	--12771
		x"ff",	--12772
		x"ff",	--12773
		x"ff",	--12774
		x"ff",	--12775
		x"ff",	--12776
		x"ff",	--12777
		x"ff",	--12778
		x"ff",	--12779
		x"ff",	--12780
		x"ff",	--12781
		x"ff",	--12782
		x"ff",	--12783
		x"ff",	--12784
		x"ff",	--12785
		x"ff",	--12786
		x"ff",	--12787
		x"ff",	--12788
		x"ff",	--12789
		x"ff",	--12790
		x"ff",	--12791
		x"ff",	--12792
		x"ff",	--12793
		x"ff",	--12794
		x"ff",	--12795
		x"ff",	--12796
		x"ff",	--12797
		x"ff",	--12798
		x"ff",	--12799
		x"ff",	--12800
		x"ff",	--12801
		x"ff",	--12802
		x"ff",	--12803
		x"ff",	--12804
		x"ff",	--12805
		x"ff",	--12806
		x"ff",	--12807
		x"ff",	--12808
		x"ff",	--12809
		x"ff",	--12810
		x"ff",	--12811
		x"ff",	--12812
		x"ff",	--12813
		x"ff",	--12814
		x"ff",	--12815
		x"ff",	--12816
		x"ff",	--12817
		x"ff",	--12818
		x"ff",	--12819
		x"ff",	--12820
		x"ff",	--12821
		x"ff",	--12822
		x"ff",	--12823
		x"ff",	--12824
		x"ff",	--12825
		x"ff",	--12826
		x"ff",	--12827
		x"ff",	--12828
		x"ff",	--12829
		x"ff",	--12830
		x"ff",	--12831
		x"ff",	--12832
		x"ff",	--12833
		x"ff",	--12834
		x"ff",	--12835
		x"ff",	--12836
		x"ff",	--12837
		x"ff",	--12838
		x"ff",	--12839
		x"ff",	--12840
		x"ff",	--12841
		x"ff",	--12842
		x"ff",	--12843
		x"ff",	--12844
		x"ff",	--12845
		x"ff",	--12846
		x"ff",	--12847
		x"ff",	--12848
		x"ff",	--12849
		x"ff",	--12850
		x"ff",	--12851
		x"ff",	--12852
		x"ff",	--12853
		x"ff",	--12854
		x"ff",	--12855
		x"ff",	--12856
		x"ff",	--12857
		x"ff",	--12858
		x"ff",	--12859
		x"ff",	--12860
		x"ff",	--12861
		x"ff",	--12862
		x"ff",	--12863
		x"ff",	--12864
		x"ff",	--12865
		x"ff",	--12866
		x"ff",	--12867
		x"ff",	--12868
		x"ff",	--12869
		x"ff",	--12870
		x"ff",	--12871
		x"ff",	--12872
		x"ff",	--12873
		x"ff",	--12874
		x"ff",	--12875
		x"ff",	--12876
		x"ff",	--12877
		x"ff",	--12878
		x"ff",	--12879
		x"ff",	--12880
		x"ff",	--12881
		x"ff",	--12882
		x"ff",	--12883
		x"ff",	--12884
		x"ff",	--12885
		x"ff",	--12886
		x"ff",	--12887
		x"ff",	--12888
		x"ff",	--12889
		x"ff",	--12890
		x"ff",	--12891
		x"ff",	--12892
		x"ff",	--12893
		x"ff",	--12894
		x"ff",	--12895
		x"ff",	--12896
		x"ff",	--12897
		x"ff",	--12898
		x"ff",	--12899
		x"ff",	--12900
		x"ff",	--12901
		x"ff",	--12902
		x"ff",	--12903
		x"ff",	--12904
		x"ff",	--12905
		x"ff",	--12906
		x"ff",	--12907
		x"ff",	--12908
		x"ff",	--12909
		x"ff",	--12910
		x"ff",	--12911
		x"ff",	--12912
		x"ff",	--12913
		x"ff",	--12914
		x"ff",	--12915
		x"ff",	--12916
		x"ff",	--12917
		x"ff",	--12918
		x"ff",	--12919
		x"ff",	--12920
		x"ff",	--12921
		x"ff",	--12922
		x"ff",	--12923
		x"ff",	--12924
		x"ff",	--12925
		x"ff",	--12926
		x"ff",	--12927
		x"ff",	--12928
		x"ff",	--12929
		x"ff",	--12930
		x"ff",	--12931
		x"ff",	--12932
		x"ff",	--12933
		x"ff",	--12934
		x"ff",	--12935
		x"ff",	--12936
		x"ff",	--12937
		x"ff",	--12938
		x"ff",	--12939
		x"ff",	--12940
		x"ff",	--12941
		x"ff",	--12942
		x"ff",	--12943
		x"ff",	--12944
		x"ff",	--12945
		x"ff",	--12946
		x"ff",	--12947
		x"ff",	--12948
		x"ff",	--12949
		x"ff",	--12950
		x"ff",	--12951
		x"ff",	--12952
		x"ff",	--12953
		x"ff",	--12954
		x"ff",	--12955
		x"ff",	--12956
		x"ff",	--12957
		x"ff",	--12958
		x"ff",	--12959
		x"ff",	--12960
		x"ff",	--12961
		x"ff",	--12962
		x"ff",	--12963
		x"ff",	--12964
		x"ff",	--12965
		x"ff",	--12966
		x"ff",	--12967
		x"ff",	--12968
		x"ff",	--12969
		x"ff",	--12970
		x"ff",	--12971
		x"ff",	--12972
		x"ff",	--12973
		x"ff",	--12974
		x"ff",	--12975
		x"ff",	--12976
		x"ff",	--12977
		x"ff",	--12978
		x"ff",	--12979
		x"ff",	--12980
		x"ff",	--12981
		x"ff",	--12982
		x"ff",	--12983
		x"ff",	--12984
		x"ff",	--12985
		x"ff",	--12986
		x"ff",	--12987
		x"ff",	--12988
		x"ff",	--12989
		x"ff",	--12990
		x"ff",	--12991
		x"ff",	--12992
		x"ff",	--12993
		x"ff",	--12994
		x"ff",	--12995
		x"ff",	--12996
		x"ff",	--12997
		x"ff",	--12998
		x"ff",	--12999
		x"ff",	--13000
		x"ff",	--13001
		x"ff",	--13002
		x"ff",	--13003
		x"ff",	--13004
		x"ff",	--13005
		x"ff",	--13006
		x"ff",	--13007
		x"ff",	--13008
		x"ff",	--13009
		x"ff",	--13010
		x"ff",	--13011
		x"ff",	--13012
		x"ff",	--13013
		x"ff",	--13014
		x"ff",	--13015
		x"ff",	--13016
		x"ff",	--13017
		x"ff",	--13018
		x"ff",	--13019
		x"ff",	--13020
		x"ff",	--13021
		x"ff",	--13022
		x"ff",	--13023
		x"ff",	--13024
		x"ff",	--13025
		x"ff",	--13026
		x"ff",	--13027
		x"ff",	--13028
		x"ff",	--13029
		x"ff",	--13030
		x"ff",	--13031
		x"ff",	--13032
		x"ff",	--13033
		x"ff",	--13034
		x"ff",	--13035
		x"ff",	--13036
		x"ff",	--13037
		x"ff",	--13038
		x"ff",	--13039
		x"ff",	--13040
		x"ff",	--13041
		x"ff",	--13042
		x"ff",	--13043
		x"ff",	--13044
		x"ff",	--13045
		x"ff",	--13046
		x"ff",	--13047
		x"ff",	--13048
		x"ff",	--13049
		x"ff",	--13050
		x"ff",	--13051
		x"ff",	--13052
		x"ff",	--13053
		x"ff",	--13054
		x"ff",	--13055
		x"ff",	--13056
		x"ff",	--13057
		x"ff",	--13058
		x"ff",	--13059
		x"ff",	--13060
		x"ff",	--13061
		x"ff",	--13062
		x"ff",	--13063
		x"ff",	--13064
		x"ff",	--13065
		x"ff",	--13066
		x"ff",	--13067
		x"ff",	--13068
		x"ff",	--13069
		x"ff",	--13070
		x"ff",	--13071
		x"ff",	--13072
		x"ff",	--13073
		x"ff",	--13074
		x"ff",	--13075
		x"ff",	--13076
		x"ff",	--13077
		x"ff",	--13078
		x"ff",	--13079
		x"ff",	--13080
		x"ff",	--13081
		x"ff",	--13082
		x"ff",	--13083
		x"ff",	--13084
		x"ff",	--13085
		x"ff",	--13086
		x"ff",	--13087
		x"ff",	--13088
		x"ff",	--13089
		x"ff",	--13090
		x"ff",	--13091
		x"ff",	--13092
		x"ff",	--13093
		x"ff",	--13094
		x"ff",	--13095
		x"ff",	--13096
		x"ff",	--13097
		x"ff",	--13098
		x"ff",	--13099
		x"ff",	--13100
		x"ff",	--13101
		x"ff",	--13102
		x"ff",	--13103
		x"ff",	--13104
		x"ff",	--13105
		x"ff",	--13106
		x"ff",	--13107
		x"ff",	--13108
		x"ff",	--13109
		x"ff",	--13110
		x"ff",	--13111
		x"ff",	--13112
		x"ff",	--13113
		x"ff",	--13114
		x"ff",	--13115
		x"ff",	--13116
		x"ff",	--13117
		x"ff",	--13118
		x"ff",	--13119
		x"ff",	--13120
		x"ff",	--13121
		x"ff",	--13122
		x"ff",	--13123
		x"ff",	--13124
		x"ff",	--13125
		x"ff",	--13126
		x"ff",	--13127
		x"ff",	--13128
		x"ff",	--13129
		x"ff",	--13130
		x"ff",	--13131
		x"ff",	--13132
		x"ff",	--13133
		x"ff",	--13134
		x"ff",	--13135
		x"ff",	--13136
		x"ff",	--13137
		x"ff",	--13138
		x"ff",	--13139
		x"ff",	--13140
		x"ff",	--13141
		x"ff",	--13142
		x"ff",	--13143
		x"ff",	--13144
		x"ff",	--13145
		x"ff",	--13146
		x"ff",	--13147
		x"ff",	--13148
		x"ff",	--13149
		x"ff",	--13150
		x"ff",	--13151
		x"ff",	--13152
		x"ff",	--13153
		x"ff",	--13154
		x"ff",	--13155
		x"ff",	--13156
		x"ff",	--13157
		x"ff",	--13158
		x"ff",	--13159
		x"ff",	--13160
		x"ff",	--13161
		x"ff",	--13162
		x"ff",	--13163
		x"ff",	--13164
		x"ff",	--13165
		x"ff",	--13166
		x"ff",	--13167
		x"ff",	--13168
		x"ff",	--13169
		x"ff",	--13170
		x"ff",	--13171
		x"ff",	--13172
		x"ff",	--13173
		x"ff",	--13174
		x"ff",	--13175
		x"ff",	--13176
		x"ff",	--13177
		x"ff",	--13178
		x"ff",	--13179
		x"ff",	--13180
		x"ff",	--13181
		x"ff",	--13182
		x"ff",	--13183
		x"ff",	--13184
		x"ff",	--13185
		x"ff",	--13186
		x"ff",	--13187
		x"ff",	--13188
		x"ff",	--13189
		x"ff",	--13190
		x"ff",	--13191
		x"ff",	--13192
		x"ff",	--13193
		x"ff",	--13194
		x"ff",	--13195
		x"ff",	--13196
		x"ff",	--13197
		x"ff",	--13198
		x"ff",	--13199
		x"ff",	--13200
		x"ff",	--13201
		x"ff",	--13202
		x"ff",	--13203
		x"ff",	--13204
		x"ff",	--13205
		x"ff",	--13206
		x"ff",	--13207
		x"ff",	--13208
		x"ff",	--13209
		x"ff",	--13210
		x"ff",	--13211
		x"ff",	--13212
		x"ff",	--13213
		x"ff",	--13214
		x"ff",	--13215
		x"ff",	--13216
		x"ff",	--13217
		x"ff",	--13218
		x"ff",	--13219
		x"ff",	--13220
		x"ff",	--13221
		x"ff",	--13222
		x"ff",	--13223
		x"ff",	--13224
		x"ff",	--13225
		x"ff",	--13226
		x"ff",	--13227
		x"ff",	--13228
		x"ff",	--13229
		x"ff",	--13230
		x"ff",	--13231
		x"ff",	--13232
		x"ff",	--13233
		x"ff",	--13234
		x"ff",	--13235
		x"ff",	--13236
		x"ff",	--13237
		x"ff",	--13238
		x"ff",	--13239
		x"ff",	--13240
		x"ff",	--13241
		x"ff",	--13242
		x"ff",	--13243
		x"ff",	--13244
		x"ff",	--13245
		x"ff",	--13246
		x"ff",	--13247
		x"ff",	--13248
		x"ff",	--13249
		x"ff",	--13250
		x"ff",	--13251
		x"ff",	--13252
		x"ff",	--13253
		x"ff",	--13254
		x"ff",	--13255
		x"ff",	--13256
		x"ff",	--13257
		x"ff",	--13258
		x"ff",	--13259
		x"ff",	--13260
		x"ff",	--13261
		x"ff",	--13262
		x"ff",	--13263
		x"ff",	--13264
		x"ff",	--13265
		x"ff",	--13266
		x"ff",	--13267
		x"ff",	--13268
		x"ff",	--13269
		x"ff",	--13270
		x"ff",	--13271
		x"ff",	--13272
		x"ff",	--13273
		x"ff",	--13274
		x"ff",	--13275
		x"ff",	--13276
		x"ff",	--13277
		x"ff",	--13278
		x"ff",	--13279
		x"ff",	--13280
		x"ff",	--13281
		x"ff",	--13282
		x"ff",	--13283
		x"ff",	--13284
		x"ff",	--13285
		x"ff",	--13286
		x"ff",	--13287
		x"ff",	--13288
		x"ff",	--13289
		x"ff",	--13290
		x"ff",	--13291
		x"ff",	--13292
		x"ff",	--13293
		x"ff",	--13294
		x"ff",	--13295
		x"ff",	--13296
		x"ff",	--13297
		x"ff",	--13298
		x"ff",	--13299
		x"ff",	--13300
		x"ff",	--13301
		x"ff",	--13302
		x"ff",	--13303
		x"ff",	--13304
		x"ff",	--13305
		x"ff",	--13306
		x"ff",	--13307
		x"ff",	--13308
		x"ff",	--13309
		x"ff",	--13310
		x"ff",	--13311
		x"ff",	--13312
		x"ff",	--13313
		x"ff",	--13314
		x"ff",	--13315
		x"ff",	--13316
		x"ff",	--13317
		x"ff",	--13318
		x"ff",	--13319
		x"ff",	--13320
		x"ff",	--13321
		x"ff",	--13322
		x"ff",	--13323
		x"ff",	--13324
		x"ff",	--13325
		x"ff",	--13326
		x"ff",	--13327
		x"ff",	--13328
		x"ff",	--13329
		x"ff",	--13330
		x"ff",	--13331
		x"ff",	--13332
		x"ff",	--13333
		x"ff",	--13334
		x"ff",	--13335
		x"ff",	--13336
		x"ff",	--13337
		x"ff",	--13338
		x"ff",	--13339
		x"ff",	--13340
		x"ff",	--13341
		x"ff",	--13342
		x"ff",	--13343
		x"ff",	--13344
		x"ff",	--13345
		x"ff",	--13346
		x"ff",	--13347
		x"ff",	--13348
		x"ff",	--13349
		x"ff",	--13350
		x"ff",	--13351
		x"ff",	--13352
		x"ff",	--13353
		x"ff",	--13354
		x"ff",	--13355
		x"ff",	--13356
		x"ff",	--13357
		x"ff",	--13358
		x"ff",	--13359
		x"ff",	--13360
		x"ff",	--13361
		x"ff",	--13362
		x"ff",	--13363
		x"ff",	--13364
		x"ff",	--13365
		x"ff",	--13366
		x"ff",	--13367
		x"ff",	--13368
		x"ff",	--13369
		x"ff",	--13370
		x"ff",	--13371
		x"ff",	--13372
		x"ff",	--13373
		x"ff",	--13374
		x"ff",	--13375
		x"ff",	--13376
		x"ff",	--13377
		x"ff",	--13378
		x"ff",	--13379
		x"ff",	--13380
		x"ff",	--13381
		x"ff",	--13382
		x"ff",	--13383
		x"ff",	--13384
		x"ff",	--13385
		x"ff",	--13386
		x"ff",	--13387
		x"ff",	--13388
		x"ff",	--13389
		x"ff",	--13390
		x"ff",	--13391
		x"ff",	--13392
		x"ff",	--13393
		x"ff",	--13394
		x"ff",	--13395
		x"ff",	--13396
		x"ff",	--13397
		x"ff",	--13398
		x"ff",	--13399
		x"ff",	--13400
		x"ff",	--13401
		x"ff",	--13402
		x"ff",	--13403
		x"ff",	--13404
		x"ff",	--13405
		x"ff",	--13406
		x"ff",	--13407
		x"ff",	--13408
		x"ff",	--13409
		x"ff",	--13410
		x"ff",	--13411
		x"ff",	--13412
		x"ff",	--13413
		x"ff",	--13414
		x"ff",	--13415
		x"ff",	--13416
		x"ff",	--13417
		x"ff",	--13418
		x"ff",	--13419
		x"ff",	--13420
		x"ff",	--13421
		x"ff",	--13422
		x"ff",	--13423
		x"ff",	--13424
		x"ff",	--13425
		x"ff",	--13426
		x"ff",	--13427
		x"ff",	--13428
		x"ff",	--13429
		x"ff",	--13430
		x"ff",	--13431
		x"ff",	--13432
		x"ff",	--13433
		x"ff",	--13434
		x"ff",	--13435
		x"ff",	--13436
		x"ff",	--13437
		x"ff",	--13438
		x"ff",	--13439
		x"ff",	--13440
		x"ff",	--13441
		x"ff",	--13442
		x"ff",	--13443
		x"ff",	--13444
		x"ff",	--13445
		x"ff",	--13446
		x"ff",	--13447
		x"ff",	--13448
		x"ff",	--13449
		x"ff",	--13450
		x"ff",	--13451
		x"ff",	--13452
		x"ff",	--13453
		x"ff",	--13454
		x"ff",	--13455
		x"ff",	--13456
		x"ff",	--13457
		x"ff",	--13458
		x"ff",	--13459
		x"ff",	--13460
		x"ff",	--13461
		x"ff",	--13462
		x"ff",	--13463
		x"ff",	--13464
		x"ff",	--13465
		x"ff",	--13466
		x"ff",	--13467
		x"ff",	--13468
		x"ff",	--13469
		x"ff",	--13470
		x"ff",	--13471
		x"ff",	--13472
		x"ff",	--13473
		x"ff",	--13474
		x"ff",	--13475
		x"ff",	--13476
		x"ff",	--13477
		x"ff",	--13478
		x"ff",	--13479
		x"ff",	--13480
		x"ff",	--13481
		x"ff",	--13482
		x"ff",	--13483
		x"ff",	--13484
		x"ff",	--13485
		x"ff",	--13486
		x"ff",	--13487
		x"ff",	--13488
		x"ff",	--13489
		x"ff",	--13490
		x"ff",	--13491
		x"ff",	--13492
		x"ff",	--13493
		x"ff",	--13494
		x"ff",	--13495
		x"ff",	--13496
		x"ff",	--13497
		x"ff",	--13498
		x"ff",	--13499
		x"ff",	--13500
		x"ff",	--13501
		x"ff",	--13502
		x"ff",	--13503
		x"ff",	--13504
		x"ff",	--13505
		x"ff",	--13506
		x"ff",	--13507
		x"ff",	--13508
		x"ff",	--13509
		x"ff",	--13510
		x"ff",	--13511
		x"ff",	--13512
		x"ff",	--13513
		x"ff",	--13514
		x"ff",	--13515
		x"ff",	--13516
		x"ff",	--13517
		x"ff",	--13518
		x"ff",	--13519
		x"ff",	--13520
		x"ff",	--13521
		x"ff",	--13522
		x"ff",	--13523
		x"ff",	--13524
		x"ff",	--13525
		x"ff",	--13526
		x"ff",	--13527
		x"ff",	--13528
		x"ff",	--13529
		x"ff",	--13530
		x"ff",	--13531
		x"ff",	--13532
		x"ff",	--13533
		x"ff",	--13534
		x"ff",	--13535
		x"ff",	--13536
		x"ff",	--13537
		x"ff",	--13538
		x"ff",	--13539
		x"ff",	--13540
		x"ff",	--13541
		x"ff",	--13542
		x"ff",	--13543
		x"ff",	--13544
		x"ff",	--13545
		x"ff",	--13546
		x"ff",	--13547
		x"ff",	--13548
		x"ff",	--13549
		x"ff",	--13550
		x"ff",	--13551
		x"ff",	--13552
		x"ff",	--13553
		x"ff",	--13554
		x"ff",	--13555
		x"ff",	--13556
		x"ff",	--13557
		x"ff",	--13558
		x"ff",	--13559
		x"ff",	--13560
		x"ff",	--13561
		x"ff",	--13562
		x"ff",	--13563
		x"ff",	--13564
		x"ff",	--13565
		x"ff",	--13566
		x"ff",	--13567
		x"ff",	--13568
		x"ff",	--13569
		x"ff",	--13570
		x"ff",	--13571
		x"ff",	--13572
		x"ff",	--13573
		x"ff",	--13574
		x"ff",	--13575
		x"ff",	--13576
		x"ff",	--13577
		x"ff",	--13578
		x"ff",	--13579
		x"ff",	--13580
		x"ff",	--13581
		x"ff",	--13582
		x"ff",	--13583
		x"ff",	--13584
		x"ff",	--13585
		x"ff",	--13586
		x"ff",	--13587
		x"ff",	--13588
		x"ff",	--13589
		x"ff",	--13590
		x"ff",	--13591
		x"ff",	--13592
		x"ff",	--13593
		x"ff",	--13594
		x"ff",	--13595
		x"ff",	--13596
		x"ff",	--13597
		x"ff",	--13598
		x"ff",	--13599
		x"ff",	--13600
		x"ff",	--13601
		x"ff",	--13602
		x"ff",	--13603
		x"ff",	--13604
		x"ff",	--13605
		x"ff",	--13606
		x"ff",	--13607
		x"ff",	--13608
		x"ff",	--13609
		x"ff",	--13610
		x"ff",	--13611
		x"ff",	--13612
		x"ff",	--13613
		x"ff",	--13614
		x"ff",	--13615
		x"ff",	--13616
		x"ff",	--13617
		x"ff",	--13618
		x"ff",	--13619
		x"ff",	--13620
		x"ff",	--13621
		x"ff",	--13622
		x"ff",	--13623
		x"ff",	--13624
		x"ff",	--13625
		x"ff",	--13626
		x"ff",	--13627
		x"ff",	--13628
		x"ff",	--13629
		x"ff",	--13630
		x"ff",	--13631
		x"ff",	--13632
		x"ff",	--13633
		x"ff",	--13634
		x"ff",	--13635
		x"ff",	--13636
		x"ff",	--13637
		x"ff",	--13638
		x"ff",	--13639
		x"ff",	--13640
		x"ff",	--13641
		x"ff",	--13642
		x"ff",	--13643
		x"ff",	--13644
		x"ff",	--13645
		x"ff",	--13646
		x"ff",	--13647
		x"ff",	--13648
		x"ff",	--13649
		x"ff",	--13650
		x"ff",	--13651
		x"ff",	--13652
		x"ff",	--13653
		x"ff",	--13654
		x"ff",	--13655
		x"ff",	--13656
		x"ff",	--13657
		x"ff",	--13658
		x"ff",	--13659
		x"ff",	--13660
		x"ff",	--13661
		x"ff",	--13662
		x"ff",	--13663
		x"ff",	--13664
		x"ff",	--13665
		x"ff",	--13666
		x"ff",	--13667
		x"ff",	--13668
		x"ff",	--13669
		x"ff",	--13670
		x"ff",	--13671
		x"ff",	--13672
		x"ff",	--13673
		x"ff",	--13674
		x"ff",	--13675
		x"ff",	--13676
		x"ff",	--13677
		x"ff",	--13678
		x"ff",	--13679
		x"ff",	--13680
		x"ff",	--13681
		x"ff",	--13682
		x"ff",	--13683
		x"ff",	--13684
		x"ff",	--13685
		x"ff",	--13686
		x"ff",	--13687
		x"ff",	--13688
		x"ff",	--13689
		x"ff",	--13690
		x"ff",	--13691
		x"ff",	--13692
		x"ff",	--13693
		x"ff",	--13694
		x"ff",	--13695
		x"ff",	--13696
		x"ff",	--13697
		x"ff",	--13698
		x"ff",	--13699
		x"ff",	--13700
		x"ff",	--13701
		x"ff",	--13702
		x"ff",	--13703
		x"ff",	--13704
		x"ff",	--13705
		x"ff",	--13706
		x"ff",	--13707
		x"ff",	--13708
		x"ff",	--13709
		x"ff",	--13710
		x"ff",	--13711
		x"ff",	--13712
		x"ff",	--13713
		x"ff",	--13714
		x"ff",	--13715
		x"ff",	--13716
		x"ff",	--13717
		x"ff",	--13718
		x"ff",	--13719
		x"ff",	--13720
		x"ff",	--13721
		x"ff",	--13722
		x"ff",	--13723
		x"ff",	--13724
		x"ff",	--13725
		x"ff",	--13726
		x"ff",	--13727
		x"ff",	--13728
		x"ff",	--13729
		x"ff",	--13730
		x"ff",	--13731
		x"ff",	--13732
		x"ff",	--13733
		x"ff",	--13734
		x"ff",	--13735
		x"ff",	--13736
		x"ff",	--13737
		x"ff",	--13738
		x"ff",	--13739
		x"ff",	--13740
		x"ff",	--13741
		x"ff",	--13742
		x"ff",	--13743
		x"ff",	--13744
		x"ff",	--13745
		x"ff",	--13746
		x"ff",	--13747
		x"ff",	--13748
		x"ff",	--13749
		x"ff",	--13750
		x"ff",	--13751
		x"ff",	--13752
		x"ff",	--13753
		x"ff",	--13754
		x"ff",	--13755
		x"ff",	--13756
		x"ff",	--13757
		x"ff",	--13758
		x"ff",	--13759
		x"ff",	--13760
		x"ff",	--13761
		x"ff",	--13762
		x"ff",	--13763
		x"ff",	--13764
		x"ff",	--13765
		x"ff",	--13766
		x"ff",	--13767
		x"ff",	--13768
		x"ff",	--13769
		x"ff",	--13770
		x"ff",	--13771
		x"ff",	--13772
		x"ff",	--13773
		x"ff",	--13774
		x"ff",	--13775
		x"ff",	--13776
		x"ff",	--13777
		x"ff",	--13778
		x"ff",	--13779
		x"ff",	--13780
		x"ff",	--13781
		x"ff",	--13782
		x"ff",	--13783
		x"ff",	--13784
		x"ff",	--13785
		x"ff",	--13786
		x"ff",	--13787
		x"ff",	--13788
		x"ff",	--13789
		x"ff",	--13790
		x"ff",	--13791
		x"ff",	--13792
		x"ff",	--13793
		x"ff",	--13794
		x"ff",	--13795
		x"ff",	--13796
		x"ff",	--13797
		x"ff",	--13798
		x"ff",	--13799
		x"ff",	--13800
		x"ff",	--13801
		x"ff",	--13802
		x"ff",	--13803
		x"ff",	--13804
		x"ff",	--13805
		x"ff",	--13806
		x"ff",	--13807
		x"ff",	--13808
		x"ff",	--13809
		x"ff",	--13810
		x"ff",	--13811
		x"ff",	--13812
		x"ff",	--13813
		x"ff",	--13814
		x"ff",	--13815
		x"ff",	--13816
		x"ff",	--13817
		x"ff",	--13818
		x"ff",	--13819
		x"ff",	--13820
		x"ff",	--13821
		x"ff",	--13822
		x"ff",	--13823
		x"ff",	--13824
		x"ff",	--13825
		x"ff",	--13826
		x"ff",	--13827
		x"ff",	--13828
		x"ff",	--13829
		x"ff",	--13830
		x"ff",	--13831
		x"ff",	--13832
		x"ff",	--13833
		x"ff",	--13834
		x"ff",	--13835
		x"ff",	--13836
		x"ff",	--13837
		x"ff",	--13838
		x"ff",	--13839
		x"ff",	--13840
		x"ff",	--13841
		x"ff",	--13842
		x"ff",	--13843
		x"ff",	--13844
		x"ff",	--13845
		x"ff",	--13846
		x"ff",	--13847
		x"ff",	--13848
		x"ff",	--13849
		x"ff",	--13850
		x"ff",	--13851
		x"ff",	--13852
		x"ff",	--13853
		x"ff",	--13854
		x"ff",	--13855
		x"ff",	--13856
		x"ff",	--13857
		x"ff",	--13858
		x"ff",	--13859
		x"ff",	--13860
		x"ff",	--13861
		x"ff",	--13862
		x"ff",	--13863
		x"ff",	--13864
		x"ff",	--13865
		x"ff",	--13866
		x"ff",	--13867
		x"ff",	--13868
		x"ff",	--13869
		x"ff",	--13870
		x"ff",	--13871
		x"ff",	--13872
		x"ff",	--13873
		x"ff",	--13874
		x"ff",	--13875
		x"ff",	--13876
		x"ff",	--13877
		x"ff",	--13878
		x"ff",	--13879
		x"ff",	--13880
		x"ff",	--13881
		x"ff",	--13882
		x"ff",	--13883
		x"ff",	--13884
		x"ff",	--13885
		x"ff",	--13886
		x"ff",	--13887
		x"ff",	--13888
		x"ff",	--13889
		x"ff",	--13890
		x"ff",	--13891
		x"ff",	--13892
		x"ff",	--13893
		x"ff",	--13894
		x"ff",	--13895
		x"ff",	--13896
		x"ff",	--13897
		x"ff",	--13898
		x"ff",	--13899
		x"ff",	--13900
		x"ff",	--13901
		x"ff",	--13902
		x"ff",	--13903
		x"ff",	--13904
		x"ff",	--13905
		x"ff",	--13906
		x"ff",	--13907
		x"ff",	--13908
		x"ff",	--13909
		x"ff",	--13910
		x"ff",	--13911
		x"ff",	--13912
		x"ff",	--13913
		x"ff",	--13914
		x"ff",	--13915
		x"ff",	--13916
		x"ff",	--13917
		x"ff",	--13918
		x"ff",	--13919
		x"ff",	--13920
		x"ff",	--13921
		x"ff",	--13922
		x"ff",	--13923
		x"ff",	--13924
		x"ff",	--13925
		x"ff",	--13926
		x"ff",	--13927
		x"ff",	--13928
		x"ff",	--13929
		x"ff",	--13930
		x"ff",	--13931
		x"ff",	--13932
		x"ff",	--13933
		x"ff",	--13934
		x"ff",	--13935
		x"ff",	--13936
		x"ff",	--13937
		x"ff",	--13938
		x"ff",	--13939
		x"ff",	--13940
		x"ff",	--13941
		x"ff",	--13942
		x"ff",	--13943
		x"ff",	--13944
		x"ff",	--13945
		x"ff",	--13946
		x"ff",	--13947
		x"ff",	--13948
		x"ff",	--13949
		x"ff",	--13950
		x"ff",	--13951
		x"ff",	--13952
		x"ff",	--13953
		x"ff",	--13954
		x"ff",	--13955
		x"ff",	--13956
		x"ff",	--13957
		x"ff",	--13958
		x"ff",	--13959
		x"ff",	--13960
		x"ff",	--13961
		x"ff",	--13962
		x"ff",	--13963
		x"ff",	--13964
		x"ff",	--13965
		x"ff",	--13966
		x"ff",	--13967
		x"ff",	--13968
		x"ff",	--13969
		x"ff",	--13970
		x"ff",	--13971
		x"ff",	--13972
		x"ff",	--13973
		x"ff",	--13974
		x"ff",	--13975
		x"ff",	--13976
		x"ff",	--13977
		x"ff",	--13978
		x"ff",	--13979
		x"ff",	--13980
		x"ff",	--13981
		x"ff",	--13982
		x"ff",	--13983
		x"ff",	--13984
		x"ff",	--13985
		x"ff",	--13986
		x"ff",	--13987
		x"ff",	--13988
		x"ff",	--13989
		x"ff",	--13990
		x"ff",	--13991
		x"ff",	--13992
		x"ff",	--13993
		x"ff",	--13994
		x"ff",	--13995
		x"ff",	--13996
		x"ff",	--13997
		x"ff",	--13998
		x"ff",	--13999
		x"ff",	--14000
		x"ff",	--14001
		x"ff",	--14002
		x"ff",	--14003
		x"ff",	--14004
		x"ff",	--14005
		x"ff",	--14006
		x"ff",	--14007
		x"ff",	--14008
		x"ff",	--14009
		x"ff",	--14010
		x"ff",	--14011
		x"ff",	--14012
		x"ff",	--14013
		x"ff",	--14014
		x"ff",	--14015
		x"ff",	--14016
		x"ff",	--14017
		x"ff",	--14018
		x"ff",	--14019
		x"ff",	--14020
		x"ff",	--14021
		x"ff",	--14022
		x"ff",	--14023
		x"ff",	--14024
		x"ff",	--14025
		x"ff",	--14026
		x"ff",	--14027
		x"ff",	--14028
		x"ff",	--14029
		x"ff",	--14030
		x"ff",	--14031
		x"ff",	--14032
		x"ff",	--14033
		x"ff",	--14034
		x"ff",	--14035
		x"ff",	--14036
		x"ff",	--14037
		x"ff",	--14038
		x"ff",	--14039
		x"ff",	--14040
		x"ff",	--14041
		x"ff",	--14042
		x"ff",	--14043
		x"ff",	--14044
		x"ff",	--14045
		x"ff",	--14046
		x"ff",	--14047
		x"ff",	--14048
		x"ff",	--14049
		x"ff",	--14050
		x"ff",	--14051
		x"ff",	--14052
		x"ff",	--14053
		x"ff",	--14054
		x"ff",	--14055
		x"ff",	--14056
		x"ff",	--14057
		x"ff",	--14058
		x"ff",	--14059
		x"ff",	--14060
		x"ff",	--14061
		x"ff",	--14062
		x"ff",	--14063
		x"ff",	--14064
		x"ff",	--14065
		x"ff",	--14066
		x"ff",	--14067
		x"ff",	--14068
		x"ff",	--14069
		x"ff",	--14070
		x"ff",	--14071
		x"ff",	--14072
		x"ff",	--14073
		x"ff",	--14074
		x"ff",	--14075
		x"ff",	--14076
		x"ff",	--14077
		x"ff",	--14078
		x"ff",	--14079
		x"ff",	--14080
		x"ff",	--14081
		x"ff",	--14082
		x"ff",	--14083
		x"ff",	--14084
		x"ff",	--14085
		x"ff",	--14086
		x"ff",	--14087
		x"ff",	--14088
		x"ff",	--14089
		x"ff",	--14090
		x"ff",	--14091
		x"ff",	--14092
		x"ff",	--14093
		x"ff",	--14094
		x"ff",	--14095
		x"ff",	--14096
		x"ff",	--14097
		x"ff",	--14098
		x"ff",	--14099
		x"ff",	--14100
		x"ff",	--14101
		x"ff",	--14102
		x"ff",	--14103
		x"ff",	--14104
		x"ff",	--14105
		x"ff",	--14106
		x"ff",	--14107
		x"ff",	--14108
		x"ff",	--14109
		x"ff",	--14110
		x"ff",	--14111
		x"ff",	--14112
		x"ff",	--14113
		x"ff",	--14114
		x"ff",	--14115
		x"ff",	--14116
		x"ff",	--14117
		x"ff",	--14118
		x"ff",	--14119
		x"ff",	--14120
		x"ff",	--14121
		x"ff",	--14122
		x"ff",	--14123
		x"ff",	--14124
		x"ff",	--14125
		x"ff",	--14126
		x"ff",	--14127
		x"ff",	--14128
		x"ff",	--14129
		x"ff",	--14130
		x"ff",	--14131
		x"ff",	--14132
		x"ff",	--14133
		x"ff",	--14134
		x"ff",	--14135
		x"ff",	--14136
		x"ff",	--14137
		x"ff",	--14138
		x"ff",	--14139
		x"ff",	--14140
		x"ff",	--14141
		x"ff",	--14142
		x"ff",	--14143
		x"ff",	--14144
		x"ff",	--14145
		x"ff",	--14146
		x"ff",	--14147
		x"ff",	--14148
		x"ff",	--14149
		x"ff",	--14150
		x"ff",	--14151
		x"ff",	--14152
		x"ff",	--14153
		x"ff",	--14154
		x"ff",	--14155
		x"ff",	--14156
		x"ff",	--14157
		x"ff",	--14158
		x"ff",	--14159
		x"ff",	--14160
		x"ff",	--14161
		x"ff",	--14162
		x"ff",	--14163
		x"ff",	--14164
		x"ff",	--14165
		x"ff",	--14166
		x"ff",	--14167
		x"ff",	--14168
		x"ff",	--14169
		x"ff",	--14170
		x"ff",	--14171
		x"ff",	--14172
		x"ff",	--14173
		x"ff",	--14174
		x"ff",	--14175
		x"ff",	--14176
		x"ff",	--14177
		x"ff",	--14178
		x"ff",	--14179
		x"ff",	--14180
		x"ff",	--14181
		x"ff",	--14182
		x"ff",	--14183
		x"ff",	--14184
		x"ff",	--14185
		x"ff",	--14186
		x"ff",	--14187
		x"ff",	--14188
		x"ff",	--14189
		x"ff",	--14190
		x"ff",	--14191
		x"ff",	--14192
		x"ff",	--14193
		x"ff",	--14194
		x"ff",	--14195
		x"ff",	--14196
		x"ff",	--14197
		x"ff",	--14198
		x"ff",	--14199
		x"ff",	--14200
		x"ff",	--14201
		x"ff",	--14202
		x"ff",	--14203
		x"ff",	--14204
		x"ff",	--14205
		x"ff",	--14206
		x"ff",	--14207
		x"ff",	--14208
		x"ff",	--14209
		x"ff",	--14210
		x"ff",	--14211
		x"ff",	--14212
		x"ff",	--14213
		x"ff",	--14214
		x"ff",	--14215
		x"ff",	--14216
		x"ff",	--14217
		x"ff",	--14218
		x"ff",	--14219
		x"ff",	--14220
		x"ff",	--14221
		x"ff",	--14222
		x"ff",	--14223
		x"ff",	--14224
		x"ff",	--14225
		x"ff",	--14226
		x"ff",	--14227
		x"ff",	--14228
		x"ff",	--14229
		x"ff",	--14230
		x"ff",	--14231
		x"ff",	--14232
		x"ff",	--14233
		x"ff",	--14234
		x"ff",	--14235
		x"ff",	--14236
		x"ff",	--14237
		x"ff",	--14238
		x"ff",	--14239
		x"ff",	--14240
		x"ff",	--14241
		x"ff",	--14242
		x"ff",	--14243
		x"ff",	--14244
		x"ff",	--14245
		x"ff",	--14246
		x"ff",	--14247
		x"ff",	--14248
		x"ff",	--14249
		x"ff",	--14250
		x"ff",	--14251
		x"ff",	--14252
		x"ff",	--14253
		x"ff",	--14254
		x"ff",	--14255
		x"ff",	--14256
		x"ff",	--14257
		x"ff",	--14258
		x"ff",	--14259
		x"ff",	--14260
		x"ff",	--14261
		x"ff",	--14262
		x"ff",	--14263
		x"ff",	--14264
		x"ff",	--14265
		x"ff",	--14266
		x"ff",	--14267
		x"ff",	--14268
		x"ff",	--14269
		x"ff",	--14270
		x"ff",	--14271
		x"ff",	--14272
		x"ff",	--14273
		x"ff",	--14274
		x"ff",	--14275
		x"ff",	--14276
		x"ff",	--14277
		x"ff",	--14278
		x"ff",	--14279
		x"ff",	--14280
		x"ff",	--14281
		x"ff",	--14282
		x"ff",	--14283
		x"ff",	--14284
		x"ff",	--14285
		x"ff",	--14286
		x"ff",	--14287
		x"ff",	--14288
		x"ff",	--14289
		x"ff",	--14290
		x"ff",	--14291
		x"ff",	--14292
		x"ff",	--14293
		x"ff",	--14294
		x"ff",	--14295
		x"ff",	--14296
		x"ff",	--14297
		x"ff",	--14298
		x"ff",	--14299
		x"ff",	--14300
		x"ff",	--14301
		x"ff",	--14302
		x"ff",	--14303
		x"ff",	--14304
		x"ff",	--14305
		x"ff",	--14306
		x"ff",	--14307
		x"ff",	--14308
		x"ff",	--14309
		x"ff",	--14310
		x"ff",	--14311
		x"ff",	--14312
		x"ff",	--14313
		x"ff",	--14314
		x"ff",	--14315
		x"ff",	--14316
		x"ff",	--14317
		x"ff",	--14318
		x"ff",	--14319
		x"ff",	--14320
		x"ff",	--14321
		x"ff",	--14322
		x"ff",	--14323
		x"ff",	--14324
		x"ff",	--14325
		x"ff",	--14326
		x"ff",	--14327
		x"ff",	--14328
		x"ff",	--14329
		x"ff",	--14330
		x"ff",	--14331
		x"ff",	--14332
		x"ff",	--14333
		x"ff",	--14334
		x"ff",	--14335
		x"ff",	--14336
		x"ff",	--14337
		x"ff",	--14338
		x"ff",	--14339
		x"ff",	--14340
		x"ff",	--14341
		x"ff",	--14342
		x"ff",	--14343
		x"ff",	--14344
		x"ff",	--14345
		x"ff",	--14346
		x"ff",	--14347
		x"ff",	--14348
		x"ff",	--14349
		x"ff",	--14350
		x"ff",	--14351
		x"ff",	--14352
		x"ff",	--14353
		x"ff",	--14354
		x"ff",	--14355
		x"ff",	--14356
		x"ff",	--14357
		x"ff",	--14358
		x"ff",	--14359
		x"ff",	--14360
		x"ff",	--14361
		x"ff",	--14362
		x"ff",	--14363
		x"ff",	--14364
		x"ff",	--14365
		x"ff",	--14366
		x"ff",	--14367
		x"ff",	--14368
		x"ff",	--14369
		x"ff",	--14370
		x"ff",	--14371
		x"ff",	--14372
		x"ff",	--14373
		x"ff",	--14374
		x"ff",	--14375
		x"ff",	--14376
		x"ff",	--14377
		x"ff",	--14378
		x"ff",	--14379
		x"ff",	--14380
		x"ff",	--14381
		x"ff",	--14382
		x"ff",	--14383
		x"ff",	--14384
		x"ff",	--14385
		x"ff",	--14386
		x"ff",	--14387
		x"ff",	--14388
		x"ff",	--14389
		x"ff",	--14390
		x"ff",	--14391
		x"ff",	--14392
		x"ff",	--14393
		x"ff",	--14394
		x"ff",	--14395
		x"ff",	--14396
		x"ff",	--14397
		x"ff",	--14398
		x"ff",	--14399
		x"ff",	--14400
		x"ff",	--14401
		x"ff",	--14402
		x"ff",	--14403
		x"ff",	--14404
		x"ff",	--14405
		x"ff",	--14406
		x"ff",	--14407
		x"ff",	--14408
		x"ff",	--14409
		x"ff",	--14410
		x"ff",	--14411
		x"ff",	--14412
		x"ff",	--14413
		x"ff",	--14414
		x"ff",	--14415
		x"ff",	--14416
		x"ff",	--14417
		x"ff",	--14418
		x"ff",	--14419
		x"ff",	--14420
		x"ff",	--14421
		x"ff",	--14422
		x"ff",	--14423
		x"ff",	--14424
		x"ff",	--14425
		x"ff",	--14426
		x"ff",	--14427
		x"ff",	--14428
		x"ff",	--14429
		x"ff",	--14430
		x"ff",	--14431
		x"ff",	--14432
		x"ff",	--14433
		x"ff",	--14434
		x"ff",	--14435
		x"ff",	--14436
		x"ff",	--14437
		x"ff",	--14438
		x"ff",	--14439
		x"ff",	--14440
		x"ff",	--14441
		x"ff",	--14442
		x"ff",	--14443
		x"ff",	--14444
		x"ff",	--14445
		x"ff",	--14446
		x"ff",	--14447
		x"ff",	--14448
		x"ff",	--14449
		x"ff",	--14450
		x"ff",	--14451
		x"ff",	--14452
		x"ff",	--14453
		x"ff",	--14454
		x"ff",	--14455
		x"ff",	--14456
		x"ff",	--14457
		x"ff",	--14458
		x"ff",	--14459
		x"ff",	--14460
		x"ff",	--14461
		x"ff",	--14462
		x"ff",	--14463
		x"ff",	--14464
		x"ff",	--14465
		x"ff",	--14466
		x"ff",	--14467
		x"ff",	--14468
		x"ff",	--14469
		x"ff",	--14470
		x"ff",	--14471
		x"ff",	--14472
		x"ff",	--14473
		x"ff",	--14474
		x"ff",	--14475
		x"ff",	--14476
		x"ff",	--14477
		x"ff",	--14478
		x"ff",	--14479
		x"ff",	--14480
		x"ff",	--14481
		x"ff",	--14482
		x"ff",	--14483
		x"ff",	--14484
		x"ff",	--14485
		x"ff",	--14486
		x"ff",	--14487
		x"ff",	--14488
		x"ff",	--14489
		x"ff",	--14490
		x"ff",	--14491
		x"ff",	--14492
		x"ff",	--14493
		x"ff",	--14494
		x"ff",	--14495
		x"ff",	--14496
		x"ff",	--14497
		x"ff",	--14498
		x"ff",	--14499
		x"ff",	--14500
		x"ff",	--14501
		x"ff",	--14502
		x"ff",	--14503
		x"ff",	--14504
		x"ff",	--14505
		x"ff",	--14506
		x"ff",	--14507
		x"ff",	--14508
		x"ff",	--14509
		x"ff",	--14510
		x"ff",	--14511
		x"ff",	--14512
		x"ff",	--14513
		x"ff",	--14514
		x"ff",	--14515
		x"ff",	--14516
		x"ff",	--14517
		x"ff",	--14518
		x"ff",	--14519
		x"ff",	--14520
		x"ff",	--14521
		x"ff",	--14522
		x"ff",	--14523
		x"ff",	--14524
		x"ff",	--14525
		x"ff",	--14526
		x"ff",	--14527
		x"ff",	--14528
		x"ff",	--14529
		x"ff",	--14530
		x"ff",	--14531
		x"ff",	--14532
		x"ff",	--14533
		x"ff",	--14534
		x"ff",	--14535
		x"ff",	--14536
		x"ff",	--14537
		x"ff",	--14538
		x"ff",	--14539
		x"ff",	--14540
		x"ff",	--14541
		x"ff",	--14542
		x"ff",	--14543
		x"ff",	--14544
		x"ff",	--14545
		x"ff",	--14546
		x"ff",	--14547
		x"ff",	--14548
		x"ff",	--14549
		x"ff",	--14550
		x"ff",	--14551
		x"ff",	--14552
		x"ff",	--14553
		x"ff",	--14554
		x"ff",	--14555
		x"ff",	--14556
		x"ff",	--14557
		x"ff",	--14558
		x"ff",	--14559
		x"ff",	--14560
		x"ff",	--14561
		x"ff",	--14562
		x"ff",	--14563
		x"ff",	--14564
		x"ff",	--14565
		x"ff",	--14566
		x"ff",	--14567
		x"ff",	--14568
		x"ff",	--14569
		x"ff",	--14570
		x"ff",	--14571
		x"ff",	--14572
		x"ff",	--14573
		x"ff",	--14574
		x"ff",	--14575
		x"ff",	--14576
		x"ff",	--14577
		x"ff",	--14578
		x"ff",	--14579
		x"ff",	--14580
		x"ff",	--14581
		x"ff",	--14582
		x"ff",	--14583
		x"ff",	--14584
		x"ff",	--14585
		x"ff",	--14586
		x"ff",	--14587
		x"ff",	--14588
		x"ff",	--14589
		x"ff",	--14590
		x"ff",	--14591
		x"ff",	--14592
		x"ff",	--14593
		x"ff",	--14594
		x"ff",	--14595
		x"ff",	--14596
		x"ff",	--14597
		x"ff",	--14598
		x"ff",	--14599
		x"ff",	--14600
		x"ff",	--14601
		x"ff",	--14602
		x"ff",	--14603
		x"ff",	--14604
		x"ff",	--14605
		x"ff",	--14606
		x"ff",	--14607
		x"ff",	--14608
		x"ff",	--14609
		x"ff",	--14610
		x"ff",	--14611
		x"ff",	--14612
		x"ff",	--14613
		x"ff",	--14614
		x"ff",	--14615
		x"ff",	--14616
		x"ff",	--14617
		x"ff",	--14618
		x"ff",	--14619
		x"ff",	--14620
		x"ff",	--14621
		x"ff",	--14622
		x"ff",	--14623
		x"ff",	--14624
		x"ff",	--14625
		x"ff",	--14626
		x"ff",	--14627
		x"ff",	--14628
		x"ff",	--14629
		x"ff",	--14630
		x"ff",	--14631
		x"ff",	--14632
		x"ff",	--14633
		x"ff",	--14634
		x"ff",	--14635
		x"ff",	--14636
		x"ff",	--14637
		x"ff",	--14638
		x"ff",	--14639
		x"ff",	--14640
		x"ff",	--14641
		x"ff",	--14642
		x"ff",	--14643
		x"ff",	--14644
		x"ff",	--14645
		x"ff",	--14646
		x"ff",	--14647
		x"ff",	--14648
		x"ff",	--14649
		x"ff",	--14650
		x"ff",	--14651
		x"ff",	--14652
		x"ff",	--14653
		x"ff",	--14654
		x"ff",	--14655
		x"ff",	--14656
		x"ff",	--14657
		x"ff",	--14658
		x"ff",	--14659
		x"ff",	--14660
		x"ff",	--14661
		x"ff",	--14662
		x"ff",	--14663
		x"ff",	--14664
		x"ff",	--14665
		x"ff",	--14666
		x"ff",	--14667
		x"ff",	--14668
		x"ff",	--14669
		x"ff",	--14670
		x"ff",	--14671
		x"ff",	--14672
		x"ff",	--14673
		x"ff",	--14674
		x"ff",	--14675
		x"ff",	--14676
		x"ff",	--14677
		x"ff",	--14678
		x"ff",	--14679
		x"ff",	--14680
		x"ff",	--14681
		x"ff",	--14682
		x"ff",	--14683
		x"ff",	--14684
		x"ff",	--14685
		x"ff",	--14686
		x"ff",	--14687
		x"ff",	--14688
		x"ff",	--14689
		x"ff",	--14690
		x"ff",	--14691
		x"ff",	--14692
		x"ff",	--14693
		x"ff",	--14694
		x"ff",	--14695
		x"ff",	--14696
		x"ff",	--14697
		x"ff",	--14698
		x"ff",	--14699
		x"ff",	--14700
		x"ff",	--14701
		x"ff",	--14702
		x"ff",	--14703
		x"ff",	--14704
		x"ff",	--14705
		x"ff",	--14706
		x"ff",	--14707
		x"ff",	--14708
		x"ff",	--14709
		x"ff",	--14710
		x"ff",	--14711
		x"ff",	--14712
		x"ff",	--14713
		x"ff",	--14714
		x"ff",	--14715
		x"ff",	--14716
		x"ff",	--14717
		x"ff",	--14718
		x"ff",	--14719
		x"ff",	--14720
		x"ff",	--14721
		x"ff",	--14722
		x"ff",	--14723
		x"ff",	--14724
		x"ff",	--14725
		x"ff",	--14726
		x"ff",	--14727
		x"ff",	--14728
		x"ff",	--14729
		x"ff",	--14730
		x"ff",	--14731
		x"ff",	--14732
		x"ff",	--14733
		x"ff",	--14734
		x"ff",	--14735
		x"ff",	--14736
		x"ff",	--14737
		x"ff",	--14738
		x"ff",	--14739
		x"ff",	--14740
		x"ff",	--14741
		x"ff",	--14742
		x"ff",	--14743
		x"ff",	--14744
		x"ff",	--14745
		x"ff",	--14746
		x"ff",	--14747
		x"ff",	--14748
		x"ff",	--14749
		x"ff",	--14750
		x"ff",	--14751
		x"ff",	--14752
		x"ff",	--14753
		x"ff",	--14754
		x"ff",	--14755
		x"ff",	--14756
		x"ff",	--14757
		x"ff",	--14758
		x"ff",	--14759
		x"ff",	--14760
		x"ff",	--14761
		x"ff",	--14762
		x"ff",	--14763
		x"ff",	--14764
		x"ff",	--14765
		x"ff",	--14766
		x"ff",	--14767
		x"ff",	--14768
		x"ff",	--14769
		x"ff",	--14770
		x"ff",	--14771
		x"ff",	--14772
		x"ff",	--14773
		x"ff",	--14774
		x"ff",	--14775
		x"ff",	--14776
		x"ff",	--14777
		x"ff",	--14778
		x"ff",	--14779
		x"ff",	--14780
		x"ff",	--14781
		x"ff",	--14782
		x"ff",	--14783
		x"ff",	--14784
		x"ff",	--14785
		x"ff",	--14786
		x"ff",	--14787
		x"ff",	--14788
		x"ff",	--14789
		x"ff",	--14790
		x"ff",	--14791
		x"ff",	--14792
		x"ff",	--14793
		x"ff",	--14794
		x"ff",	--14795
		x"ff",	--14796
		x"ff",	--14797
		x"ff",	--14798
		x"ff",	--14799
		x"ff",	--14800
		x"ff",	--14801
		x"ff",	--14802
		x"ff",	--14803
		x"ff",	--14804
		x"ff",	--14805
		x"ff",	--14806
		x"ff",	--14807
		x"ff",	--14808
		x"ff",	--14809
		x"ff",	--14810
		x"ff",	--14811
		x"ff",	--14812
		x"ff",	--14813
		x"ff",	--14814
		x"ff",	--14815
		x"ff",	--14816
		x"ff",	--14817
		x"ff",	--14818
		x"ff",	--14819
		x"ff",	--14820
		x"ff",	--14821
		x"ff",	--14822
		x"ff",	--14823
		x"ff",	--14824
		x"ff",	--14825
		x"ff",	--14826
		x"ff",	--14827
		x"ff",	--14828
		x"ff",	--14829
		x"ff",	--14830
		x"ff",	--14831
		x"ff",	--14832
		x"ff",	--14833
		x"ff",	--14834
		x"ff",	--14835
		x"ff",	--14836
		x"ff",	--14837
		x"ff",	--14838
		x"ff",	--14839
		x"ff",	--14840
		x"ff",	--14841
		x"ff",	--14842
		x"ff",	--14843
		x"ff",	--14844
		x"ff",	--14845
		x"ff",	--14846
		x"ff",	--14847
		x"ff",	--14848
		x"ff",	--14849
		x"ff",	--14850
		x"ff",	--14851
		x"ff",	--14852
		x"ff",	--14853
		x"ff",	--14854
		x"ff",	--14855
		x"ff",	--14856
		x"ff",	--14857
		x"ff",	--14858
		x"ff",	--14859
		x"ff",	--14860
		x"ff",	--14861
		x"ff",	--14862
		x"ff",	--14863
		x"ff",	--14864
		x"ff",	--14865
		x"ff",	--14866
		x"ff",	--14867
		x"ff",	--14868
		x"ff",	--14869
		x"ff",	--14870
		x"ff",	--14871
		x"ff",	--14872
		x"ff",	--14873
		x"ff",	--14874
		x"ff",	--14875
		x"ff",	--14876
		x"ff",	--14877
		x"ff",	--14878
		x"ff",	--14879
		x"ff",	--14880
		x"ff",	--14881
		x"ff",	--14882
		x"ff",	--14883
		x"ff",	--14884
		x"ff",	--14885
		x"ff",	--14886
		x"ff",	--14887
		x"ff",	--14888
		x"ff",	--14889
		x"ff",	--14890
		x"ff",	--14891
		x"ff",	--14892
		x"ff",	--14893
		x"ff",	--14894
		x"ff",	--14895
		x"ff",	--14896
		x"ff",	--14897
		x"ff",	--14898
		x"ff",	--14899
		x"ff",	--14900
		x"ff",	--14901
		x"ff",	--14902
		x"ff",	--14903
		x"ff",	--14904
		x"ff",	--14905
		x"ff",	--14906
		x"ff",	--14907
		x"ff",	--14908
		x"ff",	--14909
		x"ff",	--14910
		x"ff",	--14911
		x"ff",	--14912
		x"ff",	--14913
		x"ff",	--14914
		x"ff",	--14915
		x"ff",	--14916
		x"ff",	--14917
		x"ff",	--14918
		x"ff",	--14919
		x"ff",	--14920
		x"ff",	--14921
		x"ff",	--14922
		x"ff",	--14923
		x"ff",	--14924
		x"ff",	--14925
		x"ff",	--14926
		x"ff",	--14927
		x"ff",	--14928
		x"ff",	--14929
		x"ff",	--14930
		x"ff",	--14931
		x"ff",	--14932
		x"ff",	--14933
		x"ff",	--14934
		x"ff",	--14935
		x"ff",	--14936
		x"ff",	--14937
		x"ff",	--14938
		x"ff",	--14939
		x"ff",	--14940
		x"ff",	--14941
		x"ff",	--14942
		x"ff",	--14943
		x"ff",	--14944
		x"ff",	--14945
		x"ff",	--14946
		x"ff",	--14947
		x"ff",	--14948
		x"ff",	--14949
		x"ff",	--14950
		x"ff",	--14951
		x"ff",	--14952
		x"ff",	--14953
		x"ff",	--14954
		x"ff",	--14955
		x"ff",	--14956
		x"ff",	--14957
		x"ff",	--14958
		x"ff",	--14959
		x"ff",	--14960
		x"ff",	--14961
		x"ff",	--14962
		x"ff",	--14963
		x"ff",	--14964
		x"ff",	--14965
		x"ff",	--14966
		x"ff",	--14967
		x"ff",	--14968
		x"ff",	--14969
		x"ff",	--14970
		x"ff",	--14971
		x"ff",	--14972
		x"ff",	--14973
		x"ff",	--14974
		x"ff",	--14975
		x"ff",	--14976
		x"ff",	--14977
		x"ff",	--14978
		x"ff",	--14979
		x"ff",	--14980
		x"ff",	--14981
		x"ff",	--14982
		x"ff",	--14983
		x"ff",	--14984
		x"ff",	--14985
		x"ff",	--14986
		x"ff",	--14987
		x"ff",	--14988
		x"ff",	--14989
		x"ff",	--14990
		x"ff",	--14991
		x"ff",	--14992
		x"ff",	--14993
		x"ff",	--14994
		x"ff",	--14995
		x"ff",	--14996
		x"ff",	--14997
		x"ff",	--14998
		x"ff",	--14999
		x"ff",	--15000
		x"ff",	--15001
		x"ff",	--15002
		x"ff",	--15003
		x"ff",	--15004
		x"ff",	--15005
		x"ff",	--15006
		x"ff",	--15007
		x"ff",	--15008
		x"ff",	--15009
		x"ff",	--15010
		x"ff",	--15011
		x"ff",	--15012
		x"ff",	--15013
		x"ff",	--15014
		x"ff",	--15015
		x"ff",	--15016
		x"ff",	--15017
		x"ff",	--15018
		x"ff",	--15019
		x"ff",	--15020
		x"ff",	--15021
		x"ff",	--15022
		x"ff",	--15023
		x"ff",	--15024
		x"ff",	--15025
		x"ff",	--15026
		x"ff",	--15027
		x"ff",	--15028
		x"ff",	--15029
		x"ff",	--15030
		x"ff",	--15031
		x"ff",	--15032
		x"ff",	--15033
		x"ff",	--15034
		x"ff",	--15035
		x"ff",	--15036
		x"ff",	--15037
		x"ff",	--15038
		x"ff",	--15039
		x"ff",	--15040
		x"ff",	--15041
		x"ff",	--15042
		x"ff",	--15043
		x"ff",	--15044
		x"ff",	--15045
		x"ff",	--15046
		x"ff",	--15047
		x"ff",	--15048
		x"ff",	--15049
		x"ff",	--15050
		x"ff",	--15051
		x"ff",	--15052
		x"ff",	--15053
		x"ff",	--15054
		x"ff",	--15055
		x"ff",	--15056
		x"ff",	--15057
		x"ff",	--15058
		x"ff",	--15059
		x"ff",	--15060
		x"ff",	--15061
		x"ff",	--15062
		x"ff",	--15063
		x"ff",	--15064
		x"ff",	--15065
		x"ff",	--15066
		x"ff",	--15067
		x"ff",	--15068
		x"ff",	--15069
		x"ff",	--15070
		x"ff",	--15071
		x"ff",	--15072
		x"ff",	--15073
		x"ff",	--15074
		x"ff",	--15075
		x"ff",	--15076
		x"ff",	--15077
		x"ff",	--15078
		x"ff",	--15079
		x"ff",	--15080
		x"ff",	--15081
		x"ff",	--15082
		x"ff",	--15083
		x"ff",	--15084
		x"ff",	--15085
		x"ff",	--15086
		x"ff",	--15087
		x"ff",	--15088
		x"ff",	--15089
		x"ff",	--15090
		x"ff",	--15091
		x"ff",	--15092
		x"ff",	--15093
		x"ff",	--15094
		x"ff",	--15095
		x"ff",	--15096
		x"ff",	--15097
		x"ff",	--15098
		x"ff",	--15099
		x"ff",	--15100
		x"ff",	--15101
		x"ff",	--15102
		x"ff",	--15103
		x"ff",	--15104
		x"ff",	--15105
		x"ff",	--15106
		x"ff",	--15107
		x"ff",	--15108
		x"ff",	--15109
		x"ff",	--15110
		x"ff",	--15111
		x"ff",	--15112
		x"ff",	--15113
		x"ff",	--15114
		x"ff",	--15115
		x"ff",	--15116
		x"ff",	--15117
		x"ff",	--15118
		x"ff",	--15119
		x"ff",	--15120
		x"ff",	--15121
		x"ff",	--15122
		x"ff",	--15123
		x"ff",	--15124
		x"ff",	--15125
		x"ff",	--15126
		x"ff",	--15127
		x"ff",	--15128
		x"ff",	--15129
		x"ff",	--15130
		x"ff",	--15131
		x"ff",	--15132
		x"ff",	--15133
		x"ff",	--15134
		x"ff",	--15135
		x"ff",	--15136
		x"ff",	--15137
		x"ff",	--15138
		x"ff",	--15139
		x"ff",	--15140
		x"ff",	--15141
		x"ff",	--15142
		x"ff",	--15143
		x"ff",	--15144
		x"ff",	--15145
		x"ff",	--15146
		x"ff",	--15147
		x"ff",	--15148
		x"ff",	--15149
		x"ff",	--15150
		x"ff",	--15151
		x"ff",	--15152
		x"ff",	--15153
		x"ff",	--15154
		x"ff",	--15155
		x"ff",	--15156
		x"ff",	--15157
		x"ff",	--15158
		x"ff",	--15159
		x"ff",	--15160
		x"ff",	--15161
		x"ff",	--15162
		x"ff",	--15163
		x"ff",	--15164
		x"ff",	--15165
		x"ff",	--15166
		x"ff",	--15167
		x"ff",	--15168
		x"ff",	--15169
		x"ff",	--15170
		x"ff",	--15171
		x"ff",	--15172
		x"ff",	--15173
		x"ff",	--15174
		x"ff",	--15175
		x"ff",	--15176
		x"ff",	--15177
		x"ff",	--15178
		x"ff",	--15179
		x"ff",	--15180
		x"ff",	--15181
		x"ff",	--15182
		x"ff",	--15183
		x"ff",	--15184
		x"ff",	--15185
		x"ff",	--15186
		x"ff",	--15187
		x"ff",	--15188
		x"ff",	--15189
		x"ff",	--15190
		x"ff",	--15191
		x"ff",	--15192
		x"ff",	--15193
		x"ff",	--15194
		x"ff",	--15195
		x"ff",	--15196
		x"ff",	--15197
		x"ff",	--15198
		x"ff",	--15199
		x"ff",	--15200
		x"ff",	--15201
		x"ff",	--15202
		x"ff",	--15203
		x"ff",	--15204
		x"ff",	--15205
		x"ff",	--15206
		x"ff",	--15207
		x"ff",	--15208
		x"ff",	--15209
		x"ff",	--15210
		x"ff",	--15211
		x"ff",	--15212
		x"ff",	--15213
		x"ff",	--15214
		x"ff",	--15215
		x"ff",	--15216
		x"ff",	--15217
		x"ff",	--15218
		x"ff",	--15219
		x"ff",	--15220
		x"ff",	--15221
		x"ff",	--15222
		x"ff",	--15223
		x"ff",	--15224
		x"ff",	--15225
		x"ff",	--15226
		x"ff",	--15227
		x"ff",	--15228
		x"ff",	--15229
		x"ff",	--15230
		x"ff",	--15231
		x"ff",	--15232
		x"ff",	--15233
		x"ff",	--15234
		x"ff",	--15235
		x"ff",	--15236
		x"ff",	--15237
		x"ff",	--15238
		x"ff",	--15239
		x"ff",	--15240
		x"ff",	--15241
		x"ff",	--15242
		x"ff",	--15243
		x"ff",	--15244
		x"ff",	--15245
		x"ff",	--15246
		x"ff",	--15247
		x"ff",	--15248
		x"ff",	--15249
		x"ff",	--15250
		x"ff",	--15251
		x"ff",	--15252
		x"ff",	--15253
		x"ff",	--15254
		x"ff",	--15255
		x"ff",	--15256
		x"ff",	--15257
		x"ff",	--15258
		x"ff",	--15259
		x"ff",	--15260
		x"ff",	--15261
		x"ff",	--15262
		x"ff",	--15263
		x"ff",	--15264
		x"ff",	--15265
		x"ff",	--15266
		x"ff",	--15267
		x"ff",	--15268
		x"ff",	--15269
		x"ff",	--15270
		x"ff",	--15271
		x"ff",	--15272
		x"ff",	--15273
		x"ff",	--15274
		x"ff",	--15275
		x"ff",	--15276
		x"ff",	--15277
		x"ff",	--15278
		x"ff",	--15279
		x"ff",	--15280
		x"ff",	--15281
		x"ff",	--15282
		x"ff",	--15283
		x"ff",	--15284
		x"ff",	--15285
		x"ff",	--15286
		x"ff",	--15287
		x"ff",	--15288
		x"ff",	--15289
		x"ff",	--15290
		x"ff",	--15291
		x"ff",	--15292
		x"ff",	--15293
		x"ff",	--15294
		x"ff",	--15295
		x"ff",	--15296
		x"ff",	--15297
		x"ff",	--15298
		x"ff",	--15299
		x"ff",	--15300
		x"ff",	--15301
		x"ff",	--15302
		x"ff",	--15303
		x"ff",	--15304
		x"ff",	--15305
		x"ff",	--15306
		x"ff",	--15307
		x"ff",	--15308
		x"ff",	--15309
		x"ff",	--15310
		x"ff",	--15311
		x"ff",	--15312
		x"ff",	--15313
		x"ff",	--15314
		x"ff",	--15315
		x"ff",	--15316
		x"ff",	--15317
		x"ff",	--15318
		x"ff",	--15319
		x"ff",	--15320
		x"ff",	--15321
		x"ff",	--15322
		x"ff",	--15323
		x"ff",	--15324
		x"ff",	--15325
		x"ff",	--15326
		x"ff",	--15327
		x"ff",	--15328
		x"ff",	--15329
		x"ff",	--15330
		x"ff",	--15331
		x"ff",	--15332
		x"ff",	--15333
		x"ff",	--15334
		x"ff",	--15335
		x"ff",	--15336
		x"ff",	--15337
		x"ff",	--15338
		x"ff",	--15339
		x"ff",	--15340
		x"ff",	--15341
		x"ff",	--15342
		x"ff",	--15343
		x"ff",	--15344
		x"ff",	--15345
		x"ff",	--15346
		x"ff",	--15347
		x"ff",	--15348
		x"ff",	--15349
		x"ff",	--15350
		x"ff",	--15351
		x"ff",	--15352
		x"ff",	--15353
		x"ff",	--15354
		x"ff",	--15355
		x"ff",	--15356
		x"ff",	--15357
		x"ff",	--15358
		x"ff",	--15359
		x"ff",	--15360
		x"ff",	--15361
		x"ff",	--15362
		x"ff",	--15363
		x"ff",	--15364
		x"ff",	--15365
		x"ff",	--15366
		x"ff",	--15367
		x"ff",	--15368
		x"ff",	--15369
		x"ff",	--15370
		x"ff",	--15371
		x"ff",	--15372
		x"ff",	--15373
		x"ff",	--15374
		x"ff",	--15375
		x"ff",	--15376
		x"ff",	--15377
		x"ff",	--15378
		x"ff",	--15379
		x"ff",	--15380
		x"ff",	--15381
		x"ff",	--15382
		x"ff",	--15383
		x"ff",	--15384
		x"ff",	--15385
		x"ff",	--15386
		x"ff",	--15387
		x"ff",	--15388
		x"ff",	--15389
		x"ff",	--15390
		x"ff",	--15391
		x"ff",	--15392
		x"ff",	--15393
		x"ff",	--15394
		x"ff",	--15395
		x"ff",	--15396
		x"ff",	--15397
		x"ff",	--15398
		x"ff",	--15399
		x"ff",	--15400
		x"ff",	--15401
		x"ff",	--15402
		x"ff",	--15403
		x"ff",	--15404
		x"ff",	--15405
		x"ff",	--15406
		x"ff",	--15407
		x"ff",	--15408
		x"ff",	--15409
		x"ff",	--15410
		x"ff",	--15411
		x"ff",	--15412
		x"ff",	--15413
		x"ff",	--15414
		x"ff",	--15415
		x"ff",	--15416
		x"ff",	--15417
		x"ff",	--15418
		x"ff",	--15419
		x"ff",	--15420
		x"ff",	--15421
		x"ff",	--15422
		x"ff",	--15423
		x"ff",	--15424
		x"ff",	--15425
		x"ff",	--15426
		x"ff",	--15427
		x"ff",	--15428
		x"ff",	--15429
		x"ff",	--15430
		x"ff",	--15431
		x"ff",	--15432
		x"ff",	--15433
		x"ff",	--15434
		x"ff",	--15435
		x"ff",	--15436
		x"ff",	--15437
		x"ff",	--15438
		x"ff",	--15439
		x"ff",	--15440
		x"ff",	--15441
		x"ff",	--15442
		x"ff",	--15443
		x"ff",	--15444
		x"ff",	--15445
		x"ff",	--15446
		x"ff",	--15447
		x"ff",	--15448
		x"ff",	--15449
		x"ff",	--15450
		x"ff",	--15451
		x"ff",	--15452
		x"ff",	--15453
		x"ff",	--15454
		x"ff",	--15455
		x"ff",	--15456
		x"ff",	--15457
		x"ff",	--15458
		x"ff",	--15459
		x"ff",	--15460
		x"ff",	--15461
		x"ff",	--15462
		x"ff",	--15463
		x"ff",	--15464
		x"ff",	--15465
		x"ff",	--15466
		x"ff",	--15467
		x"ff",	--15468
		x"ff",	--15469
		x"ff",	--15470
		x"ff",	--15471
		x"ff",	--15472
		x"ff",	--15473
		x"ff",	--15474
		x"ff",	--15475
		x"ff",	--15476
		x"ff",	--15477
		x"ff",	--15478
		x"ff",	--15479
		x"ff",	--15480
		x"ff",	--15481
		x"ff",	--15482
		x"ff",	--15483
		x"ff",	--15484
		x"ff",	--15485
		x"ff",	--15486
		x"ff",	--15487
		x"ff",	--15488
		x"ff",	--15489
		x"ff",	--15490
		x"ff",	--15491
		x"ff",	--15492
		x"ff",	--15493
		x"ff",	--15494
		x"ff",	--15495
		x"ff",	--15496
		x"ff",	--15497
		x"ff",	--15498
		x"ff",	--15499
		x"ff",	--15500
		x"ff",	--15501
		x"ff",	--15502
		x"ff",	--15503
		x"ff",	--15504
		x"ff",	--15505
		x"ff",	--15506
		x"ff",	--15507
		x"ff",	--15508
		x"ff",	--15509
		x"ff",	--15510
		x"ff",	--15511
		x"ff",	--15512
		x"ff",	--15513
		x"ff",	--15514
		x"ff",	--15515
		x"ff",	--15516
		x"ff",	--15517
		x"ff",	--15518
		x"ff",	--15519
		x"ff",	--15520
		x"ff",	--15521
		x"ff",	--15522
		x"ff",	--15523
		x"ff",	--15524
		x"ff",	--15525
		x"ff",	--15526
		x"ff",	--15527
		x"ff",	--15528
		x"ff",	--15529
		x"ff",	--15530
		x"ff",	--15531
		x"ff",	--15532
		x"ff",	--15533
		x"ff",	--15534
		x"ff",	--15535
		x"ff",	--15536
		x"ff",	--15537
		x"ff",	--15538
		x"ff",	--15539
		x"ff",	--15540
		x"ff",	--15541
		x"ff",	--15542
		x"ff",	--15543
		x"ff",	--15544
		x"ff",	--15545
		x"ff",	--15546
		x"ff",	--15547
		x"ff",	--15548
		x"ff",	--15549
		x"ff",	--15550
		x"ff",	--15551
		x"ff",	--15552
		x"ff",	--15553
		x"ff",	--15554
		x"ff",	--15555
		x"ff",	--15556
		x"ff",	--15557
		x"ff",	--15558
		x"ff",	--15559
		x"ff",	--15560
		x"ff",	--15561
		x"ff",	--15562
		x"ff",	--15563
		x"ff",	--15564
		x"ff",	--15565
		x"ff",	--15566
		x"ff",	--15567
		x"ff",	--15568
		x"ff",	--15569
		x"ff",	--15570
		x"ff",	--15571
		x"ff",	--15572
		x"ff",	--15573
		x"ff",	--15574
		x"ff",	--15575
		x"ff",	--15576
		x"ff",	--15577
		x"ff",	--15578
		x"ff",	--15579
		x"ff",	--15580
		x"ff",	--15581
		x"ff",	--15582
		x"ff",	--15583
		x"ff",	--15584
		x"ff",	--15585
		x"ff",	--15586
		x"ff",	--15587
		x"ff",	--15588
		x"ff",	--15589
		x"ff",	--15590
		x"ff",	--15591
		x"ff",	--15592
		x"ff",	--15593
		x"ff",	--15594
		x"ff",	--15595
		x"ff",	--15596
		x"ff",	--15597
		x"ff",	--15598
		x"ff",	--15599
		x"ff",	--15600
		x"ff",	--15601
		x"ff",	--15602
		x"ff",	--15603
		x"ff",	--15604
		x"ff",	--15605
		x"ff",	--15606
		x"ff",	--15607
		x"ff",	--15608
		x"ff",	--15609
		x"ff",	--15610
		x"ff",	--15611
		x"ff",	--15612
		x"ff",	--15613
		x"ff",	--15614
		x"ff",	--15615
		x"ff",	--15616
		x"ff",	--15617
		x"ff",	--15618
		x"ff",	--15619
		x"ff",	--15620
		x"ff",	--15621
		x"ff",	--15622
		x"ff",	--15623
		x"ff",	--15624
		x"ff",	--15625
		x"ff",	--15626
		x"ff",	--15627
		x"ff",	--15628
		x"ff",	--15629
		x"ff",	--15630
		x"ff",	--15631
		x"ff",	--15632
		x"ff",	--15633
		x"ff",	--15634
		x"ff",	--15635
		x"ff",	--15636
		x"ff",	--15637
		x"ff",	--15638
		x"ff",	--15639
		x"ff",	--15640
		x"ff",	--15641
		x"ff",	--15642
		x"ff",	--15643
		x"ff",	--15644
		x"ff",	--15645
		x"ff",	--15646
		x"ff",	--15647
		x"ff",	--15648
		x"ff",	--15649
		x"ff",	--15650
		x"ff",	--15651
		x"ff",	--15652
		x"ff",	--15653
		x"ff",	--15654
		x"ff",	--15655
		x"ff",	--15656
		x"ff",	--15657
		x"ff",	--15658
		x"ff",	--15659
		x"ff",	--15660
		x"ff",	--15661
		x"ff",	--15662
		x"ff",	--15663
		x"ff",	--15664
		x"ff",	--15665
		x"ff",	--15666
		x"ff",	--15667
		x"ff",	--15668
		x"ff",	--15669
		x"ff",	--15670
		x"ff",	--15671
		x"ff",	--15672
		x"ff",	--15673
		x"ff",	--15674
		x"ff",	--15675
		x"ff",	--15676
		x"ff",	--15677
		x"ff",	--15678
		x"ff",	--15679
		x"ff",	--15680
		x"ff",	--15681
		x"ff",	--15682
		x"ff",	--15683
		x"ff",	--15684
		x"ff",	--15685
		x"ff",	--15686
		x"ff",	--15687
		x"ff",	--15688
		x"ff",	--15689
		x"ff",	--15690
		x"ff",	--15691
		x"ff",	--15692
		x"ff",	--15693
		x"ff",	--15694
		x"ff",	--15695
		x"ff",	--15696
		x"ff",	--15697
		x"ff",	--15698
		x"ff",	--15699
		x"ff",	--15700
		x"ff",	--15701
		x"ff",	--15702
		x"ff",	--15703
		x"ff",	--15704
		x"ff",	--15705
		x"ff",	--15706
		x"ff",	--15707
		x"ff",	--15708
		x"ff",	--15709
		x"ff",	--15710
		x"ff",	--15711
		x"ff",	--15712
		x"ff",	--15713
		x"ff",	--15714
		x"ff",	--15715
		x"ff",	--15716
		x"ff",	--15717
		x"ff",	--15718
		x"ff",	--15719
		x"ff",	--15720
		x"ff",	--15721
		x"ff",	--15722
		x"ff",	--15723
		x"ff",	--15724
		x"ff",	--15725
		x"ff",	--15726
		x"ff",	--15727
		x"ff",	--15728
		x"ff",	--15729
		x"ff",	--15730
		x"ff",	--15731
		x"ff",	--15732
		x"ff",	--15733
		x"ff",	--15734
		x"ff",	--15735
		x"ff",	--15736
		x"ff",	--15737
		x"ff",	--15738
		x"ff",	--15739
		x"ff",	--15740
		x"ff",	--15741
		x"ff",	--15742
		x"ff",	--15743
		x"ff",	--15744
		x"ff",	--15745
		x"ff",	--15746
		x"ff",	--15747
		x"ff",	--15748
		x"ff",	--15749
		x"ff",	--15750
		x"ff",	--15751
		x"ff",	--15752
		x"ff",	--15753
		x"ff",	--15754
		x"ff",	--15755
		x"ff",	--15756
		x"ff",	--15757
		x"ff",	--15758
		x"ff",	--15759
		x"ff",	--15760
		x"ff",	--15761
		x"ff",	--15762
		x"ff",	--15763
		x"ff",	--15764
		x"ff",	--15765
		x"ff",	--15766
		x"ff",	--15767
		x"ff",	--15768
		x"ff",	--15769
		x"ff",	--15770
		x"ff",	--15771
		x"ff",	--15772
		x"ff",	--15773
		x"ff",	--15774
		x"ff",	--15775
		x"ff",	--15776
		x"ff",	--15777
		x"ff",	--15778
		x"ff",	--15779
		x"ff",	--15780
		x"ff",	--15781
		x"ff",	--15782
		x"ff",	--15783
		x"ff",	--15784
		x"ff",	--15785
		x"ff",	--15786
		x"ff",	--15787
		x"ff",	--15788
		x"ff",	--15789
		x"ff",	--15790
		x"ff",	--15791
		x"ff",	--15792
		x"ff",	--15793
		x"ff",	--15794
		x"ff",	--15795
		x"ff",	--15796
		x"ff",	--15797
		x"ff",	--15798
		x"ff",	--15799
		x"ff",	--15800
		x"ff",	--15801
		x"ff",	--15802
		x"ff",	--15803
		x"ff",	--15804
		x"ff",	--15805
		x"ff",	--15806
		x"ff",	--15807
		x"ff",	--15808
		x"ff",	--15809
		x"ff",	--15810
		x"ff",	--15811
		x"ff",	--15812
		x"ff",	--15813
		x"ff",	--15814
		x"ff",	--15815
		x"ff",	--15816
		x"ff",	--15817
		x"ff",	--15818
		x"ff",	--15819
		x"ff",	--15820
		x"ff",	--15821
		x"ff",	--15822
		x"ff",	--15823
		x"ff",	--15824
		x"ff",	--15825
		x"ff",	--15826
		x"ff",	--15827
		x"ff",	--15828
		x"ff",	--15829
		x"ff",	--15830
		x"ff",	--15831
		x"ff",	--15832
		x"ff",	--15833
		x"ff",	--15834
		x"ff",	--15835
		x"ff",	--15836
		x"ff",	--15837
		x"ff",	--15838
		x"ff",	--15839
		x"ff",	--15840
		x"ff",	--15841
		x"ff",	--15842
		x"ff",	--15843
		x"ff",	--15844
		x"ff",	--15845
		x"ff",	--15846
		x"ff",	--15847
		x"ff",	--15848
		x"ff",	--15849
		x"ff",	--15850
		x"ff",	--15851
		x"ff",	--15852
		x"ff",	--15853
		x"ff",	--15854
		x"ff",	--15855
		x"ff",	--15856
		x"ff",	--15857
		x"ff",	--15858
		x"ff",	--15859
		x"ff",	--15860
		x"ff",	--15861
		x"ff",	--15862
		x"ff",	--15863
		x"ff",	--15864
		x"ff",	--15865
		x"ff",	--15866
		x"ff",	--15867
		x"ff",	--15868
		x"ff",	--15869
		x"ff",	--15870
		x"ff",	--15871
		x"ff",	--15872
		x"ff",	--15873
		x"ff",	--15874
		x"ff",	--15875
		x"ff",	--15876
		x"ff",	--15877
		x"ff",	--15878
		x"ff",	--15879
		x"ff",	--15880
		x"ff",	--15881
		x"ff",	--15882
		x"ff",	--15883
		x"ff",	--15884
		x"ff",	--15885
		x"ff",	--15886
		x"ff",	--15887
		x"ff",	--15888
		x"ff",	--15889
		x"ff",	--15890
		x"ff",	--15891
		x"ff",	--15892
		x"ff",	--15893
		x"ff",	--15894
		x"ff",	--15895
		x"ff",	--15896
		x"ff",	--15897
		x"ff",	--15898
		x"ff",	--15899
		x"ff",	--15900
		x"ff",	--15901
		x"ff",	--15902
		x"ff",	--15903
		x"ff",	--15904
		x"ff",	--15905
		x"ff",	--15906
		x"ff",	--15907
		x"ff",	--15908
		x"ff",	--15909
		x"ff",	--15910
		x"ff",	--15911
		x"ff",	--15912
		x"ff",	--15913
		x"ff",	--15914
		x"ff",	--15915
		x"ff",	--15916
		x"ff",	--15917
		x"ff",	--15918
		x"ff",	--15919
		x"ff",	--15920
		x"ff",	--15921
		x"ff",	--15922
		x"ff",	--15923
		x"ff",	--15924
		x"ff",	--15925
		x"ff",	--15926
		x"ff",	--15927
		x"ff",	--15928
		x"ff",	--15929
		x"ff",	--15930
		x"ff",	--15931
		x"ff",	--15932
		x"ff",	--15933
		x"ff",	--15934
		x"ff",	--15935
		x"ff",	--15936
		x"ff",	--15937
		x"ff",	--15938
		x"ff",	--15939
		x"ff",	--15940
		x"ff",	--15941
		x"ff",	--15942
		x"ff",	--15943
		x"ff",	--15944
		x"ff",	--15945
		x"ff",	--15946
		x"ff",	--15947
		x"ff",	--15948
		x"ff",	--15949
		x"ff",	--15950
		x"ff",	--15951
		x"ff",	--15952
		x"ff",	--15953
		x"ff",	--15954
		x"ff",	--15955
		x"ff",	--15956
		x"ff",	--15957
		x"ff",	--15958
		x"ff",	--15959
		x"ff",	--15960
		x"ff",	--15961
		x"ff",	--15962
		x"ff",	--15963
		x"ff",	--15964
		x"ff",	--15965
		x"ff",	--15966
		x"ff",	--15967
		x"ff",	--15968
		x"ff",	--15969
		x"ff",	--15970
		x"ff",	--15971
		x"ff",	--15972
		x"ff",	--15973
		x"ff",	--15974
		x"ff",	--15975
		x"ff",	--15976
		x"ff",	--15977
		x"ff",	--15978
		x"ff",	--15979
		x"ff",	--15980
		x"ff",	--15981
		x"ff",	--15982
		x"ff",	--15983
		x"ff",	--15984
		x"ff",	--15985
		x"ff",	--15986
		x"ff",	--15987
		x"ff",	--15988
		x"ff",	--15989
		x"ff",	--15990
		x"ff",	--15991
		x"ff",	--15992
		x"ff",	--15993
		x"ff",	--15994
		x"ff",	--15995
		x"ff",	--15996
		x"ff",	--15997
		x"ff",	--15998
		x"ff",	--15999
		x"ff",	--16000
		x"ff",	--16001
		x"ff",	--16002
		x"ff",	--16003
		x"ff",	--16004
		x"ff",	--16005
		x"ff",	--16006
		x"ff",	--16007
		x"ff",	--16008
		x"ff",	--16009
		x"ff",	--16010
		x"ff",	--16011
		x"ff",	--16012
		x"ff",	--16013
		x"ff",	--16014
		x"ff",	--16015
		x"ff",	--16016
		x"ff",	--16017
		x"ff",	--16018
		x"ff",	--16019
		x"ff",	--16020
		x"ff",	--16021
		x"ff",	--16022
		x"ff",	--16023
		x"ff",	--16024
		x"ff",	--16025
		x"ff",	--16026
		x"ff",	--16027
		x"ff",	--16028
		x"ff",	--16029
		x"ff",	--16030
		x"ff",	--16031
		x"ff",	--16032
		x"ff",	--16033
		x"ff",	--16034
		x"ff",	--16035
		x"ff",	--16036
		x"ff",	--16037
		x"ff",	--16038
		x"ff",	--16039
		x"ff",	--16040
		x"ff",	--16041
		x"ff",	--16042
		x"ff",	--16043
		x"ff",	--16044
		x"ff",	--16045
		x"ff",	--16046
		x"ff",	--16047
		x"ff",	--16048
		x"ff",	--16049
		x"ff",	--16050
		x"ff",	--16051
		x"ff",	--16052
		x"ff",	--16053
		x"ff",	--16054
		x"ff",	--16055
		x"ff",	--16056
		x"ff",	--16057
		x"ff",	--16058
		x"ff",	--16059
		x"ff",	--16060
		x"ff",	--16061
		x"ff",	--16062
		x"ff",	--16063
		x"ff",	--16064
		x"ff",	--16065
		x"ff",	--16066
		x"ff",	--16067
		x"ff",	--16068
		x"ff",	--16069
		x"ff",	--16070
		x"ff",	--16071
		x"ff",	--16072
		x"ff",	--16073
		x"ff",	--16074
		x"ff",	--16075
		x"ff",	--16076
		x"ff",	--16077
		x"ff",	--16078
		x"ff",	--16079
		x"ff",	--16080
		x"ff",	--16081
		x"ff",	--16082
		x"ff",	--16083
		x"ff",	--16084
		x"ff",	--16085
		x"ff",	--16086
		x"ff",	--16087
		x"ff",	--16088
		x"ff",	--16089
		x"ff",	--16090
		x"ff",	--16091
		x"ff",	--16092
		x"ff",	--16093
		x"ff",	--16094
		x"ff",	--16095
		x"ff",	--16096
		x"ff",	--16097
		x"ff",	--16098
		x"ff",	--16099
		x"ff",	--16100
		x"ff",	--16101
		x"ff",	--16102
		x"ff",	--16103
		x"ff",	--16104
		x"ff",	--16105
		x"ff",	--16106
		x"ff",	--16107
		x"ff",	--16108
		x"ff",	--16109
		x"ff",	--16110
		x"ff",	--16111
		x"ff",	--16112
		x"ff",	--16113
		x"ff",	--16114
		x"ff",	--16115
		x"ff",	--16116
		x"ff",	--16117
		x"ff",	--16118
		x"ff",	--16119
		x"ff",	--16120
		x"ff",	--16121
		x"ff",	--16122
		x"ff",	--16123
		x"ff",	--16124
		x"ff",	--16125
		x"ff",	--16126
		x"ff",	--16127
		x"ff",	--16128
		x"ff",	--16129
		x"ff",	--16130
		x"ff",	--16131
		x"ff",	--16132
		x"ff",	--16133
		x"ff",	--16134
		x"ff",	--16135
		x"ff",	--16136
		x"ff",	--16137
		x"ff",	--16138
		x"ff",	--16139
		x"ff",	--16140
		x"ff",	--16141
		x"ff",	--16142
		x"ff",	--16143
		x"ff",	--16144
		x"ff",	--16145
		x"ff",	--16146
		x"ff",	--16147
		x"ff",	--16148
		x"ff",	--16149
		x"ff",	--16150
		x"ff",	--16151
		x"ff",	--16152
		x"ff",	--16153
		x"ff",	--16154
		x"ff",	--16155
		x"ff",	--16156
		x"ff",	--16157
		x"ff",	--16158
		x"ff",	--16159
		x"ff",	--16160
		x"ff",	--16161
		x"ff",	--16162
		x"ff",	--16163
		x"ff",	--16164
		x"ff",	--16165
		x"ff",	--16166
		x"ff",	--16167
		x"ff",	--16168
		x"ff",	--16169
		x"ff",	--16170
		x"ff",	--16171
		x"ff",	--16172
		x"ff",	--16173
		x"ff",	--16174
		x"ff",	--16175
		x"ff",	--16176
		x"ff",	--16177
		x"ff",	--16178
		x"ff",	--16179
		x"ff",	--16180
		x"ff",	--16181
		x"ff",	--16182
		x"ff",	--16183
		x"ff",	--16184
		x"ff",	--16185
		x"ff",	--16186
		x"ff",	--16187
		x"ff",	--16188
		x"ff",	--16189
		x"ff",	--16190
		x"ff",	--16191
		x"ff",	--16192
		x"ff",	--16193
		x"ff",	--16194
		x"ff",	--16195
		x"ff",	--16196
		x"ff",	--16197
		x"ff",	--16198
		x"ff",	--16199
		x"ff",	--16200
		x"ff",	--16201
		x"ff",	--16202
		x"ff",	--16203
		x"ff",	--16204
		x"ff",	--16205
		x"ff",	--16206
		x"ff",	--16207
		x"ff",	--16208
		x"ff",	--16209
		x"ff",	--16210
		x"ff",	--16211
		x"ff",	--16212
		x"ff",	--16213
		x"ff",	--16214
		x"ff",	--16215
		x"ff",	--16216
		x"ff",	--16217
		x"ff",	--16218
		x"ff",	--16219
		x"ff",	--16220
		x"ff",	--16221
		x"ff",	--16222
		x"ff",	--16223
		x"ff",	--16224
		x"ff",	--16225
		x"ff",	--16226
		x"ff",	--16227
		x"ff",	--16228
		x"ff",	--16229
		x"ff",	--16230
		x"ff",	--16231
		x"ff",	--16232
		x"ff",	--16233
		x"ff",	--16234
		x"ff",	--16235
		x"ff",	--16236
		x"ff",	--16237
		x"ff",	--16238
		x"ff",	--16239
		x"ff",	--16240
		x"ff",	--16241
		x"ff",	--16242
		x"ff",	--16243
		x"ff",	--16244
		x"ff",	--16245
		x"ff",	--16246
		x"ff",	--16247
		x"ff",	--16248
		x"ff",	--16249
		x"ff",	--16250
		x"ff",	--16251
		x"ff",	--16252
		x"ff",	--16253
		x"ff",	--16254
		x"ff",	--16255
		x"ff",	--16256
		x"ff",	--16257
		x"ff",	--16258
		x"ff",	--16259
		x"ff",	--16260
		x"ff",	--16261
		x"ff",	--16262
		x"ff",	--16263
		x"ff",	--16264
		x"ff",	--16265
		x"ff",	--16266
		x"ff",	--16267
		x"ff",	--16268
		x"ff",	--16269
		x"ff",	--16270
		x"ff",	--16271
		x"ff",	--16272
		x"ff",	--16273
		x"ff",	--16274
		x"ff",	--16275
		x"ff",	--16276
		x"ff",	--16277
		x"ff",	--16278
		x"ff",	--16279
		x"ff",	--16280
		x"ff",	--16281
		x"ff",	--16282
		x"ff",	--16283
		x"ff",	--16284
		x"ff",	--16285
		x"ff",	--16286
		x"ff",	--16287
		x"ff",	--16288
		x"ff",	--16289
		x"ff",	--16290
		x"ff",	--16291
		x"ff",	--16292
		x"ff",	--16293
		x"ff",	--16294
		x"ff",	--16295
		x"ff",	--16296
		x"ff",	--16297
		x"ff",	--16298
		x"ff",	--16299
		x"ff",	--16300
		x"ff",	--16301
		x"ff",	--16302
		x"ff",	--16303
		x"ff",	--16304
		x"ff",	--16305
		x"ff",	--16306
		x"ff",	--16307
		x"ff",	--16308
		x"ff",	--16309
		x"ff",	--16310
		x"ff",	--16311
		x"ff",	--16312
		x"ff",	--16313
		x"ff",	--16314
		x"ff",	--16315
		x"ff",	--16316
		x"ff",	--16317
		x"ff",	--16318
		x"ff",	--16319
		x"ff",	--16320
		x"ff",	--16321
		x"ff",	--16322
		x"ff",	--16323
		x"ff",	--16324
		x"ff",	--16325
		x"ff",	--16326
		x"ff",	--16327
		x"ff",	--16328
		x"ff",	--16329
		x"ff",	--16330
		x"ff",	--16331
		x"ff",	--16332
		x"ff",	--16333
		x"ff",	--16334
		x"ff",	--16335
		x"ff",	--16336
		x"ff",	--16337
		x"ff",	--16338
		x"ff",	--16339
		x"ff",	--16340
		x"ff",	--16341
		x"ff",	--16342
		x"ff",	--16343
		x"ff",	--16344
		x"ff",	--16345
		x"ff",	--16346
		x"ff",	--16347
		x"ff",	--16348
		x"ff",	--16349
		x"ff",	--16350
		x"ff",	--16351
		x"ff",	--16352
		x"ff",	--16353
		x"ff",	--16354
		x"ff",	--16355
		x"ff",	--16356
		x"ff",	--16357
		x"ff",	--16358
		x"ff",	--16359
		x"ff",	--16360
		x"ff",	--16361
		x"ff",	--16362
		x"ff",	--16363
		x"ff",	--16364
		x"ff",	--16365
		x"ff",	--16366
		x"ff",	--16367
		x"83",	--16368
		x"83",	--16369
		x"83",	--16370
		x"83",	--16371
		x"83",	--16372
		x"83",	--16373
		x"83",	--16374
		x"9d",	--16375
		x"99",	--16376
		x"83",	--16377
		x"83",	--16378
		x"83",	--16379
		x"83",	--16380
		x"83",	--16381
		x"83",	--16382
		x"80");	--16383

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
