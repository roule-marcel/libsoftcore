library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"4a",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"00",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"4a",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"62",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"4a",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"4a",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"00",	--29
		x"f9",	--30
		x"31",	--31
		x"c2",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"80",	--41
		x"0f",	--42
		x"b0",	--43
		x"4a",	--44
		x"b0",	--45
		x"b6",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"d5",	--50
		x"b0",	--51
		x"08",	--52
		x"21",	--53
		x"3e",	--54
		x"8e",	--55
		x"7f",	--56
		x"77",	--57
		x"b0",	--58
		x"b8",	--59
		x"3e",	--60
		x"2e",	--61
		x"7f",	--62
		x"72",	--63
		x"b0",	--64
		x"b8",	--65
		x"3e",	--66
		x"dc",	--67
		x"7f",	--68
		x"70",	--69
		x"b0",	--70
		x"b8",	--71
		x"3e",	--72
		x"a6",	--73
		x"7f",	--74
		x"62",	--75
		x"b0",	--76
		x"b8",	--77
		x"2c",	--78
		x"3d",	--79
		x"20",	--80
		x"3e",	--81
		x"80",	--82
		x"0f",	--83
		x"3f",	--84
		x"0a",	--85
		x"b0",	--86
		x"c6",	--87
		x"0f",	--88
		x"3f",	--89
		x"0a",	--90
		x"b0",	--91
		x"0e",	--92
		x"2c",	--93
		x"3d",	--94
		x"20",	--95
		x"3e",	--96
		x"88",	--97
		x"0f",	--98
		x"b0",	--99
		x"c6",	--100
		x"0f",	--101
		x"b0",	--102
		x"0e",	--103
		x"0e",	--104
		x"0f",	--105
		x"3f",	--106
		x"0a",	--107
		x"b0",	--108
		x"d2",	--109
		x"f2",	--110
		x"80",	--111
		x"19",	--112
		x"32",	--113
		x"0b",	--114
		x"30",	--115
		x"f2",	--116
		x"b0",	--117
		x"08",	--118
		x"21",	--119
		x"0a",	--120
		x"32",	--121
		x"10",	--122
		x"1b",	--123
		x"3b",	--124
		x"09",	--125
		x"0a",	--126
		x"1f",	--127
		x"4e",	--128
		x"7e",	--129
		x"0f",	--130
		x"03",	--131
		x"0f",	--132
		x"7e",	--133
		x"fd",	--134
		x"4f",	--135
		x"02",	--136
		x"5f",	--137
		x"0b",	--138
		x"c2",	--139
		x"19",	--140
		x"b0",	--141
		x"58",	--142
		x"0f",	--143
		x"e8",	--144
		x"b0",	--145
		x"80",	--146
		x"7f",	--147
		x"1c",	--148
		x"7f",	--149
		x"0d",	--150
		x"22",	--151
		x"30",	--152
		x"f5",	--153
		x"b0",	--154
		x"08",	--155
		x"21",	--156
		x"3f",	--157
		x"14",	--158
		x"0f",	--159
		x"0a",	--160
		x"ca",	--161
		x"00",	--162
		x"0f",	--163
		x"30",	--164
		x"f8",	--165
		x"b0",	--166
		x"08",	--167
		x"21",	--168
		x"0e",	--169
		x"3e",	--170
		x"14",	--171
		x"5f",	--172
		x"14",	--173
		x"b0",	--174
		x"e2",	--175
		x"c2",	--176
		x"0a",	--177
		x"c6",	--178
		x"3a",	--179
		x"30",	--180
		x"fe",	--181
		x"b0",	--182
		x"08",	--183
		x"21",	--184
		x"bf",	--185
		x"3a",	--186
		x"28",	--187
		x"bc",	--188
		x"4e",	--189
		x"8e",	--190
		x"0e",	--191
		x"30",	--192
		x"02",	--193
		x"81",	--194
		x"40",	--195
		x"b0",	--196
		x"08",	--197
		x"21",	--198
		x"3e",	--199
		x"14",	--200
		x"0e",	--201
		x"0e",	--202
		x"1f",	--203
		x"3c",	--204
		x"ce",	--205
		x"00",	--206
		x"1a",	--207
		x"a8",	--208
		x"30",	--209
		x"54",	--210
		x"b2",	--211
		x"00",	--212
		x"92",	--213
		x"a2",	--214
		x"94",	--215
		x"b2",	--216
		x"6d",	--217
		x"96",	--218
		x"30",	--219
		x"5c",	--220
		x"b0",	--221
		x"08",	--222
		x"92",	--223
		x"90",	--224
		x"b1",	--225
		x"7a",	--226
		x"00",	--227
		x"b0",	--228
		x"08",	--229
		x"21",	--230
		x"0f",	--231
		x"30",	--232
		x"82",	--233
		x"08",	--234
		x"82",	--235
		x"06",	--236
		x"30",	--237
		x"31",	--238
		x"ff",	--239
		x"20",	--240
		x"01",	--241
		x"39",	--242
		x"cf",	--243
		x"02",	--244
		x"36",	--245
		x"0d",	--246
		x"0e",	--247
		x"2e",	--248
		x"0f",	--249
		x"2f",	--250
		x"b0",	--251
		x"ac",	--252
		x"81",	--253
		x"00",	--254
		x"40",	--255
		x"0d",	--256
		x"0e",	--257
		x"0f",	--258
		x"2f",	--259
		x"b0",	--260
		x"ac",	--261
		x"81",	--262
		x"00",	--263
		x"37",	--264
		x"1e",	--265
		x"04",	--266
		x"0f",	--267
		x"b0",	--268
		x"72",	--269
		x"0c",	--270
		x"3d",	--271
		x"c8",	--272
		x"b0",	--273
		x"42",	--274
		x"0d",	--275
		x"0e",	--276
		x"1f",	--277
		x"08",	--278
		x"b0",	--279
		x"62",	--280
		x"1e",	--281
		x"02",	--282
		x"0f",	--283
		x"b0",	--284
		x"72",	--285
		x"0c",	--286
		x"3d",	--287
		x"c8",	--288
		x"b0",	--289
		x"42",	--290
		x"0d",	--291
		x"0e",	--292
		x"1f",	--293
		x"06",	--294
		x"b0",	--295
		x"62",	--296
		x"0f",	--297
		x"31",	--298
		x"30",	--299
		x"30",	--300
		x"93",	--301
		x"81",	--302
		x"08",	--303
		x"b0",	--304
		x"08",	--305
		x"1f",	--306
		x"08",	--307
		x"6f",	--308
		x"8f",	--309
		x"81",	--310
		x"00",	--311
		x"30",	--312
		x"a4",	--313
		x"b0",	--314
		x"08",	--315
		x"21",	--316
		x"3f",	--317
		x"31",	--318
		x"30",	--319
		x"30",	--320
		x"b5",	--321
		x"b0",	--322
		x"08",	--323
		x"21",	--324
		x"3f",	--325
		x"e3",	--326
		x"0b",	--327
		x"31",	--328
		x"fa",	--329
		x"0b",	--330
		x"30",	--331
		x"05",	--332
		x"b0",	--333
		x"08",	--334
		x"21",	--335
		x"fb",	--336
		x"20",	--337
		x"01",	--338
		x"2a",	--339
		x"cb",	--340
		x"02",	--341
		x"27",	--342
		x"0d",	--343
		x"0e",	--344
		x"2e",	--345
		x"0f",	--346
		x"2f",	--347
		x"b0",	--348
		x"ac",	--349
		x"81",	--350
		x"00",	--351
		x"2f",	--352
		x"0d",	--353
		x"0e",	--354
		x"0f",	--355
		x"2f",	--356
		x"b0",	--357
		x"ac",	--358
		x"81",	--359
		x"00",	--360
		x"26",	--361
		x"11",	--362
		x"04",	--363
		x"11",	--364
		x"08",	--365
		x"30",	--366
		x"53",	--367
		x"b0",	--368
		x"08",	--369
		x"31",	--370
		x"06",	--371
		x"1f",	--372
		x"04",	--373
		x"9f",	--374
		x"02",	--375
		x"00",	--376
		x"0f",	--377
		x"31",	--378
		x"06",	--379
		x"3b",	--380
		x"30",	--381
		x"30",	--382
		x"0d",	--383
		x"b0",	--384
		x"08",	--385
		x"6f",	--386
		x"8f",	--387
		x"81",	--388
		x"00",	--389
		x"30",	--390
		x"1e",	--391
		x"b0",	--392
		x"08",	--393
		x"21",	--394
		x"3f",	--395
		x"31",	--396
		x"06",	--397
		x"3b",	--398
		x"30",	--399
		x"30",	--400
		x"33",	--401
		x"b0",	--402
		x"08",	--403
		x"21",	--404
		x"3f",	--405
		x"e3",	--406
		x"0b",	--407
		x"21",	--408
		x"0b",	--409
		x"30",	--410
		x"5f",	--411
		x"b0",	--412
		x"08",	--413
		x"21",	--414
		x"fb",	--415
		x"20",	--416
		x"01",	--417
		x"1b",	--418
		x"cb",	--419
		x"02",	--420
		x"18",	--421
		x"0d",	--422
		x"0e",	--423
		x"2e",	--424
		x"0f",	--425
		x"2f",	--426
		x"b0",	--427
		x"ac",	--428
		x"81",	--429
		x"00",	--430
		x"1f",	--431
		x"1f",	--432
		x"02",	--433
		x"2f",	--434
		x"0f",	--435
		x"30",	--436
		x"53",	--437
		x"b0",	--438
		x"08",	--439
		x"31",	--440
		x"06",	--441
		x"0f",	--442
		x"21",	--443
		x"3b",	--444
		x"30",	--445
		x"30",	--446
		x"0d",	--447
		x"b0",	--448
		x"08",	--449
		x"6f",	--450
		x"8f",	--451
		x"81",	--452
		x"00",	--453
		x"30",	--454
		x"66",	--455
		x"b0",	--456
		x"08",	--457
		x"21",	--458
		x"3f",	--459
		x"21",	--460
		x"3b",	--461
		x"30",	--462
		x"30",	--463
		x"33",	--464
		x"b0",	--465
		x"08",	--466
		x"21",	--467
		x"3f",	--468
		x"e5",	--469
		x"0b",	--470
		x"0a",	--471
		x"09",	--472
		x"08",	--473
		x"07",	--474
		x"8f",	--475
		x"00",	--476
		x"8d",	--477
		x"00",	--478
		x"6c",	--479
		x"4c",	--480
		x"5f",	--481
		x"0b",	--482
		x"1b",	--483
		x"08",	--484
		x"0a",	--485
		x"07",	--486
		x"09",	--487
		x"18",	--488
		x"7a",	--489
		x"0a",	--490
		x"35",	--491
		x"2c",	--492
		x"0c",	--493
		x"0c",	--494
		x"0c",	--495
		x"0c",	--496
		x"8f",	--497
		x"00",	--498
		x"3c",	--499
		x"d0",	--500
		x"6a",	--501
		x"8a",	--502
		x"0c",	--503
		x"8f",	--504
		x"00",	--505
		x"17",	--506
		x"19",	--507
		x"0a",	--508
		x"08",	--509
		x"7c",	--510
		x"4c",	--511
		x"40",	--512
		x"7c",	--513
		x"78",	--514
		x"1b",	--515
		x"7c",	--516
		x"20",	--517
		x"43",	--518
		x"4a",	--519
		x"7a",	--520
		x"d0",	--521
		x"07",	--522
		x"dd",	--523
		x"7a",	--524
		x"0a",	--525
		x"46",	--526
		x"2a",	--527
		x"0a",	--528
		x"0c",	--529
		x"0c",	--530
		x"0c",	--531
		x"0c",	--532
		x"8f",	--533
		x"00",	--534
		x"3c",	--535
		x"d0",	--536
		x"68",	--537
		x"88",	--538
		x"0c",	--539
		x"8f",	--540
		x"00",	--541
		x"dc",	--542
		x"17",	--543
		x"da",	--544
		x"4a",	--545
		x"7a",	--546
		x"9f",	--547
		x"7a",	--548
		x"06",	--549
		x"0a",	--550
		x"2c",	--551
		x"0c",	--552
		x"0c",	--553
		x"0c",	--554
		x"0c",	--555
		x"8f",	--556
		x"00",	--557
		x"3c",	--558
		x"a9",	--559
		x"c4",	--560
		x"4a",	--561
		x"7a",	--562
		x"bf",	--563
		x"7a",	--564
		x"06",	--565
		x"1e",	--566
		x"2c",	--567
		x"0c",	--568
		x"0c",	--569
		x"0c",	--570
		x"0c",	--571
		x"8f",	--572
		x"00",	--573
		x"3c",	--574
		x"c9",	--575
		x"b4",	--576
		x"9d",	--577
		x"00",	--578
		x"0f",	--579
		x"37",	--580
		x"38",	--581
		x"39",	--582
		x"3a",	--583
		x"3b",	--584
		x"30",	--585
		x"9d",	--586
		x"00",	--587
		x"0f",	--588
		x"1f",	--589
		x"0f",	--590
		x"37",	--591
		x"38",	--592
		x"39",	--593
		x"3a",	--594
		x"3b",	--595
		x"30",	--596
		x"8c",	--597
		x"0c",	--598
		x"30",	--599
		x"75",	--600
		x"b0",	--601
		x"08",	--602
		x"21",	--603
		x"0f",	--604
		x"37",	--605
		x"38",	--606
		x"39",	--607
		x"3a",	--608
		x"3b",	--609
		x"30",	--610
		x"0b",	--611
		x"0a",	--612
		x"0b",	--613
		x"0a",	--614
		x"8f",	--615
		x"00",	--616
		x"8f",	--617
		x"02",	--618
		x"8f",	--619
		x"04",	--620
		x"0c",	--621
		x"0d",	--622
		x"3e",	--623
		x"00",	--624
		x"3f",	--625
		x"6e",	--626
		x"b0",	--627
		x"a6",	--628
		x"8b",	--629
		x"02",	--630
		x"02",	--631
		x"32",	--632
		x"03",	--633
		x"82",	--634
		x"32",	--635
		x"b2",	--636
		x"18",	--637
		x"38",	--638
		x"9b",	--639
		x"3a",	--640
		x"06",	--641
		x"32",	--642
		x"0f",	--643
		x"3a",	--644
		x"3b",	--645
		x"30",	--646
		x"0b",	--647
		x"09",	--648
		x"08",	--649
		x"8f",	--650
		x"06",	--651
		x"bf",	--652
		x"00",	--653
		x"08",	--654
		x"2b",	--655
		x"1e",	--656
		x"02",	--657
		x"0f",	--658
		x"b0",	--659
		x"72",	--660
		x"0c",	--661
		x"3d",	--662
		x"00",	--663
		x"b0",	--664
		x"1e",	--665
		x"08",	--666
		x"09",	--667
		x"1e",	--668
		x"06",	--669
		x"0f",	--670
		x"b0",	--671
		x"72",	--672
		x"0c",	--673
		x"0d",	--674
		x"0e",	--675
		x"0f",	--676
		x"b0",	--677
		x"ce",	--678
		x"b0",	--679
		x"ae",	--680
		x"8b",	--681
		x"04",	--682
		x"9b",	--683
		x"00",	--684
		x"38",	--685
		x"39",	--686
		x"3b",	--687
		x"30",	--688
		x"0b",	--689
		x"0a",	--690
		x"09",	--691
		x"0a",	--692
		x"0b",	--693
		x"8f",	--694
		x"06",	--695
		x"8f",	--696
		x"08",	--697
		x"29",	--698
		x"1e",	--699
		x"02",	--700
		x"0f",	--701
		x"b0",	--702
		x"72",	--703
		x"0c",	--704
		x"0d",	--705
		x"0e",	--706
		x"0f",	--707
		x"b0",	--708
		x"1e",	--709
		x"0a",	--710
		x"0b",	--711
		x"1e",	--712
		x"06",	--713
		x"0f",	--714
		x"b0",	--715
		x"72",	--716
		x"0c",	--717
		x"0d",	--718
		x"0e",	--719
		x"0f",	--720
		x"b0",	--721
		x"ce",	--722
		x"b0",	--723
		x"ae",	--724
		x"89",	--725
		x"04",	--726
		x"39",	--727
		x"3a",	--728
		x"3b",	--729
		x"30",	--730
		x"30",	--731
		x"1c",	--732
		x"00",	--733
		x"3c",	--734
		x"40",	--735
		x"0e",	--736
		x"0d",	--737
		x"0d",	--738
		x"0d",	--739
		x"3d",	--740
		x"0a",	--741
		x"cd",	--742
		x"00",	--743
		x"8d",	--744
		x"02",	--745
		x"1c",	--746
		x"82",	--747
		x"00",	--748
		x"0f",	--749
		x"30",	--750
		x"3f",	--751
		x"30",	--752
		x"0b",	--753
		x"1b",	--754
		x"00",	--755
		x"1b",	--756
		x"0e",	--757
		x"5f",	--758
		x"0a",	--759
		x"13",	--760
		x"3d",	--761
		x"0e",	--762
		x"0c",	--763
		x"04",	--764
		x"2d",	--765
		x"cd",	--766
		x"fc",	--767
		x"0c",	--768
		x"1c",	--769
		x"0c",	--770
		x"f9",	--771
		x"30",	--772
		x"8a",	--773
		x"b0",	--774
		x"08",	--775
		x"21",	--776
		x"3f",	--777
		x"3b",	--778
		x"30",	--779
		x"0c",	--780
		x"0c",	--781
		x"0c",	--782
		x"3c",	--783
		x"0a",	--784
		x"0f",	--785
		x"9c",	--786
		x"02",	--787
		x"3b",	--788
		x"30",	--789
		x"5e",	--790
		x"81",	--791
		x"3e",	--792
		x"fc",	--793
		x"c2",	--794
		x"84",	--795
		x"0f",	--796
		x"30",	--797
		x"3f",	--798
		x"0f",	--799
		x"5f",	--800
		x"48",	--801
		x"8f",	--802
		x"b0",	--803
		x"2c",	--804
		x"30",	--805
		x"0b",	--806
		x"0b",	--807
		x"0e",	--808
		x"0e",	--809
		x"0e",	--810
		x"0e",	--811
		x"0e",	--812
		x"0f",	--813
		x"b0",	--814
		x"3c",	--815
		x"0f",	--816
		x"b0",	--817
		x"3c",	--818
		x"3b",	--819
		x"30",	--820
		x"0b",	--821
		x"0a",	--822
		x"0a",	--823
		x"3b",	--824
		x"07",	--825
		x"0e",	--826
		x"4d",	--827
		x"7d",	--828
		x"0f",	--829
		x"03",	--830
		x"0e",	--831
		x"7d",	--832
		x"fd",	--833
		x"1e",	--834
		x"0a",	--835
		x"3f",	--836
		x"31",	--837
		x"b0",	--838
		x"2c",	--839
		x"3b",	--840
		x"3b",	--841
		x"ef",	--842
		x"3a",	--843
		x"3b",	--844
		x"30",	--845
		x"3f",	--846
		x"30",	--847
		x"f5",	--848
		x"0b",	--849
		x"0b",	--850
		x"0e",	--851
		x"8e",	--852
		x"8e",	--853
		x"0f",	--854
		x"b0",	--855
		x"4c",	--856
		x"0f",	--857
		x"b0",	--858
		x"4c",	--859
		x"3b",	--860
		x"30",	--861
		x"0b",	--862
		x"0a",	--863
		x"0a",	--864
		x"0b",	--865
		x"0d",	--866
		x"8d",	--867
		x"8d",	--868
		x"0f",	--869
		x"b0",	--870
		x"4c",	--871
		x"0f",	--872
		x"b0",	--873
		x"4c",	--874
		x"0c",	--875
		x"0d",	--876
		x"8d",	--877
		x"8c",	--878
		x"4d",	--879
		x"0d",	--880
		x"0f",	--881
		x"b0",	--882
		x"4c",	--883
		x"0f",	--884
		x"b0",	--885
		x"4c",	--886
		x"3a",	--887
		x"3b",	--888
		x"30",	--889
		x"0b",	--890
		x"0a",	--891
		x"09",	--892
		x"0a",	--893
		x"0e",	--894
		x"19",	--895
		x"09",	--896
		x"39",	--897
		x"0b",	--898
		x"0d",	--899
		x"0d",	--900
		x"6f",	--901
		x"8f",	--902
		x"b0",	--903
		x"4c",	--904
		x"0b",	--905
		x"0e",	--906
		x"1b",	--907
		x"3b",	--908
		x"07",	--909
		x"05",	--910
		x"3f",	--911
		x"20",	--912
		x"b0",	--913
		x"2c",	--914
		x"ef",	--915
		x"3f",	--916
		x"3a",	--917
		x"b0",	--918
		x"2c",	--919
		x"ea",	--920
		x"39",	--921
		x"3a",	--922
		x"3b",	--923
		x"30",	--924
		x"0b",	--925
		x"0a",	--926
		x"09",	--927
		x"0a",	--928
		x"0e",	--929
		x"17",	--930
		x"09",	--931
		x"39",	--932
		x"0b",	--933
		x"6f",	--934
		x"8f",	--935
		x"b0",	--936
		x"3c",	--937
		x"0b",	--938
		x"0e",	--939
		x"1b",	--940
		x"3b",	--941
		x"07",	--942
		x"f6",	--943
		x"3f",	--944
		x"20",	--945
		x"b0",	--946
		x"2c",	--947
		x"6f",	--948
		x"8f",	--949
		x"b0",	--950
		x"3c",	--951
		x"0b",	--952
		x"f2",	--953
		x"39",	--954
		x"3a",	--955
		x"3b",	--956
		x"30",	--957
		x"0b",	--958
		x"0a",	--959
		x"09",	--960
		x"31",	--961
		x"ec",	--962
		x"0b",	--963
		x"0f",	--964
		x"34",	--965
		x"3b",	--966
		x"0a",	--967
		x"38",	--968
		x"09",	--969
		x"0a",	--970
		x"0a",	--971
		x"3e",	--972
		x"0a",	--973
		x"0f",	--974
		x"b0",	--975
		x"9e",	--976
		x"7f",	--977
		x"30",	--978
		x"ca",	--979
		x"00",	--980
		x"19",	--981
		x"3e",	--982
		x"0a",	--983
		x"0f",	--984
		x"b0",	--985
		x"6c",	--986
		x"0b",	--987
		x"3f",	--988
		x"0a",	--989
		x"eb",	--990
		x"0a",	--991
		x"1a",	--992
		x"09",	--993
		x"3e",	--994
		x"0a",	--995
		x"0f",	--996
		x"b0",	--997
		x"9e",	--998
		x"7f",	--999
		x"30",	--1000
		x"c9",	--1001
		x"00",	--1002
		x"3a",	--1003
		x"0f",	--1004
		x"0f",	--1005
		x"6f",	--1006
		x"8f",	--1007
		x"b0",	--1008
		x"2c",	--1009
		x"0a",	--1010
		x"f7",	--1011
		x"31",	--1012
		x"14",	--1013
		x"39",	--1014
		x"3a",	--1015
		x"3b",	--1016
		x"30",	--1017
		x"3f",	--1018
		x"2d",	--1019
		x"b0",	--1020
		x"2c",	--1021
		x"3b",	--1022
		x"1b",	--1023
		x"c5",	--1024
		x"1a",	--1025
		x"09",	--1026
		x"dd",	--1027
		x"0b",	--1028
		x"0a",	--1029
		x"09",	--1030
		x"0b",	--1031
		x"3b",	--1032
		x"39",	--1033
		x"6f",	--1034
		x"4f",	--1035
		x"0b",	--1036
		x"1a",	--1037
		x"8f",	--1038
		x"b0",	--1039
		x"2c",	--1040
		x"0a",	--1041
		x"09",	--1042
		x"19",	--1043
		x"5f",	--1044
		x"01",	--1045
		x"4f",	--1046
		x"10",	--1047
		x"7f",	--1048
		x"25",	--1049
		x"f3",	--1050
		x"0a",	--1051
		x"1a",	--1052
		x"5f",	--1053
		x"01",	--1054
		x"7f",	--1055
		x"db",	--1056
		x"7f",	--1057
		x"54",	--1058
		x"ee",	--1059
		x"4f",	--1060
		x"0f",	--1061
		x"10",	--1062
		x"a0",	--1063
		x"39",	--1064
		x"3a",	--1065
		x"3b",	--1066
		x"30",	--1067
		x"09",	--1068
		x"29",	--1069
		x"1e",	--1070
		x"02",	--1071
		x"2f",	--1072
		x"b0",	--1073
		x"f4",	--1074
		x"0b",	--1075
		x"dd",	--1076
		x"09",	--1077
		x"29",	--1078
		x"2f",	--1079
		x"b0",	--1080
		x"a2",	--1081
		x"0b",	--1082
		x"d6",	--1083
		x"0f",	--1084
		x"2b",	--1085
		x"29",	--1086
		x"6f",	--1087
		x"4f",	--1088
		x"d0",	--1089
		x"19",	--1090
		x"8f",	--1091
		x"b0",	--1092
		x"2c",	--1093
		x"7f",	--1094
		x"4f",	--1095
		x"fa",	--1096
		x"c8",	--1097
		x"09",	--1098
		x"29",	--1099
		x"1e",	--1100
		x"02",	--1101
		x"2f",	--1102
		x"b0",	--1103
		x"3a",	--1104
		x"0b",	--1105
		x"bf",	--1106
		x"09",	--1107
		x"29",	--1108
		x"2e",	--1109
		x"0f",	--1110
		x"8f",	--1111
		x"8f",	--1112
		x"8f",	--1113
		x"8f",	--1114
		x"b0",	--1115
		x"bc",	--1116
		x"0b",	--1117
		x"b3",	--1118
		x"09",	--1119
		x"29",	--1120
		x"2f",	--1121
		x"b0",	--1122
		x"7c",	--1123
		x"0b",	--1124
		x"ac",	--1125
		x"09",	--1126
		x"29",	--1127
		x"2f",	--1128
		x"b0",	--1129
		x"2c",	--1130
		x"0b",	--1131
		x"a5",	--1132
		x"09",	--1133
		x"29",	--1134
		x"2f",	--1135
		x"b0",	--1136
		x"4c",	--1137
		x"0b",	--1138
		x"9e",	--1139
		x"09",	--1140
		x"29",	--1141
		x"2f",	--1142
		x"b0",	--1143
		x"6a",	--1144
		x"0b",	--1145
		x"97",	--1146
		x"3f",	--1147
		x"25",	--1148
		x"b0",	--1149
		x"2c",	--1150
		x"92",	--1151
		x"0f",	--1152
		x"0e",	--1153
		x"1f",	--1154
		x"02",	--1155
		x"df",	--1156
		x"85",	--1157
		x"0a",	--1158
		x"1f",	--1159
		x"02",	--1160
		x"3f",	--1161
		x"3f",	--1162
		x"16",	--1163
		x"92",	--1164
		x"02",	--1165
		x"1e",	--1166
		x"02",	--1167
		x"1f",	--1168
		x"04",	--1169
		x"0e",	--1170
		x"02",	--1171
		x"92",	--1172
		x"04",	--1173
		x"f2",	--1174
		x"10",	--1175
		x"81",	--1176
		x"b1",	--1177
		x"10",	--1178
		x"04",	--1179
		x"3e",	--1180
		x"3f",	--1181
		x"b1",	--1182
		x"f0",	--1183
		x"00",	--1184
		x"00",	--1185
		x"82",	--1186
		x"02",	--1187
		x"e9",	--1188
		x"b2",	--1189
		x"c3",	--1190
		x"82",	--1191
		x"f2",	--1192
		x"11",	--1193
		x"80",	--1194
		x"30",	--1195
		x"1e",	--1196
		x"02",	--1197
		x"1f",	--1198
		x"04",	--1199
		x"0e",	--1200
		x"05",	--1201
		x"1f",	--1202
		x"02",	--1203
		x"1f",	--1204
		x"04",	--1205
		x"30",	--1206
		x"1d",	--1207
		x"02",	--1208
		x"1e",	--1209
		x"04",	--1210
		x"3f",	--1211
		x"40",	--1212
		x"0f",	--1213
		x"0f",	--1214
		x"30",	--1215
		x"1f",	--1216
		x"04",	--1217
		x"5f",	--1218
		x"0a",	--1219
		x"1d",	--1220
		x"04",	--1221
		x"1e",	--1222
		x"02",	--1223
		x"0d",	--1224
		x"0b",	--1225
		x"1e",	--1226
		x"04",	--1227
		x"3e",	--1228
		x"3f",	--1229
		x"03",	--1230
		x"82",	--1231
		x"04",	--1232
		x"30",	--1233
		x"92",	--1234
		x"04",	--1235
		x"30",	--1236
		x"4f",	--1237
		x"30",	--1238
		x"0b",	--1239
		x"0a",	--1240
		x"0a",	--1241
		x"0b",	--1242
		x"0c",	--1243
		x"3d",	--1244
		x"00",	--1245
		x"b0",	--1246
		x"92",	--1247
		x"0f",	--1248
		x"07",	--1249
		x"0e",	--1250
		x"0f",	--1251
		x"b0",	--1252
		x"e2",	--1253
		x"3a",	--1254
		x"3b",	--1255
		x"30",	--1256
		x"0c",	--1257
		x"3d",	--1258
		x"00",	--1259
		x"0e",	--1260
		x"0f",	--1261
		x"b0",	--1262
		x"ce",	--1263
		x"b0",	--1264
		x"e2",	--1265
		x"0e",	--1266
		x"3f",	--1267
		x"00",	--1268
		x"3a",	--1269
		x"3b",	--1270
		x"30",	--1271
		x"0b",	--1272
		x"0a",	--1273
		x"09",	--1274
		x"08",	--1275
		x"07",	--1276
		x"06",	--1277
		x"05",	--1278
		x"04",	--1279
		x"31",	--1280
		x"fa",	--1281
		x"08",	--1282
		x"6b",	--1283
		x"6b",	--1284
		x"67",	--1285
		x"6c",	--1286
		x"6c",	--1287
		x"e9",	--1288
		x"6b",	--1289
		x"02",	--1290
		x"30",	--1291
		x"70",	--1292
		x"6c",	--1293
		x"e3",	--1294
		x"6c",	--1295
		x"bb",	--1296
		x"6b",	--1297
		x"df",	--1298
		x"91",	--1299
		x"02",	--1300
		x"00",	--1301
		x"1b",	--1302
		x"02",	--1303
		x"14",	--1304
		x"04",	--1305
		x"15",	--1306
		x"06",	--1307
		x"16",	--1308
		x"04",	--1309
		x"17",	--1310
		x"06",	--1311
		x"2c",	--1312
		x"0c",	--1313
		x"09",	--1314
		x"0c",	--1315
		x"bf",	--1316
		x"39",	--1317
		x"20",	--1318
		x"50",	--1319
		x"1c",	--1320
		x"d7",	--1321
		x"81",	--1322
		x"02",	--1323
		x"81",	--1324
		x"04",	--1325
		x"4c",	--1326
		x"7c",	--1327
		x"1f",	--1328
		x"0b",	--1329
		x"0a",	--1330
		x"0b",	--1331
		x"12",	--1332
		x"0b",	--1333
		x"0a",	--1334
		x"7c",	--1335
		x"fb",	--1336
		x"81",	--1337
		x"02",	--1338
		x"81",	--1339
		x"04",	--1340
		x"1c",	--1341
		x"0d",	--1342
		x"79",	--1343
		x"1f",	--1344
		x"04",	--1345
		x"0c",	--1346
		x"0d",	--1347
		x"79",	--1348
		x"fc",	--1349
		x"3c",	--1350
		x"3d",	--1351
		x"0c",	--1352
		x"0d",	--1353
		x"1a",	--1354
		x"0b",	--1355
		x"0c",	--1356
		x"02",	--1357
		x"0d",	--1358
		x"e5",	--1359
		x"16",	--1360
		x"02",	--1361
		x"17",	--1362
		x"04",	--1363
		x"06",	--1364
		x"07",	--1365
		x"5f",	--1366
		x"01",	--1367
		x"5f",	--1368
		x"01",	--1369
		x"28",	--1370
		x"c8",	--1371
		x"01",	--1372
		x"a8",	--1373
		x"02",	--1374
		x"0e",	--1375
		x"0f",	--1376
		x"0e",	--1377
		x"0f",	--1378
		x"88",	--1379
		x"04",	--1380
		x"88",	--1381
		x"06",	--1382
		x"f8",	--1383
		x"03",	--1384
		x"00",	--1385
		x"0f",	--1386
		x"4d",	--1387
		x"0f",	--1388
		x"31",	--1389
		x"06",	--1390
		x"34",	--1391
		x"35",	--1392
		x"36",	--1393
		x"37",	--1394
		x"38",	--1395
		x"39",	--1396
		x"3a",	--1397
		x"3b",	--1398
		x"30",	--1399
		x"2b",	--1400
		x"67",	--1401
		x"81",	--1402
		x"00",	--1403
		x"04",	--1404
		x"05",	--1405
		x"5f",	--1406
		x"01",	--1407
		x"5f",	--1408
		x"01",	--1409
		x"d8",	--1410
		x"4f",	--1411
		x"68",	--1412
		x"0e",	--1413
		x"0f",	--1414
		x"0e",	--1415
		x"0f",	--1416
		x"0f",	--1417
		x"69",	--1418
		x"c8",	--1419
		x"01",	--1420
		x"a8",	--1421
		x"02",	--1422
		x"88",	--1423
		x"04",	--1424
		x"88",	--1425
		x"06",	--1426
		x"0c",	--1427
		x"0d",	--1428
		x"3c",	--1429
		x"3d",	--1430
		x"3d",	--1431
		x"ff",	--1432
		x"05",	--1433
		x"3d",	--1434
		x"00",	--1435
		x"17",	--1436
		x"3c",	--1437
		x"15",	--1438
		x"1b",	--1439
		x"02",	--1440
		x"3b",	--1441
		x"0e",	--1442
		x"0f",	--1443
		x"0a",	--1444
		x"3b",	--1445
		x"0c",	--1446
		x"0d",	--1447
		x"3c",	--1448
		x"3d",	--1449
		x"3d",	--1450
		x"ff",	--1451
		x"f5",	--1452
		x"3c",	--1453
		x"88",	--1454
		x"04",	--1455
		x"88",	--1456
		x"06",	--1457
		x"88",	--1458
		x"02",	--1459
		x"f8",	--1460
		x"03",	--1461
		x"00",	--1462
		x"0f",	--1463
		x"b3",	--1464
		x"0c",	--1465
		x"0d",	--1466
		x"1c",	--1467
		x"0d",	--1468
		x"12",	--1469
		x"0f",	--1470
		x"0e",	--1471
		x"0a",	--1472
		x"0b",	--1473
		x"0a",	--1474
		x"0b",	--1475
		x"88",	--1476
		x"04",	--1477
		x"88",	--1478
		x"06",	--1479
		x"98",	--1480
		x"02",	--1481
		x"0f",	--1482
		x"a1",	--1483
		x"6b",	--1484
		x"9f",	--1485
		x"ad",	--1486
		x"00",	--1487
		x"9d",	--1488
		x"02",	--1489
		x"02",	--1490
		x"9d",	--1491
		x"04",	--1492
		x"04",	--1493
		x"9d",	--1494
		x"06",	--1495
		x"06",	--1496
		x"5e",	--1497
		x"01",	--1498
		x"5e",	--1499
		x"01",	--1500
		x"cd",	--1501
		x"01",	--1502
		x"0f",	--1503
		x"8c",	--1504
		x"06",	--1505
		x"07",	--1506
		x"9a",	--1507
		x"39",	--1508
		x"19",	--1509
		x"39",	--1510
		x"20",	--1511
		x"8f",	--1512
		x"3e",	--1513
		x"3c",	--1514
		x"b6",	--1515
		x"c1",	--1516
		x"0e",	--1517
		x"0f",	--1518
		x"0e",	--1519
		x"0f",	--1520
		x"97",	--1521
		x"0f",	--1522
		x"79",	--1523
		x"d8",	--1524
		x"01",	--1525
		x"a8",	--1526
		x"02",	--1527
		x"3e",	--1528
		x"3f",	--1529
		x"1e",	--1530
		x"0f",	--1531
		x"88",	--1532
		x"04",	--1533
		x"88",	--1534
		x"06",	--1535
		x"92",	--1536
		x"0c",	--1537
		x"7b",	--1538
		x"81",	--1539
		x"00",	--1540
		x"81",	--1541
		x"02",	--1542
		x"81",	--1543
		x"04",	--1544
		x"4d",	--1545
		x"7d",	--1546
		x"1f",	--1547
		x"0c",	--1548
		x"4b",	--1549
		x"0c",	--1550
		x"0d",	--1551
		x"12",	--1552
		x"0d",	--1553
		x"0c",	--1554
		x"7b",	--1555
		x"fb",	--1556
		x"81",	--1557
		x"02",	--1558
		x"81",	--1559
		x"04",	--1560
		x"1c",	--1561
		x"0d",	--1562
		x"79",	--1563
		x"1f",	--1564
		x"04",	--1565
		x"0c",	--1566
		x"0d",	--1567
		x"79",	--1568
		x"fc",	--1569
		x"3c",	--1570
		x"3d",	--1571
		x"0c",	--1572
		x"0d",	--1573
		x"1a",	--1574
		x"0b",	--1575
		x"0c",	--1576
		x"04",	--1577
		x"0d",	--1578
		x"02",	--1579
		x"0a",	--1580
		x"0b",	--1581
		x"14",	--1582
		x"02",	--1583
		x"15",	--1584
		x"04",	--1585
		x"04",	--1586
		x"05",	--1587
		x"49",	--1588
		x"0a",	--1589
		x"0b",	--1590
		x"18",	--1591
		x"6c",	--1592
		x"33",	--1593
		x"df",	--1594
		x"01",	--1595
		x"01",	--1596
		x"2f",	--1597
		x"3f",	--1598
		x"5a",	--1599
		x"2c",	--1600
		x"31",	--1601
		x"e0",	--1602
		x"81",	--1603
		x"04",	--1604
		x"81",	--1605
		x"06",	--1606
		x"81",	--1607
		x"00",	--1608
		x"81",	--1609
		x"02",	--1610
		x"0e",	--1611
		x"3e",	--1612
		x"18",	--1613
		x"0f",	--1614
		x"2f",	--1615
		x"b0",	--1616
		x"a4",	--1617
		x"0e",	--1618
		x"3e",	--1619
		x"10",	--1620
		x"0f",	--1621
		x"b0",	--1622
		x"a4",	--1623
		x"0d",	--1624
		x"3d",	--1625
		x"0e",	--1626
		x"3e",	--1627
		x"10",	--1628
		x"0f",	--1629
		x"3f",	--1630
		x"18",	--1631
		x"b0",	--1632
		x"f0",	--1633
		x"b0",	--1634
		x"c6",	--1635
		x"31",	--1636
		x"20",	--1637
		x"30",	--1638
		x"31",	--1639
		x"e0",	--1640
		x"81",	--1641
		x"04",	--1642
		x"81",	--1643
		x"06",	--1644
		x"81",	--1645
		x"00",	--1646
		x"81",	--1647
		x"02",	--1648
		x"0e",	--1649
		x"3e",	--1650
		x"18",	--1651
		x"0f",	--1652
		x"2f",	--1653
		x"b0",	--1654
		x"a4",	--1655
		x"0e",	--1656
		x"3e",	--1657
		x"10",	--1658
		x"0f",	--1659
		x"b0",	--1660
		x"a4",	--1661
		x"d1",	--1662
		x"11",	--1663
		x"0d",	--1664
		x"3d",	--1665
		x"0e",	--1666
		x"3e",	--1667
		x"10",	--1668
		x"0f",	--1669
		x"3f",	--1670
		x"18",	--1671
		x"b0",	--1672
		x"f0",	--1673
		x"b0",	--1674
		x"c6",	--1675
		x"31",	--1676
		x"20",	--1677
		x"30",	--1678
		x"0b",	--1679
		x"0a",	--1680
		x"09",	--1681
		x"08",	--1682
		x"07",	--1683
		x"06",	--1684
		x"05",	--1685
		x"04",	--1686
		x"31",	--1687
		x"dc",	--1688
		x"81",	--1689
		x"04",	--1690
		x"81",	--1691
		x"06",	--1692
		x"81",	--1693
		x"00",	--1694
		x"81",	--1695
		x"02",	--1696
		x"0e",	--1697
		x"3e",	--1698
		x"18",	--1699
		x"0f",	--1700
		x"2f",	--1701
		x"b0",	--1702
		x"a4",	--1703
		x"0e",	--1704
		x"3e",	--1705
		x"10",	--1706
		x"0f",	--1707
		x"b0",	--1708
		x"a4",	--1709
		x"5f",	--1710
		x"18",	--1711
		x"6f",	--1712
		x"b6",	--1713
		x"5e",	--1714
		x"10",	--1715
		x"6e",	--1716
		x"d9",	--1717
		x"6f",	--1718
		x"ae",	--1719
		x"6e",	--1720
		x"e2",	--1721
		x"6f",	--1722
		x"ac",	--1723
		x"6e",	--1724
		x"d1",	--1725
		x"14",	--1726
		x"1c",	--1727
		x"15",	--1728
		x"1e",	--1729
		x"18",	--1730
		x"14",	--1731
		x"19",	--1732
		x"16",	--1733
		x"3c",	--1734
		x"20",	--1735
		x"0e",	--1736
		x"0f",	--1737
		x"06",	--1738
		x"07",	--1739
		x"81",	--1740
		x"20",	--1741
		x"81",	--1742
		x"22",	--1743
		x"0a",	--1744
		x"0b",	--1745
		x"81",	--1746
		x"20",	--1747
		x"08",	--1748
		x"08",	--1749
		x"09",	--1750
		x"12",	--1751
		x"05",	--1752
		x"04",	--1753
		x"b1",	--1754
		x"20",	--1755
		x"19",	--1756
		x"14",	--1757
		x"0d",	--1758
		x"0a",	--1759
		x"0b",	--1760
		x"0e",	--1761
		x"0f",	--1762
		x"1c",	--1763
		x"0d",	--1764
		x"0b",	--1765
		x"03",	--1766
		x"0b",	--1767
		x"0c",	--1768
		x"0d",	--1769
		x"0e",	--1770
		x"0f",	--1771
		x"06",	--1772
		x"07",	--1773
		x"09",	--1774
		x"e5",	--1775
		x"16",	--1776
		x"07",	--1777
		x"e2",	--1778
		x"0a",	--1779
		x"f5",	--1780
		x"f2",	--1781
		x"81",	--1782
		x"20",	--1783
		x"81",	--1784
		x"22",	--1785
		x"0c",	--1786
		x"1a",	--1787
		x"1a",	--1788
		x"1a",	--1789
		x"12",	--1790
		x"06",	--1791
		x"26",	--1792
		x"81",	--1793
		x"0a",	--1794
		x"5d",	--1795
		x"d1",	--1796
		x"11",	--1797
		x"19",	--1798
		x"83",	--1799
		x"c1",	--1800
		x"09",	--1801
		x"0c",	--1802
		x"3c",	--1803
		x"3f",	--1804
		x"00",	--1805
		x"18",	--1806
		x"1d",	--1807
		x"0a",	--1808
		x"3d",	--1809
		x"1a",	--1810
		x"20",	--1811
		x"1b",	--1812
		x"22",	--1813
		x"0c",	--1814
		x"0e",	--1815
		x"0f",	--1816
		x"0b",	--1817
		x"2a",	--1818
		x"0a",	--1819
		x"0b",	--1820
		x"3d",	--1821
		x"3f",	--1822
		x"00",	--1823
		x"f5",	--1824
		x"81",	--1825
		x"20",	--1826
		x"81",	--1827
		x"22",	--1828
		x"81",	--1829
		x"0a",	--1830
		x"0c",	--1831
		x"0d",	--1832
		x"3c",	--1833
		x"7f",	--1834
		x"0d",	--1835
		x"3c",	--1836
		x"40",	--1837
		x"44",	--1838
		x"81",	--1839
		x"0c",	--1840
		x"81",	--1841
		x"0e",	--1842
		x"f1",	--1843
		x"03",	--1844
		x"08",	--1845
		x"0f",	--1846
		x"3f",	--1847
		x"b0",	--1848
		x"c6",	--1849
		x"31",	--1850
		x"24",	--1851
		x"34",	--1852
		x"35",	--1853
		x"36",	--1854
		x"37",	--1855
		x"38",	--1856
		x"39",	--1857
		x"3a",	--1858
		x"3b",	--1859
		x"30",	--1860
		x"1e",	--1861
		x"0f",	--1862
		x"d3",	--1863
		x"3a",	--1864
		x"03",	--1865
		x"08",	--1866
		x"1e",	--1867
		x"10",	--1868
		x"1c",	--1869
		x"20",	--1870
		x"1d",	--1871
		x"22",	--1872
		x"12",	--1873
		x"0d",	--1874
		x"0c",	--1875
		x"06",	--1876
		x"07",	--1877
		x"06",	--1878
		x"37",	--1879
		x"00",	--1880
		x"81",	--1881
		x"20",	--1882
		x"81",	--1883
		x"22",	--1884
		x"12",	--1885
		x"0f",	--1886
		x"0e",	--1887
		x"1a",	--1888
		x"0f",	--1889
		x"e7",	--1890
		x"81",	--1891
		x"0a",	--1892
		x"a6",	--1893
		x"6e",	--1894
		x"36",	--1895
		x"5f",	--1896
		x"d1",	--1897
		x"11",	--1898
		x"19",	--1899
		x"20",	--1900
		x"c1",	--1901
		x"19",	--1902
		x"0f",	--1903
		x"3f",	--1904
		x"18",	--1905
		x"c5",	--1906
		x"0d",	--1907
		x"ba",	--1908
		x"0c",	--1909
		x"0d",	--1910
		x"3c",	--1911
		x"80",	--1912
		x"0d",	--1913
		x"0c",	--1914
		x"b3",	--1915
		x"0d",	--1916
		x"b1",	--1917
		x"81",	--1918
		x"20",	--1919
		x"03",	--1920
		x"81",	--1921
		x"22",	--1922
		x"ab",	--1923
		x"3e",	--1924
		x"40",	--1925
		x"0f",	--1926
		x"3e",	--1927
		x"80",	--1928
		x"3f",	--1929
		x"a4",	--1930
		x"4d",	--1931
		x"7b",	--1932
		x"4f",	--1933
		x"de",	--1934
		x"5f",	--1935
		x"d1",	--1936
		x"11",	--1937
		x"19",	--1938
		x"06",	--1939
		x"c1",	--1940
		x"11",	--1941
		x"0f",	--1942
		x"3f",	--1943
		x"10",	--1944
		x"9e",	--1945
		x"4f",	--1946
		x"f8",	--1947
		x"6f",	--1948
		x"f1",	--1949
		x"3f",	--1950
		x"5a",	--1951
		x"97",	--1952
		x"0b",	--1953
		x"0a",	--1954
		x"09",	--1955
		x"08",	--1956
		x"07",	--1957
		x"31",	--1958
		x"e8",	--1959
		x"81",	--1960
		x"04",	--1961
		x"81",	--1962
		x"06",	--1963
		x"81",	--1964
		x"00",	--1965
		x"81",	--1966
		x"02",	--1967
		x"0e",	--1968
		x"3e",	--1969
		x"10",	--1970
		x"0f",	--1971
		x"2f",	--1972
		x"b0",	--1973
		x"a4",	--1974
		x"0e",	--1975
		x"3e",	--1976
		x"0f",	--1977
		x"b0",	--1978
		x"a4",	--1979
		x"5f",	--1980
		x"10",	--1981
		x"6f",	--1982
		x"5d",	--1983
		x"5e",	--1984
		x"08",	--1985
		x"6e",	--1986
		x"82",	--1987
		x"d1",	--1988
		x"09",	--1989
		x"11",	--1990
		x"6f",	--1991
		x"58",	--1992
		x"6f",	--1993
		x"56",	--1994
		x"6e",	--1995
		x"6f",	--1996
		x"6e",	--1997
		x"4c",	--1998
		x"1d",	--1999
		x"12",	--2000
		x"1d",	--2001
		x"0a",	--2002
		x"81",	--2003
		x"12",	--2004
		x"1e",	--2005
		x"14",	--2006
		x"1f",	--2007
		x"16",	--2008
		x"18",	--2009
		x"0c",	--2010
		x"19",	--2011
		x"0e",	--2012
		x"0f",	--2013
		x"1e",	--2014
		x"0e",	--2015
		x"0f",	--2016
		x"3d",	--2017
		x"81",	--2018
		x"12",	--2019
		x"37",	--2020
		x"1f",	--2021
		x"0c",	--2022
		x"3d",	--2023
		x"00",	--2024
		x"0a",	--2025
		x"0b",	--2026
		x"0b",	--2027
		x"0a",	--2028
		x"0b",	--2029
		x"0e",	--2030
		x"0f",	--2031
		x"12",	--2032
		x"0d",	--2033
		x"0c",	--2034
		x"0e",	--2035
		x"0f",	--2036
		x"37",	--2037
		x"0b",	--2038
		x"0f",	--2039
		x"f7",	--2040
		x"f2",	--2041
		x"0e",	--2042
		x"f4",	--2043
		x"ef",	--2044
		x"09",	--2045
		x"e5",	--2046
		x"0e",	--2047
		x"e3",	--2048
		x"dd",	--2049
		x"0c",	--2050
		x"0d",	--2051
		x"3c",	--2052
		x"7f",	--2053
		x"0d",	--2054
		x"3c",	--2055
		x"40",	--2056
		x"1c",	--2057
		x"81",	--2058
		x"14",	--2059
		x"81",	--2060
		x"16",	--2061
		x"0f",	--2062
		x"3f",	--2063
		x"10",	--2064
		x"b0",	--2065
		x"c6",	--2066
		x"31",	--2067
		x"18",	--2068
		x"37",	--2069
		x"38",	--2070
		x"39",	--2071
		x"3a",	--2072
		x"3b",	--2073
		x"30",	--2074
		x"e1",	--2075
		x"10",	--2076
		x"0f",	--2077
		x"3f",	--2078
		x"10",	--2079
		x"f0",	--2080
		x"4f",	--2081
		x"fa",	--2082
		x"3f",	--2083
		x"5a",	--2084
		x"eb",	--2085
		x"0d",	--2086
		x"e2",	--2087
		x"0c",	--2088
		x"0d",	--2089
		x"3c",	--2090
		x"80",	--2091
		x"0d",	--2092
		x"0c",	--2093
		x"db",	--2094
		x"0d",	--2095
		x"d9",	--2096
		x"0e",	--2097
		x"02",	--2098
		x"0f",	--2099
		x"d5",	--2100
		x"3a",	--2101
		x"40",	--2102
		x"0b",	--2103
		x"3a",	--2104
		x"80",	--2105
		x"3b",	--2106
		x"ce",	--2107
		x"81",	--2108
		x"14",	--2109
		x"81",	--2110
		x"16",	--2111
		x"81",	--2112
		x"12",	--2113
		x"0f",	--2114
		x"3f",	--2115
		x"10",	--2116
		x"cb",	--2117
		x"0f",	--2118
		x"3f",	--2119
		x"c8",	--2120
		x"31",	--2121
		x"e8",	--2122
		x"81",	--2123
		x"04",	--2124
		x"81",	--2125
		x"06",	--2126
		x"81",	--2127
		x"00",	--2128
		x"81",	--2129
		x"02",	--2130
		x"0e",	--2131
		x"3e",	--2132
		x"10",	--2133
		x"0f",	--2134
		x"2f",	--2135
		x"b0",	--2136
		x"a4",	--2137
		x"0e",	--2138
		x"3e",	--2139
		x"0f",	--2140
		x"b0",	--2141
		x"a4",	--2142
		x"e1",	--2143
		x"10",	--2144
		x"0d",	--2145
		x"e1",	--2146
		x"08",	--2147
		x"0a",	--2148
		x"0e",	--2149
		x"3e",	--2150
		x"0f",	--2151
		x"3f",	--2152
		x"10",	--2153
		x"b0",	--2154
		x"c8",	--2155
		x"31",	--2156
		x"18",	--2157
		x"30",	--2158
		x"3f",	--2159
		x"fb",	--2160
		x"31",	--2161
		x"f4",	--2162
		x"81",	--2163
		x"00",	--2164
		x"81",	--2165
		x"02",	--2166
		x"0e",	--2167
		x"2e",	--2168
		x"0f",	--2169
		x"b0",	--2170
		x"a4",	--2171
		x"5f",	--2172
		x"04",	--2173
		x"6f",	--2174
		x"28",	--2175
		x"27",	--2176
		x"6f",	--2177
		x"07",	--2178
		x"1d",	--2179
		x"06",	--2180
		x"0d",	--2181
		x"21",	--2182
		x"3d",	--2183
		x"1f",	--2184
		x"09",	--2185
		x"c1",	--2186
		x"05",	--2187
		x"26",	--2188
		x"3e",	--2189
		x"3f",	--2190
		x"ff",	--2191
		x"31",	--2192
		x"0c",	--2193
		x"30",	--2194
		x"1e",	--2195
		x"08",	--2196
		x"1f",	--2197
		x"0a",	--2198
		x"3c",	--2199
		x"1e",	--2200
		x"4c",	--2201
		x"4d",	--2202
		x"7d",	--2203
		x"1f",	--2204
		x"0f",	--2205
		x"c1",	--2206
		x"05",	--2207
		x"ef",	--2208
		x"3e",	--2209
		x"3f",	--2210
		x"1e",	--2211
		x"0f",	--2212
		x"31",	--2213
		x"0c",	--2214
		x"30",	--2215
		x"0e",	--2216
		x"0f",	--2217
		x"31",	--2218
		x"0c",	--2219
		x"30",	--2220
		x"12",	--2221
		x"0f",	--2222
		x"0e",	--2223
		x"7d",	--2224
		x"fb",	--2225
		x"eb",	--2226
		x"0e",	--2227
		x"3f",	--2228
		x"00",	--2229
		x"31",	--2230
		x"0c",	--2231
		x"30",	--2232
		x"0b",	--2233
		x"0a",	--2234
		x"09",	--2235
		x"08",	--2236
		x"31",	--2237
		x"0a",	--2238
		x"0b",	--2239
		x"c1",	--2240
		x"01",	--2241
		x"0e",	--2242
		x"0d",	--2243
		x"0b",	--2244
		x"0b",	--2245
		x"e1",	--2246
		x"00",	--2247
		x"0f",	--2248
		x"b0",	--2249
		x"c6",	--2250
		x"31",	--2251
		x"38",	--2252
		x"39",	--2253
		x"3a",	--2254
		x"3b",	--2255
		x"30",	--2256
		x"f1",	--2257
		x"03",	--2258
		x"00",	--2259
		x"b1",	--2260
		x"1e",	--2261
		x"02",	--2262
		x"81",	--2263
		x"04",	--2264
		x"81",	--2265
		x"06",	--2266
		x"0e",	--2267
		x"0f",	--2268
		x"b0",	--2269
		x"54",	--2270
		x"3f",	--2271
		x"0f",	--2272
		x"18",	--2273
		x"e5",	--2274
		x"81",	--2275
		x"04",	--2276
		x"81",	--2277
		x"06",	--2278
		x"4e",	--2279
		x"7e",	--2280
		x"1f",	--2281
		x"06",	--2282
		x"3e",	--2283
		x"1e",	--2284
		x"0e",	--2285
		x"81",	--2286
		x"02",	--2287
		x"d7",	--2288
		x"91",	--2289
		x"04",	--2290
		x"04",	--2291
		x"91",	--2292
		x"06",	--2293
		x"06",	--2294
		x"7e",	--2295
		x"f8",	--2296
		x"f1",	--2297
		x"0e",	--2298
		x"3e",	--2299
		x"1e",	--2300
		x"1c",	--2301
		x"0d",	--2302
		x"48",	--2303
		x"78",	--2304
		x"1f",	--2305
		x"04",	--2306
		x"0c",	--2307
		x"0d",	--2308
		x"78",	--2309
		x"fc",	--2310
		x"3c",	--2311
		x"3d",	--2312
		x"0c",	--2313
		x"0d",	--2314
		x"18",	--2315
		x"09",	--2316
		x"0c",	--2317
		x"04",	--2318
		x"0d",	--2319
		x"02",	--2320
		x"08",	--2321
		x"09",	--2322
		x"7e",	--2323
		x"1f",	--2324
		x"0e",	--2325
		x"0d",	--2326
		x"0e",	--2327
		x"0d",	--2328
		x"0e",	--2329
		x"81",	--2330
		x"04",	--2331
		x"81",	--2332
		x"06",	--2333
		x"3e",	--2334
		x"1e",	--2335
		x"0e",	--2336
		x"81",	--2337
		x"02",	--2338
		x"a4",	--2339
		x"12",	--2340
		x"0b",	--2341
		x"0a",	--2342
		x"7e",	--2343
		x"fb",	--2344
		x"ec",	--2345
		x"0b",	--2346
		x"0a",	--2347
		x"09",	--2348
		x"1f",	--2349
		x"17",	--2350
		x"3e",	--2351
		x"00",	--2352
		x"2c",	--2353
		x"3a",	--2354
		x"18",	--2355
		x"0b",	--2356
		x"39",	--2357
		x"0c",	--2358
		x"0d",	--2359
		x"4f",	--2360
		x"4f",	--2361
		x"17",	--2362
		x"3c",	--2363
		x"62",	--2364
		x"6e",	--2365
		x"0f",	--2366
		x"0a",	--2367
		x"0b",	--2368
		x"0f",	--2369
		x"39",	--2370
		x"3a",	--2371
		x"3b",	--2372
		x"30",	--2373
		x"3f",	--2374
		x"00",	--2375
		x"0f",	--2376
		x"3a",	--2377
		x"0b",	--2378
		x"39",	--2379
		x"18",	--2380
		x"0c",	--2381
		x"0d",	--2382
		x"4f",	--2383
		x"4f",	--2384
		x"e9",	--2385
		x"12",	--2386
		x"0d",	--2387
		x"0c",	--2388
		x"7f",	--2389
		x"fb",	--2390
		x"e3",	--2391
		x"3a",	--2392
		x"10",	--2393
		x"0b",	--2394
		x"39",	--2395
		x"10",	--2396
		x"ef",	--2397
		x"3a",	--2398
		x"20",	--2399
		x"0b",	--2400
		x"09",	--2401
		x"ea",	--2402
		x"0b",	--2403
		x"0a",	--2404
		x"09",	--2405
		x"08",	--2406
		x"07",	--2407
		x"0d",	--2408
		x"1e",	--2409
		x"04",	--2410
		x"1f",	--2411
		x"06",	--2412
		x"5a",	--2413
		x"01",	--2414
		x"6c",	--2415
		x"6c",	--2416
		x"70",	--2417
		x"6c",	--2418
		x"6a",	--2419
		x"6c",	--2420
		x"36",	--2421
		x"0e",	--2422
		x"32",	--2423
		x"1b",	--2424
		x"02",	--2425
		x"3b",	--2426
		x"82",	--2427
		x"6d",	--2428
		x"3b",	--2429
		x"80",	--2430
		x"5e",	--2431
		x"0c",	--2432
		x"0d",	--2433
		x"3c",	--2434
		x"7f",	--2435
		x"0d",	--2436
		x"3c",	--2437
		x"40",	--2438
		x"40",	--2439
		x"3e",	--2440
		x"3f",	--2441
		x"0f",	--2442
		x"0f",	--2443
		x"4a",	--2444
		x"0d",	--2445
		x"3d",	--2446
		x"7f",	--2447
		x"12",	--2448
		x"0f",	--2449
		x"0e",	--2450
		x"12",	--2451
		x"0f",	--2452
		x"0e",	--2453
		x"12",	--2454
		x"0f",	--2455
		x"0e",	--2456
		x"12",	--2457
		x"0f",	--2458
		x"0e",	--2459
		x"12",	--2460
		x"0f",	--2461
		x"0e",	--2462
		x"12",	--2463
		x"0f",	--2464
		x"0e",	--2465
		x"12",	--2466
		x"0f",	--2467
		x"0e",	--2468
		x"3e",	--2469
		x"3f",	--2470
		x"7f",	--2471
		x"4d",	--2472
		x"05",	--2473
		x"0f",	--2474
		x"cc",	--2475
		x"4d",	--2476
		x"0e",	--2477
		x"0f",	--2478
		x"4d",	--2479
		x"0d",	--2480
		x"0d",	--2481
		x"0d",	--2482
		x"0d",	--2483
		x"0d",	--2484
		x"0d",	--2485
		x"0d",	--2486
		x"0c",	--2487
		x"3c",	--2488
		x"7f",	--2489
		x"0c",	--2490
		x"4f",	--2491
		x"0f",	--2492
		x"0f",	--2493
		x"0f",	--2494
		x"0d",	--2495
		x"0d",	--2496
		x"0f",	--2497
		x"37",	--2498
		x"38",	--2499
		x"39",	--2500
		x"3a",	--2501
		x"3b",	--2502
		x"30",	--2503
		x"0d",	--2504
		x"be",	--2505
		x"0c",	--2506
		x"0d",	--2507
		x"3c",	--2508
		x"80",	--2509
		x"0d",	--2510
		x"0c",	--2511
		x"02",	--2512
		x"0d",	--2513
		x"b8",	--2514
		x"3e",	--2515
		x"40",	--2516
		x"0f",	--2517
		x"b4",	--2518
		x"12",	--2519
		x"0f",	--2520
		x"0e",	--2521
		x"0d",	--2522
		x"3d",	--2523
		x"80",	--2524
		x"b2",	--2525
		x"7d",	--2526
		x"0e",	--2527
		x"0f",	--2528
		x"cd",	--2529
		x"0e",	--2530
		x"3f",	--2531
		x"10",	--2532
		x"3e",	--2533
		x"3f",	--2534
		x"7f",	--2535
		x"7d",	--2536
		x"c5",	--2537
		x"37",	--2538
		x"82",	--2539
		x"07",	--2540
		x"37",	--2541
		x"1a",	--2542
		x"4f",	--2543
		x"0c",	--2544
		x"0d",	--2545
		x"4b",	--2546
		x"7b",	--2547
		x"1f",	--2548
		x"05",	--2549
		x"12",	--2550
		x"0d",	--2551
		x"0c",	--2552
		x"7b",	--2553
		x"fb",	--2554
		x"18",	--2555
		x"09",	--2556
		x"77",	--2557
		x"1f",	--2558
		x"04",	--2559
		x"08",	--2560
		x"09",	--2561
		x"77",	--2562
		x"fc",	--2563
		x"38",	--2564
		x"39",	--2565
		x"08",	--2566
		x"09",	--2567
		x"1e",	--2568
		x"0f",	--2569
		x"08",	--2570
		x"04",	--2571
		x"09",	--2572
		x"02",	--2573
		x"0e",	--2574
		x"0f",	--2575
		x"08",	--2576
		x"09",	--2577
		x"08",	--2578
		x"09",	--2579
		x"0e",	--2580
		x"0f",	--2581
		x"3e",	--2582
		x"7f",	--2583
		x"0f",	--2584
		x"3e",	--2585
		x"40",	--2586
		x"26",	--2587
		x"38",	--2588
		x"3f",	--2589
		x"09",	--2590
		x"0e",	--2591
		x"0f",	--2592
		x"12",	--2593
		x"0f",	--2594
		x"0e",	--2595
		x"12",	--2596
		x"0f",	--2597
		x"0e",	--2598
		x"12",	--2599
		x"0f",	--2600
		x"0e",	--2601
		x"12",	--2602
		x"0f",	--2603
		x"0e",	--2604
		x"12",	--2605
		x"0f",	--2606
		x"0e",	--2607
		x"12",	--2608
		x"0f",	--2609
		x"0e",	--2610
		x"12",	--2611
		x"0f",	--2612
		x"0e",	--2613
		x"3e",	--2614
		x"3f",	--2615
		x"7f",	--2616
		x"5d",	--2617
		x"39",	--2618
		x"00",	--2619
		x"72",	--2620
		x"4d",	--2621
		x"70",	--2622
		x"08",	--2623
		x"09",	--2624
		x"da",	--2625
		x"0f",	--2626
		x"d8",	--2627
		x"0e",	--2628
		x"0f",	--2629
		x"3e",	--2630
		x"80",	--2631
		x"0f",	--2632
		x"0e",	--2633
		x"04",	--2634
		x"38",	--2635
		x"40",	--2636
		x"09",	--2637
		x"d0",	--2638
		x"0f",	--2639
		x"ce",	--2640
		x"f9",	--2641
		x"0b",	--2642
		x"0a",	--2643
		x"2a",	--2644
		x"5b",	--2645
		x"02",	--2646
		x"3b",	--2647
		x"7f",	--2648
		x"1d",	--2649
		x"02",	--2650
		x"12",	--2651
		x"0d",	--2652
		x"12",	--2653
		x"0d",	--2654
		x"12",	--2655
		x"0d",	--2656
		x"12",	--2657
		x"0d",	--2658
		x"12",	--2659
		x"0d",	--2660
		x"12",	--2661
		x"0d",	--2662
		x"12",	--2663
		x"0d",	--2664
		x"4d",	--2665
		x"5f",	--2666
		x"03",	--2667
		x"3f",	--2668
		x"80",	--2669
		x"0f",	--2670
		x"0f",	--2671
		x"ce",	--2672
		x"01",	--2673
		x"0d",	--2674
		x"2d",	--2675
		x"0a",	--2676
		x"51",	--2677
		x"be",	--2678
		x"82",	--2679
		x"02",	--2680
		x"0c",	--2681
		x"0d",	--2682
		x"0c",	--2683
		x"0d",	--2684
		x"0c",	--2685
		x"0d",	--2686
		x"0c",	--2687
		x"0d",	--2688
		x"0c",	--2689
		x"0d",	--2690
		x"0c",	--2691
		x"0d",	--2692
		x"0c",	--2693
		x"0d",	--2694
		x"0c",	--2695
		x"0d",	--2696
		x"fe",	--2697
		x"03",	--2698
		x"00",	--2699
		x"3d",	--2700
		x"00",	--2701
		x"0b",	--2702
		x"3f",	--2703
		x"81",	--2704
		x"0c",	--2705
		x"0d",	--2706
		x"0a",	--2707
		x"3f",	--2708
		x"3d",	--2709
		x"00",	--2710
		x"f9",	--2711
		x"8e",	--2712
		x"02",	--2713
		x"8e",	--2714
		x"04",	--2715
		x"8e",	--2716
		x"06",	--2717
		x"3a",	--2718
		x"3b",	--2719
		x"30",	--2720
		x"3d",	--2721
		x"ff",	--2722
		x"2a",	--2723
		x"3d",	--2724
		x"81",	--2725
		x"8e",	--2726
		x"02",	--2727
		x"fe",	--2728
		x"03",	--2729
		x"00",	--2730
		x"0c",	--2731
		x"0d",	--2732
		x"0c",	--2733
		x"0d",	--2734
		x"0c",	--2735
		x"0d",	--2736
		x"0c",	--2737
		x"0d",	--2738
		x"0c",	--2739
		x"0d",	--2740
		x"0c",	--2741
		x"0d",	--2742
		x"0c",	--2743
		x"0d",	--2744
		x"0c",	--2745
		x"0d",	--2746
		x"0a",	--2747
		x"0b",	--2748
		x"0a",	--2749
		x"3b",	--2750
		x"00",	--2751
		x"8e",	--2752
		x"04",	--2753
		x"8e",	--2754
		x"06",	--2755
		x"3a",	--2756
		x"3b",	--2757
		x"30",	--2758
		x"0b",	--2759
		x"ad",	--2760
		x"ee",	--2761
		x"00",	--2762
		x"3a",	--2763
		x"3b",	--2764
		x"30",	--2765
		x"0a",	--2766
		x"0c",	--2767
		x"0c",	--2768
		x"0d",	--2769
		x"0c",	--2770
		x"3d",	--2771
		x"10",	--2772
		x"0c",	--2773
		x"02",	--2774
		x"0d",	--2775
		x"08",	--2776
		x"de",	--2777
		x"00",	--2778
		x"e4",	--2779
		x"0b",	--2780
		x"f2",	--2781
		x"ee",	--2782
		x"00",	--2783
		x"e3",	--2784
		x"ce",	--2785
		x"00",	--2786
		x"dc",	--2787
		x"0b",	--2788
		x"6d",	--2789
		x"6d",	--2790
		x"12",	--2791
		x"6c",	--2792
		x"6c",	--2793
		x"0f",	--2794
		x"6d",	--2795
		x"41",	--2796
		x"6c",	--2797
		x"11",	--2798
		x"6d",	--2799
		x"0d",	--2800
		x"6c",	--2801
		x"14",	--2802
		x"5d",	--2803
		x"01",	--2804
		x"5d",	--2805
		x"01",	--2806
		x"14",	--2807
		x"4d",	--2808
		x"09",	--2809
		x"1e",	--2810
		x"0f",	--2811
		x"3b",	--2812
		x"30",	--2813
		x"6c",	--2814
		x"28",	--2815
		x"ce",	--2816
		x"01",	--2817
		x"f7",	--2818
		x"3e",	--2819
		x"0f",	--2820
		x"3b",	--2821
		x"30",	--2822
		x"cf",	--2823
		x"01",	--2824
		x"f0",	--2825
		x"3e",	--2826
		x"f8",	--2827
		x"1b",	--2828
		x"02",	--2829
		x"1c",	--2830
		x"02",	--2831
		x"0c",	--2832
		x"e6",	--2833
		x"0b",	--2834
		x"16",	--2835
		x"1b",	--2836
		x"04",	--2837
		x"1f",	--2838
		x"06",	--2839
		x"1c",	--2840
		x"04",	--2841
		x"1e",	--2842
		x"06",	--2843
		x"0e",	--2844
		x"da",	--2845
		x"0f",	--2846
		x"02",	--2847
		x"0c",	--2848
		x"d6",	--2849
		x"0f",	--2850
		x"06",	--2851
		x"0e",	--2852
		x"02",	--2853
		x"0b",	--2854
		x"02",	--2855
		x"0e",	--2856
		x"d1",	--2857
		x"4d",	--2858
		x"ce",	--2859
		x"3e",	--2860
		x"d6",	--2861
		x"6c",	--2862
		x"d7",	--2863
		x"5e",	--2864
		x"01",	--2865
		x"5f",	--2866
		x"01",	--2867
		x"0e",	--2868
		x"c5",	--2869
		x"0d",	--2870
		x"0f",	--2871
		x"04",	--2872
		x"3d",	--2873
		x"03",	--2874
		x"3f",	--2875
		x"1f",	--2876
		x"0e",	--2877
		x"03",	--2878
		x"5d",	--2879
		x"3e",	--2880
		x"1e",	--2881
		x"0d",	--2882
		x"b0",	--2883
		x"f2",	--2884
		x"3d",	--2885
		x"6d",	--2886
		x"02",	--2887
		x"3e",	--2888
		x"1e",	--2889
		x"5d",	--2890
		x"02",	--2891
		x"3f",	--2892
		x"1f",	--2893
		x"30",	--2894
		x"b0",	--2895
		x"6c",	--2896
		x"0f",	--2897
		x"30",	--2898
		x"0b",	--2899
		x"0b",	--2900
		x"0f",	--2901
		x"06",	--2902
		x"3b",	--2903
		x"03",	--2904
		x"3e",	--2905
		x"3f",	--2906
		x"1e",	--2907
		x"0f",	--2908
		x"0d",	--2909
		x"05",	--2910
		x"5b",	--2911
		x"3c",	--2912
		x"3d",	--2913
		x"1c",	--2914
		x"0d",	--2915
		x"b0",	--2916
		x"14",	--2917
		x"6b",	--2918
		x"04",	--2919
		x"3c",	--2920
		x"3d",	--2921
		x"1c",	--2922
		x"0d",	--2923
		x"5b",	--2924
		x"04",	--2925
		x"3e",	--2926
		x"3f",	--2927
		x"1e",	--2928
		x"0f",	--2929
		x"3b",	--2930
		x"30",	--2931
		x"b0",	--2932
		x"a6",	--2933
		x"0e",	--2934
		x"0f",	--2935
		x"30",	--2936
		x"7c",	--2937
		x"10",	--2938
		x"0d",	--2939
		x"0e",	--2940
		x"0f",	--2941
		x"0e",	--2942
		x"0e",	--2943
		x"02",	--2944
		x"0e",	--2945
		x"1f",	--2946
		x"1c",	--2947
		x"f8",	--2948
		x"30",	--2949
		x"b0",	--2950
		x"f2",	--2951
		x"0f",	--2952
		x"30",	--2953
		x"0b",	--2954
		x"0a",	--2955
		x"09",	--2956
		x"79",	--2957
		x"20",	--2958
		x"0a",	--2959
		x"0b",	--2960
		x"0c",	--2961
		x"0d",	--2962
		x"0e",	--2963
		x"0f",	--2964
		x"0c",	--2965
		x"0d",	--2966
		x"0d",	--2967
		x"06",	--2968
		x"02",	--2969
		x"0c",	--2970
		x"03",	--2971
		x"0c",	--2972
		x"0d",	--2973
		x"1e",	--2974
		x"19",	--2975
		x"f2",	--2976
		x"39",	--2977
		x"3a",	--2978
		x"3b",	--2979
		x"30",	--2980
		x"b0",	--2981
		x"14",	--2982
		x"0e",	--2983
		x"0f",	--2984
		x"30",	--2985
		x"00",	--2986
		x"32",	--2987
		x"f0",	--2988
		x"fd",	--2989
		x"57",	--2990
		x"69",	--2991
		x"69",	--2992
		x"67",	--2993
		x"66",	--2994
		x"72",	--2995
		x"61",	--2996
		x"6e",	--2997
		x"77",	--2998
		x"2e",	--2999
		x"69",	--3000
		x"20",	--3001
		x"69",	--3002
		x"65",	--3003
		x"0a",	--3004
		x"57",	--3005
		x"20",	--3006
		x"68",	--3007
		x"75",	--3008
		x"64",	--3009
		x"6e",	--3010
		x"74",	--3011
		x"73",	--3012
		x"65",	--3013
		x"74",	--3014
		x"61",	--3015
		x"0d",	--3016
		x"00",	--3017
		x"6f",	--3018
		x"72",	--3019
		x"63",	--3020
		x"20",	--3021
		x"73",	--3022
		x"67",	--3023
		x"3a",	--3024
		x"0a",	--3025
		x"09",	--3026
		x"63",	--3027
		x"4c",	--3028
		x"46",	--3029
		x"20",	--3030
		x"49",	--3031
		x"48",	--3032
		x"0d",	--3033
		x"00",	--3034
		x"6f",	--3035
		x"65",	--3036
		x"68",	--3037
		x"6e",	--3038
		x"20",	--3039
		x"65",	--3040
		x"74",	--3041
		x"74",	--3042
		x"72",	--3043
		x"69",	--3044
		x"6c",	--3045
		x"20",	--3046
		x"72",	--3047
		x"6e",	--3048
		x"0d",	--3049
		x"00",	--3050
		x"0a",	--3051
		x"3d",	--3052
		x"3d",	--3053
		x"3d",	--3054
		x"4d",	--3055
		x"72",	--3056
		x"65",	--3057
		x"20",	--3058
		x"43",	--3059
		x"20",	--3060
		x"3d",	--3061
		x"3d",	--3062
		x"3d",	--3063
		x"0a",	--3064
		x"3e",	--3065
		x"00",	--3066
		x"0a",	--3067
		x"3a",	--3068
		x"73",	--3069
		x"0a",	--3070
		x"08",	--3071
		x"08",	--3072
		x"25",	--3073
		x"00",	--3074
		x"72",	--3075
		x"74",	--3076
		x"0a",	--3077
		x"00",	--3078
		x"6f",	--3079
		x"72",	--3080
		x"63",	--3081
		x"20",	--3082
		x"73",	--3083
		x"67",	--3084
		x"3a",	--3085
		x"0a",	--3086
		x"09",	--3087
		x"63",	--3088
		x"52",	--3089
		x"47",	--3090
		x"53",	--3091
		x"45",	--3092
		x"20",	--3093
		x"41",	--3094
		x"55",	--3095
		x"0d",	--3096
		x"00",	--3097
		x"6f",	--3098
		x"65",	--3099
		x"68",	--3100
		x"6e",	--3101
		x"20",	--3102
		x"65",	--3103
		x"74",	--3104
		x"74",	--3105
		x"72",	--3106
		x"69",	--3107
		x"6c",	--3108
		x"20",	--3109
		x"72",	--3110
		x"6e",	--3111
		x"0d",	--3112
		x"00",	--3113
		x"3d",	--3114
		x"64",	--3115
		x"76",	--3116
		x"25",	--3117
		x"0d",	--3118
		x"00",	--3119
		x"65",	--3120
		x"64",	--3121
		x"0d",	--3122
		x"09",	--3123
		x"63",	--3124
		x"52",	--3125
		x"47",	--3126
		x"53",	--3127
		x"45",	--3128
		x"0d",	--3129
		x"00",	--3130
		x"63",	--3131
		x"69",	--3132
		x"20",	--3133
		x"6f",	--3134
		x"20",	--3135
		x"20",	--3136
		x"75",	--3137
		x"62",	--3138
		x"72",	--3139
		x"0a",	--3140
		x"25",	--3141
		x"3a",	--3142
		x"6e",	--3143
		x"20",	--3144
		x"75",	--3145
		x"68",	--3146
		x"63",	--3147
		x"6d",	--3148
		x"61",	--3149
		x"64",	--3150
		x"0a",	--3151
		x"f6",	--3152
		x"24",	--3153
		x"24",	--3154
		x"24",	--3155
		x"24",	--3156
		x"24",	--3157
		x"24",	--3158
		x"24",	--3159
		x"24",	--3160
		x"24",	--3161
		x"24",	--3162
		x"24",	--3163
		x"24",	--3164
		x"24",	--3165
		x"24",	--3166
		x"24",	--3167
		x"24",	--3168
		x"24",	--3169
		x"24",	--3170
		x"24",	--3171
		x"24",	--3172
		x"24",	--3173
		x"24",	--3174
		x"24",	--3175
		x"24",	--3176
		x"24",	--3177
		x"24",	--3178
		x"24",	--3179
		x"24",	--3180
		x"e8",	--3181
		x"24",	--3182
		x"24",	--3183
		x"24",	--3184
		x"24",	--3185
		x"24",	--3186
		x"24",	--3187
		x"24",	--3188
		x"24",	--3189
		x"24",	--3190
		x"24",	--3191
		x"24",	--3192
		x"24",	--3193
		x"24",	--3194
		x"24",	--3195
		x"24",	--3196
		x"24",	--3197
		x"24",	--3198
		x"24",	--3199
		x"24",	--3200
		x"24",	--3201
		x"24",	--3202
		x"24",	--3203
		x"24",	--3204
		x"24",	--3205
		x"24",	--3206
		x"24",	--3207
		x"24",	--3208
		x"24",	--3209
		x"24",	--3210
		x"24",	--3211
		x"24",	--3212
		x"da",	--3213
		x"cc",	--3214
		x"be",	--3215
		x"24",	--3216
		x"24",	--3217
		x"24",	--3218
		x"24",	--3219
		x"24",	--3220
		x"24",	--3221
		x"24",	--3222
		x"a6",	--3223
		x"24",	--3224
		x"94",	--3225
		x"24",	--3226
		x"24",	--3227
		x"24",	--3228
		x"24",	--3229
		x"78",	--3230
		x"24",	--3231
		x"24",	--3232
		x"24",	--3233
		x"6a",	--3234
		x"58",	--3235
		x"30",	--3236
		x"32",	--3237
		x"34",	--3238
		x"36",	--3239
		x"38",	--3240
		x"61",	--3241
		x"63",	--3242
		x"65",	--3243
		x"00",	--3244
		x"00",	--3245
		x"00",	--3246
		x"00",	--3247
		x"00",	--3248
		x"00",	--3249
		x"02",	--3250
		x"03",	--3251
		x"03",	--3252
		x"04",	--3253
		x"04",	--3254
		x"04",	--3255
		x"04",	--3256
		x"05",	--3257
		x"05",	--3258
		x"05",	--3259
		x"05",	--3260
		x"05",	--3261
		x"05",	--3262
		x"05",	--3263
		x"05",	--3264
		x"06",	--3265
		x"06",	--3266
		x"06",	--3267
		x"06",	--3268
		x"06",	--3269
		x"06",	--3270
		x"06",	--3271
		x"06",	--3272
		x"06",	--3273
		x"06",	--3274
		x"06",	--3275
		x"06",	--3276
		x"06",	--3277
		x"06",	--3278
		x"06",	--3279
		x"06",	--3280
		x"07",	--3281
		x"07",	--3282
		x"07",	--3283
		x"07",	--3284
		x"07",	--3285
		x"07",	--3286
		x"07",	--3287
		x"07",	--3288
		x"07",	--3289
		x"07",	--3290
		x"07",	--3291
		x"07",	--3292
		x"07",	--3293
		x"07",	--3294
		x"07",	--3295
		x"07",	--3296
		x"07",	--3297
		x"07",	--3298
		x"07",	--3299
		x"07",	--3300
		x"07",	--3301
		x"07",	--3302
		x"07",	--3303
		x"07",	--3304
		x"07",	--3305
		x"07",	--3306
		x"07",	--3307
		x"07",	--3308
		x"07",	--3309
		x"07",	--3310
		x"07",	--3311
		x"07",	--3312
		x"08",	--3313
		x"08",	--3314
		x"08",	--3315
		x"08",	--3316
		x"08",	--3317
		x"08",	--3318
		x"08",	--3319
		x"08",	--3320
		x"08",	--3321
		x"08",	--3322
		x"08",	--3323
		x"08",	--3324
		x"08",	--3325
		x"08",	--3326
		x"08",	--3327
		x"08",	--3328
		x"08",	--3329
		x"08",	--3330
		x"08",	--3331
		x"08",	--3332
		x"08",	--3333
		x"08",	--3334
		x"08",	--3335
		x"08",	--3336
		x"08",	--3337
		x"08",	--3338
		x"08",	--3339
		x"08",	--3340
		x"08",	--3341
		x"08",	--3342
		x"08",	--3343
		x"08",	--3344
		x"08",	--3345
		x"08",	--3346
		x"08",	--3347
		x"08",	--3348
		x"08",	--3349
		x"08",	--3350
		x"08",	--3351
		x"08",	--3352
		x"08",	--3353
		x"08",	--3354
		x"08",	--3355
		x"08",	--3356
		x"08",	--3357
		x"08",	--3358
		x"08",	--3359
		x"08",	--3360
		x"08",	--3361
		x"08",	--3362
		x"08",	--3363
		x"08",	--3364
		x"08",	--3365
		x"08",	--3366
		x"08",	--3367
		x"08",	--3368
		x"08",	--3369
		x"08",	--3370
		x"08",	--3371
		x"08",	--3372
		x"08",	--3373
		x"08",	--3374
		x"08",	--3375
		x"08",	--3376
		x"ff",	--3377
		x"ff",	--3378
		x"ff",	--3379
		x"ff",	--3380
		x"ff",	--3381
		x"ff",	--3382
		x"ff",	--3383
		x"ff",	--3384
		x"ff",	--3385
		x"ff",	--3386
		x"ff",	--3387
		x"ff",	--3388
		x"ff",	--3389
		x"ff",	--3390
		x"ff",	--3391
		x"ff",	--3392
		x"ff",	--3393
		x"ff",	--3394
		x"ff",	--3395
		x"ff",	--3396
		x"ff",	--3397
		x"ff",	--3398
		x"ff",	--3399
		x"ff",	--3400
		x"ff",	--3401
		x"ff",	--3402
		x"ff",	--3403
		x"ff",	--3404
		x"ff",	--3405
		x"ff",	--3406
		x"ff",	--3407
		x"ff",	--3408
		x"ff",	--3409
		x"ff",	--3410
		x"ff",	--3411
		x"ff",	--3412
		x"ff",	--3413
		x"ff",	--3414
		x"ff",	--3415
		x"ff",	--3416
		x"ff",	--3417
		x"ff",	--3418
		x"ff",	--3419
		x"ff",	--3420
		x"ff",	--3421
		x"ff",	--3422
		x"ff",	--3423
		x"ff",	--3424
		x"ff",	--3425
		x"ff",	--3426
		x"ff",	--3427
		x"ff",	--3428
		x"ff",	--3429
		x"ff",	--3430
		x"ff",	--3431
		x"ff",	--3432
		x"ff",	--3433
		x"ff",	--3434
		x"ff",	--3435
		x"ff",	--3436
		x"ff",	--3437
		x"ff",	--3438
		x"ff",	--3439
		x"ff",	--3440
		x"ff",	--3441
		x"ff",	--3442
		x"ff",	--3443
		x"ff",	--3444
		x"ff",	--3445
		x"ff",	--3446
		x"ff",	--3447
		x"ff",	--3448
		x"ff",	--3449
		x"ff",	--3450
		x"ff",	--3451
		x"ff",	--3452
		x"ff",	--3453
		x"ff",	--3454
		x"ff",	--3455
		x"ff",	--3456
		x"ff",	--3457
		x"ff",	--3458
		x"ff",	--3459
		x"ff",	--3460
		x"ff",	--3461
		x"ff",	--3462
		x"ff",	--3463
		x"ff",	--3464
		x"ff",	--3465
		x"ff",	--3466
		x"ff",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"a2",	--4080
		x"a2",	--4081
		x"a2",	--4082
		x"a2",	--4083
		x"a2",	--4084
		x"a2",	--4085
		x"a2",	--4086
		x"00",	--4087
		x"a2",	--4088
		x"a2",	--4089
		x"a2",	--4090
		x"a2",	--4091
		x"a2",	--4092
		x"a2",	--4093
		x"a2",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"03",	--5
		x"40",	--6
		x"06",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"03",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fa",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"01",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"03",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"25",	--41
		x"43",	--42
		x"12",	--43
		x"e9",	--44
		x"12",	--45
		x"e5",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"f7",	--50
		x"12",	--51
		x"e8",	--52
		x"53",	--53
		x"40",	--54
		x"e2",	--55
		x"40",	--56
		x"00",	--57
		x"12",	--58
		x"e5",	--59
		x"40",	--60
		x"e3",	--61
		x"40",	--62
		x"00",	--63
		x"12",	--64
		x"e5",	--65
		x"40",	--66
		x"e1",	--67
		x"40",	--68
		x"00",	--69
		x"12",	--70
		x"e5",	--71
		x"40",	--72
		x"e1",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"e5",	--77
		x"43",	--78
		x"40",	--79
		x"4e",	--80
		x"40",	--81
		x"01",	--82
		x"41",	--83
		x"50",	--84
		x"00",	--85
		x"12",	--86
		x"e4",	--87
		x"41",	--88
		x"50",	--89
		x"00",	--90
		x"12",	--91
		x"e5",	--92
		x"43",	--93
		x"40",	--94
		x"4e",	--95
		x"40",	--96
		x"01",	--97
		x"41",	--98
		x"12",	--99
		x"e4",	--100
		x"41",	--101
		x"12",	--102
		x"e5",	--103
		x"41",	--104
		x"41",	--105
		x"50",	--106
		x"00",	--107
		x"12",	--108
		x"e1",	--109
		x"40",	--110
		x"ff",	--111
		x"00",	--112
		x"d2",	--113
		x"43",	--114
		x"12",	--115
		x"f7",	--116
		x"12",	--117
		x"e8",	--118
		x"53",	--119
		x"43",	--120
		x"d0",	--121
		x"00",	--122
		x"53",	--123
		x"90",	--124
		x"00",	--125
		x"24",	--126
		x"43",	--127
		x"4b",	--128
		x"f0",	--129
		x"00",	--130
		x"24",	--131
		x"5f",	--132
		x"53",	--133
		x"23",	--134
		x"4f",	--135
		x"3c",	--136
		x"43",	--137
		x"43",	--138
		x"4f",	--139
		x"00",	--140
		x"12",	--141
		x"e9",	--142
		x"93",	--143
		x"27",	--144
		x"12",	--145
		x"e9",	--146
		x"92",	--147
		x"24",	--148
		x"90",	--149
		x"00",	--150
		x"20",	--151
		x"12",	--152
		x"f7",	--153
		x"12",	--154
		x"e8",	--155
		x"53",	--156
		x"40",	--157
		x"00",	--158
		x"51",	--159
		x"5f",	--160
		x"43",	--161
		x"00",	--162
		x"12",	--163
		x"12",	--164
		x"f7",	--165
		x"12",	--166
		x"e8",	--167
		x"52",	--168
		x"41",	--169
		x"50",	--170
		x"00",	--171
		x"41",	--172
		x"00",	--173
		x"12",	--174
		x"e5",	--175
		x"3f",	--176
		x"93",	--177
		x"27",	--178
		x"53",	--179
		x"12",	--180
		x"f7",	--181
		x"12",	--182
		x"e8",	--183
		x"53",	--184
		x"3f",	--185
		x"90",	--186
		x"00",	--187
		x"2f",	--188
		x"4f",	--189
		x"11",	--190
		x"12",	--191
		x"12",	--192
		x"f8",	--193
		x"4f",	--194
		x"00",	--195
		x"12",	--196
		x"e8",	--197
		x"52",	--198
		x"40",	--199
		x"00",	--200
		x"51",	--201
		x"5a",	--202
		x"41",	--203
		x"00",	--204
		x"4f",	--205
		x"00",	--206
		x"53",	--207
		x"3f",	--208
		x"40",	--209
		x"f7",	--210
		x"40",	--211
		x"e0",	--212
		x"01",	--213
		x"42",	--214
		x"01",	--215
		x"40",	--216
		x"02",	--217
		x"01",	--218
		x"12",	--219
		x"f7",	--220
		x"12",	--221
		x"e8",	--222
		x"43",	--223
		x"01",	--224
		x"40",	--225
		x"f7",	--226
		x"00",	--227
		x"12",	--228
		x"e8",	--229
		x"53",	--230
		x"43",	--231
		x"41",	--232
		x"4f",	--233
		x"02",	--234
		x"4e",	--235
		x"02",	--236
		x"41",	--237
		x"82",	--238
		x"90",	--239
		x"00",	--240
		x"00",	--241
		x"20",	--242
		x"93",	--243
		x"00",	--244
		x"24",	--245
		x"41",	--246
		x"4f",	--247
		x"53",	--248
		x"41",	--249
		x"52",	--250
		x"12",	--251
		x"e3",	--252
		x"93",	--253
		x"00",	--254
		x"24",	--255
		x"41",	--256
		x"4f",	--257
		x"41",	--258
		x"53",	--259
		x"12",	--260
		x"e3",	--261
		x"93",	--262
		x"00",	--263
		x"24",	--264
		x"41",	--265
		x"00",	--266
		x"43",	--267
		x"12",	--268
		x"f1",	--269
		x"43",	--270
		x"40",	--271
		x"42",	--272
		x"12",	--273
		x"ef",	--274
		x"4e",	--275
		x"4f",	--276
		x"42",	--277
		x"02",	--278
		x"12",	--279
		x"e5",	--280
		x"41",	--281
		x"00",	--282
		x"43",	--283
		x"12",	--284
		x"f1",	--285
		x"43",	--286
		x"40",	--287
		x"42",	--288
		x"12",	--289
		x"ef",	--290
		x"4e",	--291
		x"4f",	--292
		x"42",	--293
		x"02",	--294
		x"12",	--295
		x"e5",	--296
		x"43",	--297
		x"52",	--298
		x"41",	--299
		x"12",	--300
		x"f7",	--301
		x"4f",	--302
		x"00",	--303
		x"12",	--304
		x"e8",	--305
		x"41",	--306
		x"00",	--307
		x"4f",	--308
		x"11",	--309
		x"4f",	--310
		x"00",	--311
		x"12",	--312
		x"f7",	--313
		x"12",	--314
		x"e8",	--315
		x"52",	--316
		x"43",	--317
		x"52",	--318
		x"41",	--319
		x"12",	--320
		x"f7",	--321
		x"12",	--322
		x"e8",	--323
		x"53",	--324
		x"43",	--325
		x"3f",	--326
		x"12",	--327
		x"50",	--328
		x"ff",	--329
		x"4f",	--330
		x"12",	--331
		x"f8",	--332
		x"12",	--333
		x"e8",	--334
		x"53",	--335
		x"90",	--336
		x"00",	--337
		x"00",	--338
		x"20",	--339
		x"93",	--340
		x"00",	--341
		x"24",	--342
		x"41",	--343
		x"4b",	--344
		x"53",	--345
		x"41",	--346
		x"52",	--347
		x"12",	--348
		x"e3",	--349
		x"93",	--350
		x"00",	--351
		x"24",	--352
		x"41",	--353
		x"4f",	--354
		x"41",	--355
		x"53",	--356
		x"12",	--357
		x"e3",	--358
		x"93",	--359
		x"00",	--360
		x"24",	--361
		x"12",	--362
		x"00",	--363
		x"12",	--364
		x"00",	--365
		x"12",	--366
		x"f8",	--367
		x"12",	--368
		x"e8",	--369
		x"50",	--370
		x"00",	--371
		x"41",	--372
		x"00",	--373
		x"41",	--374
		x"00",	--375
		x"00",	--376
		x"43",	--377
		x"50",	--378
		x"00",	--379
		x"41",	--380
		x"41",	--381
		x"12",	--382
		x"f8",	--383
		x"12",	--384
		x"e8",	--385
		x"4b",	--386
		x"11",	--387
		x"4f",	--388
		x"00",	--389
		x"12",	--390
		x"f8",	--391
		x"12",	--392
		x"e8",	--393
		x"52",	--394
		x"43",	--395
		x"50",	--396
		x"00",	--397
		x"41",	--398
		x"41",	--399
		x"12",	--400
		x"f8",	--401
		x"12",	--402
		x"e8",	--403
		x"53",	--404
		x"43",	--405
		x"3f",	--406
		x"12",	--407
		x"82",	--408
		x"4f",	--409
		x"12",	--410
		x"f8",	--411
		x"12",	--412
		x"e8",	--413
		x"53",	--414
		x"90",	--415
		x"00",	--416
		x"00",	--417
		x"20",	--418
		x"93",	--419
		x"00",	--420
		x"24",	--421
		x"41",	--422
		x"4b",	--423
		x"53",	--424
		x"41",	--425
		x"53",	--426
		x"12",	--427
		x"e3",	--428
		x"93",	--429
		x"00",	--430
		x"24",	--431
		x"41",	--432
		x"00",	--433
		x"12",	--434
		x"12",	--435
		x"12",	--436
		x"f8",	--437
		x"12",	--438
		x"e8",	--439
		x"50",	--440
		x"00",	--441
		x"43",	--442
		x"52",	--443
		x"41",	--444
		x"41",	--445
		x"12",	--446
		x"f8",	--447
		x"12",	--448
		x"e8",	--449
		x"4b",	--450
		x"11",	--451
		x"4f",	--452
		x"00",	--453
		x"12",	--454
		x"f8",	--455
		x"12",	--456
		x"e8",	--457
		x"52",	--458
		x"43",	--459
		x"52",	--460
		x"41",	--461
		x"41",	--462
		x"12",	--463
		x"f8",	--464
		x"12",	--465
		x"e8",	--466
		x"53",	--467
		x"43",	--468
		x"3f",	--469
		x"12",	--470
		x"12",	--471
		x"12",	--472
		x"12",	--473
		x"12",	--474
		x"43",	--475
		x"00",	--476
		x"43",	--477
		x"00",	--478
		x"4e",	--479
		x"93",	--480
		x"24",	--481
		x"4e",	--482
		x"53",	--483
		x"4e",	--484
		x"43",	--485
		x"43",	--486
		x"43",	--487
		x"3c",	--488
		x"90",	--489
		x"00",	--490
		x"2c",	--491
		x"4f",	--492
		x"5c",	--493
		x"5c",	--494
		x"5c",	--495
		x"5c",	--496
		x"4c",	--497
		x"00",	--498
		x"50",	--499
		x"ff",	--500
		x"48",	--501
		x"11",	--502
		x"5a",	--503
		x"4c",	--504
		x"00",	--505
		x"43",	--506
		x"53",	--507
		x"49",	--508
		x"4b",	--509
		x"4b",	--510
		x"93",	--511
		x"24",	--512
		x"90",	--513
		x"00",	--514
		x"24",	--515
		x"90",	--516
		x"00",	--517
		x"24",	--518
		x"4c",	--519
		x"50",	--520
		x"ff",	--521
		x"93",	--522
		x"23",	--523
		x"90",	--524
		x"00",	--525
		x"2c",	--526
		x"4f",	--527
		x"5a",	--528
		x"4a",	--529
		x"5c",	--530
		x"5c",	--531
		x"5a",	--532
		x"4c",	--533
		x"00",	--534
		x"50",	--535
		x"ff",	--536
		x"48",	--537
		x"11",	--538
		x"58",	--539
		x"4c",	--540
		x"00",	--541
		x"3f",	--542
		x"43",	--543
		x"3f",	--544
		x"4c",	--545
		x"50",	--546
		x"ff",	--547
		x"90",	--548
		x"00",	--549
		x"2c",	--550
		x"4f",	--551
		x"5c",	--552
		x"5c",	--553
		x"5c",	--554
		x"5c",	--555
		x"4c",	--556
		x"00",	--557
		x"50",	--558
		x"ff",	--559
		x"3f",	--560
		x"4c",	--561
		x"50",	--562
		x"ff",	--563
		x"90",	--564
		x"00",	--565
		x"2c",	--566
		x"4f",	--567
		x"5c",	--568
		x"5c",	--569
		x"5c",	--570
		x"5c",	--571
		x"4c",	--572
		x"00",	--573
		x"50",	--574
		x"ff",	--575
		x"3f",	--576
		x"43",	--577
		x"00",	--578
		x"43",	--579
		x"41",	--580
		x"41",	--581
		x"41",	--582
		x"41",	--583
		x"41",	--584
		x"41",	--585
		x"43",	--586
		x"00",	--587
		x"4a",	--588
		x"53",	--589
		x"5e",	--590
		x"41",	--591
		x"41",	--592
		x"41",	--593
		x"41",	--594
		x"41",	--595
		x"41",	--596
		x"11",	--597
		x"12",	--598
		x"12",	--599
		x"f8",	--600
		x"12",	--601
		x"e8",	--602
		x"52",	--603
		x"43",	--604
		x"41",	--605
		x"41",	--606
		x"41",	--607
		x"41",	--608
		x"41",	--609
		x"41",	--610
		x"12",	--611
		x"12",	--612
		x"4e",	--613
		x"4c",	--614
		x"4e",	--615
		x"00",	--616
		x"4d",	--617
		x"00",	--618
		x"4c",	--619
		x"00",	--620
		x"4d",	--621
		x"43",	--622
		x"40",	--623
		x"36",	--624
		x"40",	--625
		x"01",	--626
		x"12",	--627
		x"f6",	--628
		x"4e",	--629
		x"00",	--630
		x"12",	--631
		x"c2",	--632
		x"43",	--633
		x"4a",	--634
		x"01",	--635
		x"40",	--636
		x"00",	--637
		x"01",	--638
		x"42",	--639
		x"01",	--640
		x"00",	--641
		x"41",	--642
		x"43",	--643
		x"41",	--644
		x"41",	--645
		x"41",	--646
		x"12",	--647
		x"12",	--648
		x"12",	--649
		x"43",	--650
		x"00",	--651
		x"40",	--652
		x"3f",	--653
		x"00",	--654
		x"4f",	--655
		x"4b",	--656
		x"00",	--657
		x"43",	--658
		x"12",	--659
		x"f1",	--660
		x"43",	--661
		x"40",	--662
		x"3f",	--663
		x"12",	--664
		x"ed",	--665
		x"4e",	--666
		x"4f",	--667
		x"4b",	--668
		x"00",	--669
		x"43",	--670
		x"12",	--671
		x"f1",	--672
		x"4e",	--673
		x"4f",	--674
		x"48",	--675
		x"49",	--676
		x"12",	--677
		x"ec",	--678
		x"12",	--679
		x"e9",	--680
		x"4e",	--681
		x"00",	--682
		x"43",	--683
		x"00",	--684
		x"41",	--685
		x"41",	--686
		x"41",	--687
		x"41",	--688
		x"12",	--689
		x"12",	--690
		x"12",	--691
		x"4d",	--692
		x"4e",	--693
		x"4d",	--694
		x"00",	--695
		x"4e",	--696
		x"00",	--697
		x"4f",	--698
		x"49",	--699
		x"00",	--700
		x"43",	--701
		x"12",	--702
		x"f1",	--703
		x"4e",	--704
		x"4f",	--705
		x"4a",	--706
		x"4b",	--707
		x"12",	--708
		x"ed",	--709
		x"4e",	--710
		x"4f",	--711
		x"49",	--712
		x"00",	--713
		x"43",	--714
		x"12",	--715
		x"f1",	--716
		x"4e",	--717
		x"4f",	--718
		x"4a",	--719
		x"4b",	--720
		x"12",	--721
		x"ec",	--722
		x"12",	--723
		x"e9",	--724
		x"4e",	--725
		x"00",	--726
		x"41",	--727
		x"41",	--728
		x"41",	--729
		x"41",	--730
		x"41",	--731
		x"42",	--732
		x"02",	--733
		x"90",	--734
		x"00",	--735
		x"34",	--736
		x"4c",	--737
		x"5d",	--738
		x"5d",	--739
		x"50",	--740
		x"02",	--741
		x"4f",	--742
		x"00",	--743
		x"4e",	--744
		x"00",	--745
		x"53",	--746
		x"4c",	--747
		x"02",	--748
		x"43",	--749
		x"41",	--750
		x"43",	--751
		x"41",	--752
		x"12",	--753
		x"42",	--754
		x"02",	--755
		x"93",	--756
		x"38",	--757
		x"92",	--758
		x"02",	--759
		x"24",	--760
		x"40",	--761
		x"02",	--762
		x"43",	--763
		x"3c",	--764
		x"52",	--765
		x"9f",	--766
		x"ff",	--767
		x"24",	--768
		x"53",	--769
		x"9b",	--770
		x"23",	--771
		x"12",	--772
		x"f8",	--773
		x"12",	--774
		x"e8",	--775
		x"53",	--776
		x"43",	--777
		x"41",	--778
		x"41",	--779
		x"43",	--780
		x"5c",	--781
		x"5c",	--782
		x"50",	--783
		x"02",	--784
		x"4e",	--785
		x"12",	--786
		x"00",	--787
		x"41",	--788
		x"41",	--789
		x"42",	--790
		x"00",	--791
		x"f2",	--792
		x"23",	--793
		x"4f",	--794
		x"00",	--795
		x"43",	--796
		x"41",	--797
		x"f0",	--798
		x"00",	--799
		x"4f",	--800
		x"f9",	--801
		x"11",	--802
		x"12",	--803
		x"e6",	--804
		x"41",	--805
		x"12",	--806
		x"4f",	--807
		x"4f",	--808
		x"11",	--809
		x"11",	--810
		x"11",	--811
		x"11",	--812
		x"4e",	--813
		x"12",	--814
		x"e6",	--815
		x"4b",	--816
		x"12",	--817
		x"e6",	--818
		x"41",	--819
		x"41",	--820
		x"12",	--821
		x"12",	--822
		x"4f",	--823
		x"40",	--824
		x"00",	--825
		x"4a",	--826
		x"4b",	--827
		x"f0",	--828
		x"00",	--829
		x"24",	--830
		x"11",	--831
		x"53",	--832
		x"23",	--833
		x"f3",	--834
		x"24",	--835
		x"40",	--836
		x"00",	--837
		x"12",	--838
		x"e6",	--839
		x"53",	--840
		x"93",	--841
		x"23",	--842
		x"41",	--843
		x"41",	--844
		x"41",	--845
		x"40",	--846
		x"00",	--847
		x"3f",	--848
		x"12",	--849
		x"4f",	--850
		x"4f",	--851
		x"10",	--852
		x"11",	--853
		x"4e",	--854
		x"12",	--855
		x"e6",	--856
		x"4b",	--857
		x"12",	--858
		x"e6",	--859
		x"41",	--860
		x"41",	--861
		x"12",	--862
		x"12",	--863
		x"4e",	--864
		x"4f",	--865
		x"4f",	--866
		x"10",	--867
		x"11",	--868
		x"4d",	--869
		x"12",	--870
		x"e6",	--871
		x"4b",	--872
		x"12",	--873
		x"e6",	--874
		x"4b",	--875
		x"4a",	--876
		x"10",	--877
		x"10",	--878
		x"ec",	--879
		x"ec",	--880
		x"4d",	--881
		x"12",	--882
		x"e6",	--883
		x"4a",	--884
		x"12",	--885
		x"e6",	--886
		x"41",	--887
		x"41",	--888
		x"41",	--889
		x"12",	--890
		x"12",	--891
		x"12",	--892
		x"4f",	--893
		x"93",	--894
		x"24",	--895
		x"4e",	--896
		x"53",	--897
		x"43",	--898
		x"4a",	--899
		x"5b",	--900
		x"4d",	--901
		x"11",	--902
		x"12",	--903
		x"e6",	--904
		x"99",	--905
		x"24",	--906
		x"53",	--907
		x"b0",	--908
		x"00",	--909
		x"20",	--910
		x"40",	--911
		x"00",	--912
		x"12",	--913
		x"e6",	--914
		x"3f",	--915
		x"40",	--916
		x"00",	--917
		x"12",	--918
		x"e6",	--919
		x"3f",	--920
		x"41",	--921
		x"41",	--922
		x"41",	--923
		x"41",	--924
		x"12",	--925
		x"12",	--926
		x"12",	--927
		x"4f",	--928
		x"93",	--929
		x"24",	--930
		x"4e",	--931
		x"53",	--932
		x"43",	--933
		x"4a",	--934
		x"11",	--935
		x"12",	--936
		x"e6",	--937
		x"99",	--938
		x"24",	--939
		x"53",	--940
		x"b0",	--941
		x"00",	--942
		x"23",	--943
		x"40",	--944
		x"00",	--945
		x"12",	--946
		x"e6",	--947
		x"4a",	--948
		x"11",	--949
		x"12",	--950
		x"e6",	--951
		x"99",	--952
		x"23",	--953
		x"41",	--954
		x"41",	--955
		x"41",	--956
		x"41",	--957
		x"12",	--958
		x"12",	--959
		x"12",	--960
		x"50",	--961
		x"ff",	--962
		x"4f",	--963
		x"93",	--964
		x"38",	--965
		x"90",	--966
		x"00",	--967
		x"38",	--968
		x"43",	--969
		x"41",	--970
		x"59",	--971
		x"40",	--972
		x"00",	--973
		x"4b",	--974
		x"12",	--975
		x"f6",	--976
		x"50",	--977
		x"00",	--978
		x"4f",	--979
		x"00",	--980
		x"53",	--981
		x"40",	--982
		x"00",	--983
		x"4b",	--984
		x"12",	--985
		x"f6",	--986
		x"4f",	--987
		x"90",	--988
		x"00",	--989
		x"37",	--990
		x"49",	--991
		x"53",	--992
		x"51",	--993
		x"40",	--994
		x"00",	--995
		x"4b",	--996
		x"12",	--997
		x"f6",	--998
		x"50",	--999
		x"00",	--1000
		x"4f",	--1001
		x"00",	--1002
		x"53",	--1003
		x"41",	--1004
		x"5a",	--1005
		x"4f",	--1006
		x"11",	--1007
		x"12",	--1008
		x"e6",	--1009
		x"93",	--1010
		x"23",	--1011
		x"50",	--1012
		x"00",	--1013
		x"41",	--1014
		x"41",	--1015
		x"41",	--1016
		x"41",	--1017
		x"40",	--1018
		x"00",	--1019
		x"12",	--1020
		x"e6",	--1021
		x"e3",	--1022
		x"53",	--1023
		x"3f",	--1024
		x"43",	--1025
		x"43",	--1026
		x"3f",	--1027
		x"12",	--1028
		x"12",	--1029
		x"12",	--1030
		x"41",	--1031
		x"52",	--1032
		x"4b",	--1033
		x"49",	--1034
		x"93",	--1035
		x"20",	--1036
		x"3c",	--1037
		x"11",	--1038
		x"12",	--1039
		x"e6",	--1040
		x"49",	--1041
		x"4a",	--1042
		x"53",	--1043
		x"4a",	--1044
		x"00",	--1045
		x"93",	--1046
		x"24",	--1047
		x"90",	--1048
		x"00",	--1049
		x"23",	--1050
		x"49",	--1051
		x"53",	--1052
		x"49",	--1053
		x"00",	--1054
		x"50",	--1055
		x"ff",	--1056
		x"90",	--1057
		x"00",	--1058
		x"2f",	--1059
		x"4f",	--1060
		x"5f",	--1061
		x"4f",	--1062
		x"f8",	--1063
		x"41",	--1064
		x"41",	--1065
		x"41",	--1066
		x"41",	--1067
		x"4b",	--1068
		x"52",	--1069
		x"4b",	--1070
		x"00",	--1071
		x"4b",	--1072
		x"12",	--1073
		x"e6",	--1074
		x"49",	--1075
		x"3f",	--1076
		x"4b",	--1077
		x"53",	--1078
		x"4b",	--1079
		x"12",	--1080
		x"e6",	--1081
		x"49",	--1082
		x"3f",	--1083
		x"4b",	--1084
		x"53",	--1085
		x"4f",	--1086
		x"49",	--1087
		x"93",	--1088
		x"27",	--1089
		x"53",	--1090
		x"11",	--1091
		x"12",	--1092
		x"e6",	--1093
		x"49",	--1094
		x"93",	--1095
		x"23",	--1096
		x"3f",	--1097
		x"4b",	--1098
		x"52",	--1099
		x"4b",	--1100
		x"00",	--1101
		x"4b",	--1102
		x"12",	--1103
		x"e7",	--1104
		x"49",	--1105
		x"3f",	--1106
		x"4b",	--1107
		x"53",	--1108
		x"4b",	--1109
		x"4e",	--1110
		x"10",	--1111
		x"11",	--1112
		x"10",	--1113
		x"11",	--1114
		x"12",	--1115
		x"e6",	--1116
		x"49",	--1117
		x"3f",	--1118
		x"4b",	--1119
		x"53",	--1120
		x"4b",	--1121
		x"12",	--1122
		x"e7",	--1123
		x"49",	--1124
		x"3f",	--1125
		x"4b",	--1126
		x"53",	--1127
		x"4b",	--1128
		x"12",	--1129
		x"e6",	--1130
		x"49",	--1131
		x"3f",	--1132
		x"4b",	--1133
		x"53",	--1134
		x"4b",	--1135
		x"12",	--1136
		x"e6",	--1137
		x"49",	--1138
		x"3f",	--1139
		x"4b",	--1140
		x"53",	--1141
		x"4b",	--1142
		x"12",	--1143
		x"e6",	--1144
		x"49",	--1145
		x"3f",	--1146
		x"40",	--1147
		x"00",	--1148
		x"12",	--1149
		x"e6",	--1150
		x"3f",	--1151
		x"12",	--1152
		x"12",	--1153
		x"42",	--1154
		x"02",	--1155
		x"42",	--1156
		x"00",	--1157
		x"03",	--1158
		x"42",	--1159
		x"02",	--1160
		x"90",	--1161
		x"00",	--1162
		x"34",	--1163
		x"53",	--1164
		x"02",	--1165
		x"42",	--1166
		x"02",	--1167
		x"42",	--1168
		x"02",	--1169
		x"9f",	--1170
		x"20",	--1171
		x"53",	--1172
		x"02",	--1173
		x"40",	--1174
		x"00",	--1175
		x"00",	--1176
		x"c0",	--1177
		x"00",	--1178
		x"00",	--1179
		x"41",	--1180
		x"41",	--1181
		x"c0",	--1182
		x"00",	--1183
		x"00",	--1184
		x"13",	--1185
		x"43",	--1186
		x"02",	--1187
		x"3f",	--1188
		x"40",	--1189
		x"09",	--1190
		x"00",	--1191
		x"40",	--1192
		x"00",	--1193
		x"00",	--1194
		x"41",	--1195
		x"42",	--1196
		x"02",	--1197
		x"42",	--1198
		x"02",	--1199
		x"9f",	--1200
		x"38",	--1201
		x"42",	--1202
		x"02",	--1203
		x"82",	--1204
		x"02",	--1205
		x"41",	--1206
		x"42",	--1207
		x"02",	--1208
		x"42",	--1209
		x"02",	--1210
		x"40",	--1211
		x"00",	--1212
		x"8d",	--1213
		x"8e",	--1214
		x"41",	--1215
		x"42",	--1216
		x"02",	--1217
		x"4f",	--1218
		x"03",	--1219
		x"42",	--1220
		x"02",	--1221
		x"42",	--1222
		x"02",	--1223
		x"9e",	--1224
		x"24",	--1225
		x"42",	--1226
		x"02",	--1227
		x"90",	--1228
		x"00",	--1229
		x"38",	--1230
		x"43",	--1231
		x"02",	--1232
		x"41",	--1233
		x"53",	--1234
		x"02",	--1235
		x"41",	--1236
		x"43",	--1237
		x"41",	--1238
		x"12",	--1239
		x"12",	--1240
		x"4e",	--1241
		x"4f",	--1242
		x"43",	--1243
		x"40",	--1244
		x"4f",	--1245
		x"12",	--1246
		x"f0",	--1247
		x"93",	--1248
		x"34",	--1249
		x"4a",	--1250
		x"4b",	--1251
		x"12",	--1252
		x"f0",	--1253
		x"41",	--1254
		x"41",	--1255
		x"41",	--1256
		x"43",	--1257
		x"40",	--1258
		x"4f",	--1259
		x"4a",	--1260
		x"4b",	--1261
		x"12",	--1262
		x"ec",	--1263
		x"12",	--1264
		x"f0",	--1265
		x"53",	--1266
		x"60",	--1267
		x"80",	--1268
		x"41",	--1269
		x"41",	--1270
		x"41",	--1271
		x"12",	--1272
		x"12",	--1273
		x"12",	--1274
		x"12",	--1275
		x"12",	--1276
		x"12",	--1277
		x"12",	--1278
		x"12",	--1279
		x"50",	--1280
		x"ff",	--1281
		x"4d",	--1282
		x"4f",	--1283
		x"93",	--1284
		x"28",	--1285
		x"4e",	--1286
		x"93",	--1287
		x"28",	--1288
		x"92",	--1289
		x"20",	--1290
		x"40",	--1291
		x"ec",	--1292
		x"92",	--1293
		x"24",	--1294
		x"93",	--1295
		x"24",	--1296
		x"93",	--1297
		x"24",	--1298
		x"4f",	--1299
		x"00",	--1300
		x"00",	--1301
		x"4e",	--1302
		x"00",	--1303
		x"4f",	--1304
		x"00",	--1305
		x"4f",	--1306
		x"00",	--1307
		x"4e",	--1308
		x"00",	--1309
		x"4e",	--1310
		x"00",	--1311
		x"41",	--1312
		x"8b",	--1313
		x"4c",	--1314
		x"93",	--1315
		x"38",	--1316
		x"90",	--1317
		x"00",	--1318
		x"34",	--1319
		x"93",	--1320
		x"38",	--1321
		x"46",	--1322
		x"00",	--1323
		x"47",	--1324
		x"00",	--1325
		x"49",	--1326
		x"f0",	--1327
		x"00",	--1328
		x"24",	--1329
		x"46",	--1330
		x"47",	--1331
		x"c3",	--1332
		x"10",	--1333
		x"10",	--1334
		x"53",	--1335
		x"23",	--1336
		x"4a",	--1337
		x"00",	--1338
		x"4b",	--1339
		x"00",	--1340
		x"43",	--1341
		x"43",	--1342
		x"f0",	--1343
		x"00",	--1344
		x"24",	--1345
		x"5c",	--1346
		x"6d",	--1347
		x"53",	--1348
		x"23",	--1349
		x"53",	--1350
		x"63",	--1351
		x"f6",	--1352
		x"f7",	--1353
		x"43",	--1354
		x"43",	--1355
		x"93",	--1356
		x"20",	--1357
		x"93",	--1358
		x"24",	--1359
		x"41",	--1360
		x"00",	--1361
		x"41",	--1362
		x"00",	--1363
		x"da",	--1364
		x"db",	--1365
		x"4f",	--1366
		x"00",	--1367
		x"9e",	--1368
		x"00",	--1369
		x"20",	--1370
		x"4f",	--1371
		x"00",	--1372
		x"41",	--1373
		x"00",	--1374
		x"46",	--1375
		x"47",	--1376
		x"54",	--1377
		x"65",	--1378
		x"4e",	--1379
		x"00",	--1380
		x"4f",	--1381
		x"00",	--1382
		x"40",	--1383
		x"00",	--1384
		x"00",	--1385
		x"93",	--1386
		x"38",	--1387
		x"48",	--1388
		x"50",	--1389
		x"00",	--1390
		x"41",	--1391
		x"41",	--1392
		x"41",	--1393
		x"41",	--1394
		x"41",	--1395
		x"41",	--1396
		x"41",	--1397
		x"41",	--1398
		x"41",	--1399
		x"91",	--1400
		x"38",	--1401
		x"4b",	--1402
		x"00",	--1403
		x"43",	--1404
		x"43",	--1405
		x"4f",	--1406
		x"00",	--1407
		x"9e",	--1408
		x"00",	--1409
		x"27",	--1410
		x"93",	--1411
		x"24",	--1412
		x"46",	--1413
		x"47",	--1414
		x"84",	--1415
		x"75",	--1416
		x"93",	--1417
		x"38",	--1418
		x"43",	--1419
		x"00",	--1420
		x"41",	--1421
		x"00",	--1422
		x"4e",	--1423
		x"00",	--1424
		x"4f",	--1425
		x"00",	--1426
		x"4e",	--1427
		x"4f",	--1428
		x"53",	--1429
		x"63",	--1430
		x"90",	--1431
		x"3f",	--1432
		x"28",	--1433
		x"90",	--1434
		x"40",	--1435
		x"2c",	--1436
		x"93",	--1437
		x"2c",	--1438
		x"48",	--1439
		x"00",	--1440
		x"53",	--1441
		x"5e",	--1442
		x"6f",	--1443
		x"4b",	--1444
		x"53",	--1445
		x"4e",	--1446
		x"4f",	--1447
		x"53",	--1448
		x"63",	--1449
		x"90",	--1450
		x"3f",	--1451
		x"2b",	--1452
		x"24",	--1453
		x"4e",	--1454
		x"00",	--1455
		x"4f",	--1456
		x"00",	--1457
		x"4a",	--1458
		x"00",	--1459
		x"40",	--1460
		x"00",	--1461
		x"00",	--1462
		x"93",	--1463
		x"37",	--1464
		x"4e",	--1465
		x"4f",	--1466
		x"f3",	--1467
		x"f3",	--1468
		x"c3",	--1469
		x"10",	--1470
		x"10",	--1471
		x"4c",	--1472
		x"4d",	--1473
		x"de",	--1474
		x"df",	--1475
		x"4a",	--1476
		x"00",	--1477
		x"4b",	--1478
		x"00",	--1479
		x"53",	--1480
		x"00",	--1481
		x"48",	--1482
		x"3f",	--1483
		x"93",	--1484
		x"23",	--1485
		x"4f",	--1486
		x"00",	--1487
		x"4f",	--1488
		x"00",	--1489
		x"00",	--1490
		x"4f",	--1491
		x"00",	--1492
		x"00",	--1493
		x"4f",	--1494
		x"00",	--1495
		x"00",	--1496
		x"4e",	--1497
		x"00",	--1498
		x"ff",	--1499
		x"00",	--1500
		x"4e",	--1501
		x"00",	--1502
		x"4d",	--1503
		x"3f",	--1504
		x"43",	--1505
		x"43",	--1506
		x"3f",	--1507
		x"e3",	--1508
		x"53",	--1509
		x"90",	--1510
		x"00",	--1511
		x"37",	--1512
		x"3f",	--1513
		x"93",	--1514
		x"2b",	--1515
		x"3f",	--1516
		x"44",	--1517
		x"45",	--1518
		x"86",	--1519
		x"77",	--1520
		x"3f",	--1521
		x"4e",	--1522
		x"3f",	--1523
		x"43",	--1524
		x"00",	--1525
		x"41",	--1526
		x"00",	--1527
		x"e3",	--1528
		x"e3",	--1529
		x"53",	--1530
		x"63",	--1531
		x"4e",	--1532
		x"00",	--1533
		x"4f",	--1534
		x"00",	--1535
		x"3f",	--1536
		x"93",	--1537
		x"27",	--1538
		x"59",	--1539
		x"00",	--1540
		x"44",	--1541
		x"00",	--1542
		x"45",	--1543
		x"00",	--1544
		x"49",	--1545
		x"f0",	--1546
		x"00",	--1547
		x"24",	--1548
		x"4d",	--1549
		x"44",	--1550
		x"45",	--1551
		x"c3",	--1552
		x"10",	--1553
		x"10",	--1554
		x"53",	--1555
		x"23",	--1556
		x"4c",	--1557
		x"00",	--1558
		x"4d",	--1559
		x"00",	--1560
		x"43",	--1561
		x"43",	--1562
		x"f0",	--1563
		x"00",	--1564
		x"24",	--1565
		x"5c",	--1566
		x"6d",	--1567
		x"53",	--1568
		x"23",	--1569
		x"53",	--1570
		x"63",	--1571
		x"f4",	--1572
		x"f5",	--1573
		x"43",	--1574
		x"43",	--1575
		x"93",	--1576
		x"20",	--1577
		x"93",	--1578
		x"20",	--1579
		x"43",	--1580
		x"43",	--1581
		x"41",	--1582
		x"00",	--1583
		x"41",	--1584
		x"00",	--1585
		x"da",	--1586
		x"db",	--1587
		x"3f",	--1588
		x"43",	--1589
		x"43",	--1590
		x"3f",	--1591
		x"92",	--1592
		x"23",	--1593
		x"9e",	--1594
		x"00",	--1595
		x"00",	--1596
		x"27",	--1597
		x"40",	--1598
		x"f9",	--1599
		x"3f",	--1600
		x"50",	--1601
		x"ff",	--1602
		x"4e",	--1603
		x"00",	--1604
		x"4f",	--1605
		x"00",	--1606
		x"4c",	--1607
		x"00",	--1608
		x"4d",	--1609
		x"00",	--1610
		x"41",	--1611
		x"50",	--1612
		x"00",	--1613
		x"41",	--1614
		x"52",	--1615
		x"12",	--1616
		x"f4",	--1617
		x"41",	--1618
		x"50",	--1619
		x"00",	--1620
		x"41",	--1621
		x"12",	--1622
		x"f4",	--1623
		x"41",	--1624
		x"52",	--1625
		x"41",	--1626
		x"50",	--1627
		x"00",	--1628
		x"41",	--1629
		x"50",	--1630
		x"00",	--1631
		x"12",	--1632
		x"e9",	--1633
		x"12",	--1634
		x"f2",	--1635
		x"50",	--1636
		x"00",	--1637
		x"41",	--1638
		x"50",	--1639
		x"ff",	--1640
		x"4e",	--1641
		x"00",	--1642
		x"4f",	--1643
		x"00",	--1644
		x"4c",	--1645
		x"00",	--1646
		x"4d",	--1647
		x"00",	--1648
		x"41",	--1649
		x"50",	--1650
		x"00",	--1651
		x"41",	--1652
		x"52",	--1653
		x"12",	--1654
		x"f4",	--1655
		x"41",	--1656
		x"50",	--1657
		x"00",	--1658
		x"41",	--1659
		x"12",	--1660
		x"f4",	--1661
		x"e3",	--1662
		x"00",	--1663
		x"41",	--1664
		x"52",	--1665
		x"41",	--1666
		x"50",	--1667
		x"00",	--1668
		x"41",	--1669
		x"50",	--1670
		x"00",	--1671
		x"12",	--1672
		x"e9",	--1673
		x"12",	--1674
		x"f2",	--1675
		x"50",	--1676
		x"00",	--1677
		x"41",	--1678
		x"12",	--1679
		x"12",	--1680
		x"12",	--1681
		x"12",	--1682
		x"12",	--1683
		x"12",	--1684
		x"12",	--1685
		x"12",	--1686
		x"50",	--1687
		x"ff",	--1688
		x"4e",	--1689
		x"00",	--1690
		x"4f",	--1691
		x"00",	--1692
		x"4c",	--1693
		x"00",	--1694
		x"4d",	--1695
		x"00",	--1696
		x"41",	--1697
		x"50",	--1698
		x"00",	--1699
		x"41",	--1700
		x"52",	--1701
		x"12",	--1702
		x"f4",	--1703
		x"41",	--1704
		x"50",	--1705
		x"00",	--1706
		x"41",	--1707
		x"12",	--1708
		x"f4",	--1709
		x"41",	--1710
		x"00",	--1711
		x"93",	--1712
		x"28",	--1713
		x"41",	--1714
		x"00",	--1715
		x"93",	--1716
		x"28",	--1717
		x"92",	--1718
		x"24",	--1719
		x"92",	--1720
		x"24",	--1721
		x"93",	--1722
		x"24",	--1723
		x"93",	--1724
		x"24",	--1725
		x"41",	--1726
		x"00",	--1727
		x"41",	--1728
		x"00",	--1729
		x"41",	--1730
		x"00",	--1731
		x"41",	--1732
		x"00",	--1733
		x"40",	--1734
		x"00",	--1735
		x"43",	--1736
		x"43",	--1737
		x"43",	--1738
		x"43",	--1739
		x"43",	--1740
		x"00",	--1741
		x"43",	--1742
		x"00",	--1743
		x"43",	--1744
		x"43",	--1745
		x"4c",	--1746
		x"00",	--1747
		x"3c",	--1748
		x"58",	--1749
		x"69",	--1750
		x"c3",	--1751
		x"10",	--1752
		x"10",	--1753
		x"53",	--1754
		x"00",	--1755
		x"24",	--1756
		x"b3",	--1757
		x"24",	--1758
		x"58",	--1759
		x"69",	--1760
		x"56",	--1761
		x"67",	--1762
		x"43",	--1763
		x"43",	--1764
		x"99",	--1765
		x"28",	--1766
		x"24",	--1767
		x"43",	--1768
		x"43",	--1769
		x"5c",	--1770
		x"6d",	--1771
		x"56",	--1772
		x"67",	--1773
		x"93",	--1774
		x"37",	--1775
		x"d3",	--1776
		x"d3",	--1777
		x"3f",	--1778
		x"98",	--1779
		x"2b",	--1780
		x"3f",	--1781
		x"4a",	--1782
		x"00",	--1783
		x"4b",	--1784
		x"00",	--1785
		x"4f",	--1786
		x"41",	--1787
		x"00",	--1788
		x"51",	--1789
		x"00",	--1790
		x"4a",	--1791
		x"53",	--1792
		x"46",	--1793
		x"00",	--1794
		x"43",	--1795
		x"91",	--1796
		x"00",	--1797
		x"00",	--1798
		x"24",	--1799
		x"4d",	--1800
		x"00",	--1801
		x"93",	--1802
		x"38",	--1803
		x"90",	--1804
		x"40",	--1805
		x"2c",	--1806
		x"41",	--1807
		x"00",	--1808
		x"53",	--1809
		x"41",	--1810
		x"00",	--1811
		x"41",	--1812
		x"00",	--1813
		x"4d",	--1814
		x"5e",	--1815
		x"6f",	--1816
		x"93",	--1817
		x"38",	--1818
		x"5a",	--1819
		x"6b",	--1820
		x"53",	--1821
		x"90",	--1822
		x"40",	--1823
		x"2b",	--1824
		x"4a",	--1825
		x"00",	--1826
		x"4b",	--1827
		x"00",	--1828
		x"4c",	--1829
		x"00",	--1830
		x"4e",	--1831
		x"4f",	--1832
		x"f0",	--1833
		x"00",	--1834
		x"f3",	--1835
		x"90",	--1836
		x"00",	--1837
		x"24",	--1838
		x"4e",	--1839
		x"00",	--1840
		x"4f",	--1841
		x"00",	--1842
		x"40",	--1843
		x"00",	--1844
		x"00",	--1845
		x"41",	--1846
		x"52",	--1847
		x"12",	--1848
		x"f2",	--1849
		x"50",	--1850
		x"00",	--1851
		x"41",	--1852
		x"41",	--1853
		x"41",	--1854
		x"41",	--1855
		x"41",	--1856
		x"41",	--1857
		x"41",	--1858
		x"41",	--1859
		x"41",	--1860
		x"d3",	--1861
		x"d3",	--1862
		x"3f",	--1863
		x"50",	--1864
		x"00",	--1865
		x"4a",	--1866
		x"b3",	--1867
		x"24",	--1868
		x"41",	--1869
		x"00",	--1870
		x"41",	--1871
		x"00",	--1872
		x"c3",	--1873
		x"10",	--1874
		x"10",	--1875
		x"4c",	--1876
		x"4d",	--1877
		x"d3",	--1878
		x"d0",	--1879
		x"80",	--1880
		x"46",	--1881
		x"00",	--1882
		x"47",	--1883
		x"00",	--1884
		x"c3",	--1885
		x"10",	--1886
		x"10",	--1887
		x"53",	--1888
		x"93",	--1889
		x"3b",	--1890
		x"48",	--1891
		x"00",	--1892
		x"3f",	--1893
		x"93",	--1894
		x"24",	--1895
		x"43",	--1896
		x"91",	--1897
		x"00",	--1898
		x"00",	--1899
		x"24",	--1900
		x"4f",	--1901
		x"00",	--1902
		x"41",	--1903
		x"50",	--1904
		x"00",	--1905
		x"3f",	--1906
		x"93",	--1907
		x"23",	--1908
		x"4e",	--1909
		x"4f",	--1910
		x"f0",	--1911
		x"00",	--1912
		x"f3",	--1913
		x"93",	--1914
		x"23",	--1915
		x"93",	--1916
		x"23",	--1917
		x"93",	--1918
		x"00",	--1919
		x"20",	--1920
		x"93",	--1921
		x"00",	--1922
		x"27",	--1923
		x"50",	--1924
		x"00",	--1925
		x"63",	--1926
		x"f0",	--1927
		x"ff",	--1928
		x"f3",	--1929
		x"3f",	--1930
		x"43",	--1931
		x"3f",	--1932
		x"43",	--1933
		x"3f",	--1934
		x"43",	--1935
		x"91",	--1936
		x"00",	--1937
		x"00",	--1938
		x"24",	--1939
		x"4f",	--1940
		x"00",	--1941
		x"41",	--1942
		x"50",	--1943
		x"00",	--1944
		x"3f",	--1945
		x"43",	--1946
		x"3f",	--1947
		x"93",	--1948
		x"23",	--1949
		x"40",	--1950
		x"f9",	--1951
		x"3f",	--1952
		x"12",	--1953
		x"12",	--1954
		x"12",	--1955
		x"12",	--1956
		x"12",	--1957
		x"50",	--1958
		x"ff",	--1959
		x"4e",	--1960
		x"00",	--1961
		x"4f",	--1962
		x"00",	--1963
		x"4c",	--1964
		x"00",	--1965
		x"4d",	--1966
		x"00",	--1967
		x"41",	--1968
		x"50",	--1969
		x"00",	--1970
		x"41",	--1971
		x"52",	--1972
		x"12",	--1973
		x"f4",	--1974
		x"41",	--1975
		x"52",	--1976
		x"41",	--1977
		x"12",	--1978
		x"f4",	--1979
		x"41",	--1980
		x"00",	--1981
		x"93",	--1982
		x"28",	--1983
		x"41",	--1984
		x"00",	--1985
		x"93",	--1986
		x"28",	--1987
		x"e1",	--1988
		x"00",	--1989
		x"00",	--1990
		x"92",	--1991
		x"24",	--1992
		x"93",	--1993
		x"24",	--1994
		x"92",	--1995
		x"24",	--1996
		x"93",	--1997
		x"24",	--1998
		x"41",	--1999
		x"00",	--2000
		x"81",	--2001
		x"00",	--2002
		x"4d",	--2003
		x"00",	--2004
		x"41",	--2005
		x"00",	--2006
		x"41",	--2007
		x"00",	--2008
		x"41",	--2009
		x"00",	--2010
		x"41",	--2011
		x"00",	--2012
		x"99",	--2013
		x"2c",	--2014
		x"5e",	--2015
		x"6f",	--2016
		x"53",	--2017
		x"4d",	--2018
		x"00",	--2019
		x"40",	--2020
		x"00",	--2021
		x"43",	--2022
		x"40",	--2023
		x"40",	--2024
		x"43",	--2025
		x"43",	--2026
		x"3c",	--2027
		x"dc",	--2028
		x"dd",	--2029
		x"88",	--2030
		x"79",	--2031
		x"c3",	--2032
		x"10",	--2033
		x"10",	--2034
		x"5e",	--2035
		x"6f",	--2036
		x"53",	--2037
		x"24",	--2038
		x"99",	--2039
		x"2b",	--2040
		x"23",	--2041
		x"98",	--2042
		x"2b",	--2043
		x"3f",	--2044
		x"9f",	--2045
		x"2b",	--2046
		x"98",	--2047
		x"2f",	--2048
		x"3f",	--2049
		x"4a",	--2050
		x"4b",	--2051
		x"f0",	--2052
		x"00",	--2053
		x"f3",	--2054
		x"90",	--2055
		x"00",	--2056
		x"24",	--2057
		x"4a",	--2058
		x"00",	--2059
		x"4b",	--2060
		x"00",	--2061
		x"41",	--2062
		x"50",	--2063
		x"00",	--2064
		x"12",	--2065
		x"f2",	--2066
		x"50",	--2067
		x"00",	--2068
		x"41",	--2069
		x"41",	--2070
		x"41",	--2071
		x"41",	--2072
		x"41",	--2073
		x"41",	--2074
		x"42",	--2075
		x"00",	--2076
		x"41",	--2077
		x"50",	--2078
		x"00",	--2079
		x"3f",	--2080
		x"9e",	--2081
		x"23",	--2082
		x"40",	--2083
		x"f9",	--2084
		x"3f",	--2085
		x"93",	--2086
		x"23",	--2087
		x"4a",	--2088
		x"4b",	--2089
		x"f0",	--2090
		x"00",	--2091
		x"f3",	--2092
		x"93",	--2093
		x"23",	--2094
		x"93",	--2095
		x"23",	--2096
		x"93",	--2097
		x"20",	--2098
		x"93",	--2099
		x"27",	--2100
		x"50",	--2101
		x"00",	--2102
		x"63",	--2103
		x"f0",	--2104
		x"ff",	--2105
		x"f3",	--2106
		x"3f",	--2107
		x"43",	--2108
		x"00",	--2109
		x"43",	--2110
		x"00",	--2111
		x"43",	--2112
		x"00",	--2113
		x"41",	--2114
		x"50",	--2115
		x"00",	--2116
		x"3f",	--2117
		x"41",	--2118
		x"52",	--2119
		x"3f",	--2120
		x"50",	--2121
		x"ff",	--2122
		x"4e",	--2123
		x"00",	--2124
		x"4f",	--2125
		x"00",	--2126
		x"4c",	--2127
		x"00",	--2128
		x"4d",	--2129
		x"00",	--2130
		x"41",	--2131
		x"50",	--2132
		x"00",	--2133
		x"41",	--2134
		x"52",	--2135
		x"12",	--2136
		x"f4",	--2137
		x"41",	--2138
		x"52",	--2139
		x"41",	--2140
		x"12",	--2141
		x"f4",	--2142
		x"93",	--2143
		x"00",	--2144
		x"28",	--2145
		x"93",	--2146
		x"00",	--2147
		x"28",	--2148
		x"41",	--2149
		x"52",	--2150
		x"41",	--2151
		x"50",	--2152
		x"00",	--2153
		x"12",	--2154
		x"f5",	--2155
		x"50",	--2156
		x"00",	--2157
		x"41",	--2158
		x"43",	--2159
		x"3f",	--2160
		x"50",	--2161
		x"ff",	--2162
		x"4e",	--2163
		x"00",	--2164
		x"4f",	--2165
		x"00",	--2166
		x"41",	--2167
		x"52",	--2168
		x"41",	--2169
		x"12",	--2170
		x"f4",	--2171
		x"41",	--2172
		x"00",	--2173
		x"93",	--2174
		x"24",	--2175
		x"28",	--2176
		x"92",	--2177
		x"24",	--2178
		x"41",	--2179
		x"00",	--2180
		x"93",	--2181
		x"38",	--2182
		x"90",	--2183
		x"00",	--2184
		x"38",	--2185
		x"93",	--2186
		x"00",	--2187
		x"20",	--2188
		x"43",	--2189
		x"40",	--2190
		x"7f",	--2191
		x"50",	--2192
		x"00",	--2193
		x"41",	--2194
		x"41",	--2195
		x"00",	--2196
		x"41",	--2197
		x"00",	--2198
		x"40",	--2199
		x"00",	--2200
		x"8d",	--2201
		x"4c",	--2202
		x"f0",	--2203
		x"00",	--2204
		x"20",	--2205
		x"93",	--2206
		x"00",	--2207
		x"27",	--2208
		x"e3",	--2209
		x"e3",	--2210
		x"53",	--2211
		x"63",	--2212
		x"50",	--2213
		x"00",	--2214
		x"41",	--2215
		x"43",	--2216
		x"43",	--2217
		x"50",	--2218
		x"00",	--2219
		x"41",	--2220
		x"c3",	--2221
		x"10",	--2222
		x"10",	--2223
		x"53",	--2224
		x"23",	--2225
		x"3f",	--2226
		x"43",	--2227
		x"40",	--2228
		x"80",	--2229
		x"50",	--2230
		x"00",	--2231
		x"41",	--2232
		x"12",	--2233
		x"12",	--2234
		x"12",	--2235
		x"12",	--2236
		x"82",	--2237
		x"4e",	--2238
		x"4f",	--2239
		x"43",	--2240
		x"00",	--2241
		x"93",	--2242
		x"20",	--2243
		x"93",	--2244
		x"20",	--2245
		x"43",	--2246
		x"00",	--2247
		x"41",	--2248
		x"12",	--2249
		x"f2",	--2250
		x"52",	--2251
		x"41",	--2252
		x"41",	--2253
		x"41",	--2254
		x"41",	--2255
		x"41",	--2256
		x"40",	--2257
		x"00",	--2258
		x"00",	--2259
		x"40",	--2260
		x"00",	--2261
		x"00",	--2262
		x"4a",	--2263
		x"00",	--2264
		x"4b",	--2265
		x"00",	--2266
		x"4a",	--2267
		x"4b",	--2268
		x"12",	--2269
		x"f2",	--2270
		x"53",	--2271
		x"93",	--2272
		x"38",	--2273
		x"27",	--2274
		x"4a",	--2275
		x"00",	--2276
		x"4b",	--2277
		x"00",	--2278
		x"4f",	--2279
		x"f0",	--2280
		x"00",	--2281
		x"20",	--2282
		x"40",	--2283
		x"00",	--2284
		x"8f",	--2285
		x"4e",	--2286
		x"00",	--2287
		x"3f",	--2288
		x"51",	--2289
		x"00",	--2290
		x"00",	--2291
		x"61",	--2292
		x"00",	--2293
		x"00",	--2294
		x"53",	--2295
		x"23",	--2296
		x"3f",	--2297
		x"4f",	--2298
		x"e3",	--2299
		x"53",	--2300
		x"43",	--2301
		x"43",	--2302
		x"4e",	--2303
		x"f0",	--2304
		x"00",	--2305
		x"24",	--2306
		x"5c",	--2307
		x"6d",	--2308
		x"53",	--2309
		x"23",	--2310
		x"53",	--2311
		x"63",	--2312
		x"fa",	--2313
		x"fb",	--2314
		x"43",	--2315
		x"43",	--2316
		x"93",	--2317
		x"20",	--2318
		x"93",	--2319
		x"20",	--2320
		x"43",	--2321
		x"43",	--2322
		x"f0",	--2323
		x"00",	--2324
		x"20",	--2325
		x"48",	--2326
		x"49",	--2327
		x"da",	--2328
		x"db",	--2329
		x"4d",	--2330
		x"00",	--2331
		x"4e",	--2332
		x"00",	--2333
		x"40",	--2334
		x"00",	--2335
		x"8f",	--2336
		x"4e",	--2337
		x"00",	--2338
		x"3f",	--2339
		x"c3",	--2340
		x"10",	--2341
		x"10",	--2342
		x"53",	--2343
		x"23",	--2344
		x"3f",	--2345
		x"12",	--2346
		x"12",	--2347
		x"12",	--2348
		x"93",	--2349
		x"2c",	--2350
		x"90",	--2351
		x"01",	--2352
		x"28",	--2353
		x"40",	--2354
		x"00",	--2355
		x"43",	--2356
		x"42",	--2357
		x"4e",	--2358
		x"4f",	--2359
		x"49",	--2360
		x"93",	--2361
		x"20",	--2362
		x"50",	--2363
		x"f9",	--2364
		x"4c",	--2365
		x"43",	--2366
		x"8e",	--2367
		x"7f",	--2368
		x"4a",	--2369
		x"41",	--2370
		x"41",	--2371
		x"41",	--2372
		x"41",	--2373
		x"90",	--2374
		x"01",	--2375
		x"28",	--2376
		x"42",	--2377
		x"43",	--2378
		x"40",	--2379
		x"00",	--2380
		x"4e",	--2381
		x"4f",	--2382
		x"49",	--2383
		x"93",	--2384
		x"27",	--2385
		x"c3",	--2386
		x"10",	--2387
		x"10",	--2388
		x"53",	--2389
		x"23",	--2390
		x"3f",	--2391
		x"40",	--2392
		x"00",	--2393
		x"43",	--2394
		x"40",	--2395
		x"00",	--2396
		x"3f",	--2397
		x"40",	--2398
		x"00",	--2399
		x"43",	--2400
		x"43",	--2401
		x"3f",	--2402
		x"12",	--2403
		x"12",	--2404
		x"12",	--2405
		x"12",	--2406
		x"12",	--2407
		x"4f",	--2408
		x"4f",	--2409
		x"00",	--2410
		x"4f",	--2411
		x"00",	--2412
		x"4d",	--2413
		x"00",	--2414
		x"4d",	--2415
		x"93",	--2416
		x"28",	--2417
		x"92",	--2418
		x"24",	--2419
		x"93",	--2420
		x"24",	--2421
		x"93",	--2422
		x"24",	--2423
		x"4d",	--2424
		x"00",	--2425
		x"90",	--2426
		x"ff",	--2427
		x"38",	--2428
		x"90",	--2429
		x"00",	--2430
		x"34",	--2431
		x"4e",	--2432
		x"4f",	--2433
		x"f0",	--2434
		x"00",	--2435
		x"f3",	--2436
		x"90",	--2437
		x"00",	--2438
		x"24",	--2439
		x"50",	--2440
		x"00",	--2441
		x"63",	--2442
		x"93",	--2443
		x"38",	--2444
		x"4b",	--2445
		x"50",	--2446
		x"00",	--2447
		x"c3",	--2448
		x"10",	--2449
		x"10",	--2450
		x"c3",	--2451
		x"10",	--2452
		x"10",	--2453
		x"c3",	--2454
		x"10",	--2455
		x"10",	--2456
		x"c3",	--2457
		x"10",	--2458
		x"10",	--2459
		x"c3",	--2460
		x"10",	--2461
		x"10",	--2462
		x"c3",	--2463
		x"10",	--2464
		x"10",	--2465
		x"c3",	--2466
		x"10",	--2467
		x"10",	--2468
		x"f3",	--2469
		x"f0",	--2470
		x"00",	--2471
		x"4d",	--2472
		x"3c",	--2473
		x"93",	--2474
		x"23",	--2475
		x"43",	--2476
		x"43",	--2477
		x"43",	--2478
		x"4d",	--2479
		x"5d",	--2480
		x"5d",	--2481
		x"5d",	--2482
		x"5d",	--2483
		x"5d",	--2484
		x"5d",	--2485
		x"5d",	--2486
		x"4f",	--2487
		x"f0",	--2488
		x"00",	--2489
		x"dd",	--2490
		x"4a",	--2491
		x"11",	--2492
		x"43",	--2493
		x"10",	--2494
		x"4c",	--2495
		x"df",	--2496
		x"4d",	--2497
		x"41",	--2498
		x"41",	--2499
		x"41",	--2500
		x"41",	--2501
		x"41",	--2502
		x"41",	--2503
		x"93",	--2504
		x"23",	--2505
		x"4e",	--2506
		x"4f",	--2507
		x"f0",	--2508
		x"00",	--2509
		x"f3",	--2510
		x"93",	--2511
		x"20",	--2512
		x"93",	--2513
		x"27",	--2514
		x"50",	--2515
		x"00",	--2516
		x"63",	--2517
		x"3f",	--2518
		x"c3",	--2519
		x"10",	--2520
		x"10",	--2521
		x"4b",	--2522
		x"50",	--2523
		x"00",	--2524
		x"3f",	--2525
		x"43",	--2526
		x"43",	--2527
		x"43",	--2528
		x"3f",	--2529
		x"d3",	--2530
		x"d0",	--2531
		x"00",	--2532
		x"f3",	--2533
		x"f0",	--2534
		x"00",	--2535
		x"43",	--2536
		x"3f",	--2537
		x"40",	--2538
		x"ff",	--2539
		x"8b",	--2540
		x"90",	--2541
		x"00",	--2542
		x"34",	--2543
		x"4e",	--2544
		x"4f",	--2545
		x"47",	--2546
		x"f0",	--2547
		x"00",	--2548
		x"24",	--2549
		x"c3",	--2550
		x"10",	--2551
		x"10",	--2552
		x"53",	--2553
		x"23",	--2554
		x"43",	--2555
		x"43",	--2556
		x"f0",	--2557
		x"00",	--2558
		x"24",	--2559
		x"58",	--2560
		x"69",	--2561
		x"53",	--2562
		x"23",	--2563
		x"53",	--2564
		x"63",	--2565
		x"fe",	--2566
		x"ff",	--2567
		x"43",	--2568
		x"43",	--2569
		x"93",	--2570
		x"20",	--2571
		x"93",	--2572
		x"20",	--2573
		x"43",	--2574
		x"43",	--2575
		x"4e",	--2576
		x"4f",	--2577
		x"dc",	--2578
		x"dd",	--2579
		x"48",	--2580
		x"49",	--2581
		x"f0",	--2582
		x"00",	--2583
		x"f3",	--2584
		x"90",	--2585
		x"00",	--2586
		x"24",	--2587
		x"50",	--2588
		x"00",	--2589
		x"63",	--2590
		x"48",	--2591
		x"49",	--2592
		x"c3",	--2593
		x"10",	--2594
		x"10",	--2595
		x"c3",	--2596
		x"10",	--2597
		x"10",	--2598
		x"c3",	--2599
		x"10",	--2600
		x"10",	--2601
		x"c3",	--2602
		x"10",	--2603
		x"10",	--2604
		x"c3",	--2605
		x"10",	--2606
		x"10",	--2607
		x"c3",	--2608
		x"10",	--2609
		x"10",	--2610
		x"c3",	--2611
		x"10",	--2612
		x"10",	--2613
		x"f3",	--2614
		x"f0",	--2615
		x"00",	--2616
		x"43",	--2617
		x"90",	--2618
		x"40",	--2619
		x"2f",	--2620
		x"43",	--2621
		x"3f",	--2622
		x"43",	--2623
		x"43",	--2624
		x"3f",	--2625
		x"93",	--2626
		x"23",	--2627
		x"48",	--2628
		x"49",	--2629
		x"f0",	--2630
		x"00",	--2631
		x"f3",	--2632
		x"93",	--2633
		x"24",	--2634
		x"50",	--2635
		x"00",	--2636
		x"63",	--2637
		x"3f",	--2638
		x"93",	--2639
		x"27",	--2640
		x"3f",	--2641
		x"12",	--2642
		x"12",	--2643
		x"4f",	--2644
		x"4f",	--2645
		x"00",	--2646
		x"f0",	--2647
		x"00",	--2648
		x"4f",	--2649
		x"00",	--2650
		x"c3",	--2651
		x"10",	--2652
		x"c3",	--2653
		x"10",	--2654
		x"c3",	--2655
		x"10",	--2656
		x"c3",	--2657
		x"10",	--2658
		x"c3",	--2659
		x"10",	--2660
		x"c3",	--2661
		x"10",	--2662
		x"c3",	--2663
		x"10",	--2664
		x"4d",	--2665
		x"4f",	--2666
		x"00",	--2667
		x"b0",	--2668
		x"00",	--2669
		x"43",	--2670
		x"6f",	--2671
		x"4f",	--2672
		x"00",	--2673
		x"93",	--2674
		x"20",	--2675
		x"93",	--2676
		x"24",	--2677
		x"40",	--2678
		x"ff",	--2679
		x"00",	--2680
		x"4a",	--2681
		x"4b",	--2682
		x"5c",	--2683
		x"6d",	--2684
		x"5c",	--2685
		x"6d",	--2686
		x"5c",	--2687
		x"6d",	--2688
		x"5c",	--2689
		x"6d",	--2690
		x"5c",	--2691
		x"6d",	--2692
		x"5c",	--2693
		x"6d",	--2694
		x"5c",	--2695
		x"6d",	--2696
		x"40",	--2697
		x"00",	--2698
		x"00",	--2699
		x"90",	--2700
		x"40",	--2701
		x"2c",	--2702
		x"40",	--2703
		x"ff",	--2704
		x"5c",	--2705
		x"6d",	--2706
		x"4f",	--2707
		x"53",	--2708
		x"90",	--2709
		x"40",	--2710
		x"2b",	--2711
		x"4a",	--2712
		x"00",	--2713
		x"4c",	--2714
		x"00",	--2715
		x"4d",	--2716
		x"00",	--2717
		x"41",	--2718
		x"41",	--2719
		x"41",	--2720
		x"90",	--2721
		x"00",	--2722
		x"24",	--2723
		x"50",	--2724
		x"ff",	--2725
		x"4d",	--2726
		x"00",	--2727
		x"40",	--2728
		x"00",	--2729
		x"00",	--2730
		x"4a",	--2731
		x"4b",	--2732
		x"5c",	--2733
		x"6d",	--2734
		x"5c",	--2735
		x"6d",	--2736
		x"5c",	--2737
		x"6d",	--2738
		x"5c",	--2739
		x"6d",	--2740
		x"5c",	--2741
		x"6d",	--2742
		x"5c",	--2743
		x"6d",	--2744
		x"5c",	--2745
		x"6d",	--2746
		x"4c",	--2747
		x"4d",	--2748
		x"d3",	--2749
		x"d0",	--2750
		x"40",	--2751
		x"4a",	--2752
		x"00",	--2753
		x"4b",	--2754
		x"00",	--2755
		x"41",	--2756
		x"41",	--2757
		x"41",	--2758
		x"93",	--2759
		x"23",	--2760
		x"43",	--2761
		x"00",	--2762
		x"41",	--2763
		x"41",	--2764
		x"41",	--2765
		x"93",	--2766
		x"24",	--2767
		x"4a",	--2768
		x"4b",	--2769
		x"f3",	--2770
		x"f0",	--2771
		x"00",	--2772
		x"93",	--2773
		x"20",	--2774
		x"93",	--2775
		x"24",	--2776
		x"43",	--2777
		x"00",	--2778
		x"3f",	--2779
		x"93",	--2780
		x"23",	--2781
		x"42",	--2782
		x"00",	--2783
		x"3f",	--2784
		x"43",	--2785
		x"00",	--2786
		x"3f",	--2787
		x"12",	--2788
		x"4f",	--2789
		x"93",	--2790
		x"28",	--2791
		x"4e",	--2792
		x"93",	--2793
		x"28",	--2794
		x"92",	--2795
		x"24",	--2796
		x"92",	--2797
		x"24",	--2798
		x"93",	--2799
		x"24",	--2800
		x"93",	--2801
		x"24",	--2802
		x"4f",	--2803
		x"00",	--2804
		x"9e",	--2805
		x"00",	--2806
		x"24",	--2807
		x"93",	--2808
		x"20",	--2809
		x"43",	--2810
		x"4e",	--2811
		x"41",	--2812
		x"41",	--2813
		x"93",	--2814
		x"24",	--2815
		x"93",	--2816
		x"00",	--2817
		x"23",	--2818
		x"43",	--2819
		x"4e",	--2820
		x"41",	--2821
		x"41",	--2822
		x"93",	--2823
		x"00",	--2824
		x"27",	--2825
		x"43",	--2826
		x"3f",	--2827
		x"4f",	--2828
		x"00",	--2829
		x"4e",	--2830
		x"00",	--2831
		x"9b",	--2832
		x"3b",	--2833
		x"9c",	--2834
		x"38",	--2835
		x"4f",	--2836
		x"00",	--2837
		x"4f",	--2838
		x"00",	--2839
		x"4e",	--2840
		x"00",	--2841
		x"4e",	--2842
		x"00",	--2843
		x"9f",	--2844
		x"2b",	--2845
		x"9e",	--2846
		x"28",	--2847
		x"9b",	--2848
		x"2b",	--2849
		x"9e",	--2850
		x"28",	--2851
		x"9f",	--2852
		x"28",	--2853
		x"9c",	--2854
		x"28",	--2855
		x"43",	--2856
		x"3f",	--2857
		x"93",	--2858
		x"23",	--2859
		x"43",	--2860
		x"3f",	--2861
		x"92",	--2862
		x"23",	--2863
		x"4e",	--2864
		x"00",	--2865
		x"4f",	--2866
		x"00",	--2867
		x"8f",	--2868
		x"3f",	--2869
		x"43",	--2870
		x"93",	--2871
		x"34",	--2872
		x"40",	--2873
		x"00",	--2874
		x"e3",	--2875
		x"53",	--2876
		x"93",	--2877
		x"34",	--2878
		x"e3",	--2879
		x"e3",	--2880
		x"53",	--2881
		x"12",	--2882
		x"12",	--2883
		x"f6",	--2884
		x"41",	--2885
		x"b3",	--2886
		x"24",	--2887
		x"e3",	--2888
		x"53",	--2889
		x"b3",	--2890
		x"24",	--2891
		x"e3",	--2892
		x"53",	--2893
		x"41",	--2894
		x"12",	--2895
		x"f6",	--2896
		x"4e",	--2897
		x"41",	--2898
		x"12",	--2899
		x"43",	--2900
		x"93",	--2901
		x"34",	--2902
		x"40",	--2903
		x"00",	--2904
		x"e3",	--2905
		x"e3",	--2906
		x"53",	--2907
		x"63",	--2908
		x"93",	--2909
		x"34",	--2910
		x"e3",	--2911
		x"e3",	--2912
		x"e3",	--2913
		x"53",	--2914
		x"63",	--2915
		x"12",	--2916
		x"f7",	--2917
		x"b3",	--2918
		x"24",	--2919
		x"e3",	--2920
		x"e3",	--2921
		x"53",	--2922
		x"63",	--2923
		x"b3",	--2924
		x"24",	--2925
		x"e3",	--2926
		x"e3",	--2927
		x"53",	--2928
		x"63",	--2929
		x"41",	--2930
		x"41",	--2931
		x"12",	--2932
		x"f6",	--2933
		x"4c",	--2934
		x"4d",	--2935
		x"41",	--2936
		x"40",	--2937
		x"00",	--2938
		x"4e",	--2939
		x"43",	--2940
		x"5f",	--2941
		x"6e",	--2942
		x"9d",	--2943
		x"28",	--2944
		x"8d",	--2945
		x"d3",	--2946
		x"83",	--2947
		x"23",	--2948
		x"41",	--2949
		x"12",	--2950
		x"f6",	--2951
		x"4e",	--2952
		x"41",	--2953
		x"12",	--2954
		x"12",	--2955
		x"12",	--2956
		x"40",	--2957
		x"00",	--2958
		x"4c",	--2959
		x"4d",	--2960
		x"43",	--2961
		x"43",	--2962
		x"5e",	--2963
		x"6f",	--2964
		x"6c",	--2965
		x"6d",	--2966
		x"9b",	--2967
		x"28",	--2968
		x"20",	--2969
		x"9a",	--2970
		x"28",	--2971
		x"8a",	--2972
		x"7b",	--2973
		x"d3",	--2974
		x"83",	--2975
		x"23",	--2976
		x"41",	--2977
		x"41",	--2978
		x"41",	--2979
		x"41",	--2980
		x"12",	--2981
		x"f7",	--2982
		x"4c",	--2983
		x"4d",	--2984
		x"41",	--2985
		x"13",	--2986
		x"d0",	--2987
		x"00",	--2988
		x"3f",	--2989
		x"61",	--2990
		x"74",	--2991
		x"6e",	--2992
		x"20",	--2993
		x"6f",	--2994
		x"20",	--2995
		x"20",	--2996
		x"65",	--2997
		x"20",	--2998
		x"62",	--2999
		x"6e",	--3000
		x"66",	--3001
		x"6c",	--3002
		x"0d",	--3003
		x"00",	--3004
		x"65",	--3005
		x"73",	--3006
		x"6f",	--3007
		x"6c",	--3008
		x"20",	--3009
		x"6f",	--3010
		x"20",	--3011
		x"65",	--3012
		x"20",	--3013
		x"68",	--3014
		x"74",	--3015
		x"0a",	--3016
		x"63",	--3017
		x"72",	--3018
		x"65",	--3019
		x"74",	--3020
		x"75",	--3021
		x"61",	--3022
		x"65",	--3023
		x"0d",	--3024
		x"00",	--3025
		x"25",	--3026
		x"20",	--3027
		x"45",	--3028
		x"54",	--3029
		x"52",	--3030
		x"47",	--3031
		x"54",	--3032
		x"0a",	--3033
		x"53",	--3034
		x"6d",	--3035
		x"74",	--3036
		x"69",	--3037
		x"67",	--3038
		x"77",	--3039
		x"6e",	--3040
		x"20",	--3041
		x"65",	--3042
		x"72",	--3043
		x"62",	--3044
		x"79",	--3045
		x"77",	--3046
		x"6f",	--3047
		x"67",	--3048
		x"0a",	--3049
		x"0d",	--3050
		x"3d",	--3051
		x"3d",	--3052
		x"3d",	--3053
		x"20",	--3054
		x"61",	--3055
		x"63",	--3056
		x"6c",	--3057
		x"4d",	--3058
		x"55",	--3059
		x"3d",	--3060
		x"3d",	--3061
		x"3d",	--3062
		x"0d",	--3063
		x"00",	--3064
		x"20",	--3065
		x"0d",	--3066
		x"00",	--3067
		x"25",	--3068
		x"0d",	--3069
		x"00",	--3070
		x"20",	--3071
		x"00",	--3072
		x"63",	--3073
		x"77",	--3074
		x"69",	--3075
		x"65",	--3076
		x"0d",	--3077
		x"63",	--3078
		x"72",	--3079
		x"65",	--3080
		x"74",	--3081
		x"75",	--3082
		x"61",	--3083
		x"65",	--3084
		x"0d",	--3085
		x"00",	--3086
		x"25",	--3087
		x"20",	--3088
		x"45",	--3089
		x"49",	--3090
		x"54",	--3091
		x"52",	--3092
		x"56",	--3093
		x"4c",	--3094
		x"45",	--3095
		x"0a",	--3096
		x"53",	--3097
		x"6d",	--3098
		x"74",	--3099
		x"69",	--3100
		x"67",	--3101
		x"77",	--3102
		x"6e",	--3103
		x"20",	--3104
		x"65",	--3105
		x"72",	--3106
		x"62",	--3107
		x"79",	--3108
		x"77",	--3109
		x"6f",	--3110
		x"67",	--3111
		x"0a",	--3112
		x"72",	--3113
		x"25",	--3114
		x"20",	--3115
		x"3d",	--3116
		x"64",	--3117
		x"0a",	--3118
		x"72",	--3119
		x"61",	--3120
		x"0a",	--3121
		x"00",	--3122
		x"25",	--3123
		x"20",	--3124
		x"45",	--3125
		x"49",	--3126
		x"54",	--3127
		x"52",	--3128
		x"0a",	--3129
		x"25",	--3130
		x"20",	--3131
		x"73",	--3132
		x"6e",	--3133
		x"74",	--3134
		x"61",	--3135
		x"6e",	--3136
		x"6d",	--3137
		x"65",	--3138
		x"0d",	--3139
		x"00",	--3140
		x"63",	--3141
		x"20",	--3142
		x"6f",	--3143
		x"73",	--3144
		x"63",	--3145
		x"20",	--3146
		x"6f",	--3147
		x"6d",	--3148
		x"6e",	--3149
		x"0d",	--3150
		x"00",	--3151
		x"e8",	--3152
		x"e8",	--3153
		x"e8",	--3154
		x"e8",	--3155
		x"e8",	--3156
		x"e8",	--3157
		x"e8",	--3158
		x"e8",	--3159
		x"e8",	--3160
		x"e8",	--3161
		x"e8",	--3162
		x"e8",	--3163
		x"e8",	--3164
		x"e8",	--3165
		x"e8",	--3166
		x"e8",	--3167
		x"e8",	--3168
		x"e8",	--3169
		x"e8",	--3170
		x"e8",	--3171
		x"e8",	--3172
		x"e8",	--3173
		x"e8",	--3174
		x"e8",	--3175
		x"e8",	--3176
		x"e8",	--3177
		x"e8",	--3178
		x"e8",	--3179
		x"e8",	--3180
		x"e8",	--3181
		x"e8",	--3182
		x"e8",	--3183
		x"e8",	--3184
		x"e8",	--3185
		x"e8",	--3186
		x"e8",	--3187
		x"e8",	--3188
		x"e8",	--3189
		x"e8",	--3190
		x"e8",	--3191
		x"e8",	--3192
		x"e8",	--3193
		x"e8",	--3194
		x"e8",	--3195
		x"e8",	--3196
		x"e8",	--3197
		x"e8",	--3198
		x"e8",	--3199
		x"e8",	--3200
		x"e8",	--3201
		x"e8",	--3202
		x"e8",	--3203
		x"e8",	--3204
		x"e8",	--3205
		x"e8",	--3206
		x"e8",	--3207
		x"e8",	--3208
		x"e8",	--3209
		x"e8",	--3210
		x"e8",	--3211
		x"e8",	--3212
		x"e8",	--3213
		x"e8",	--3214
		x"e8",	--3215
		x"e8",	--3216
		x"e8",	--3217
		x"e8",	--3218
		x"e8",	--3219
		x"e8",	--3220
		x"e8",	--3221
		x"e8",	--3222
		x"e8",	--3223
		x"e8",	--3224
		x"e8",	--3225
		x"e8",	--3226
		x"e8",	--3227
		x"e8",	--3228
		x"e8",	--3229
		x"e8",	--3230
		x"e8",	--3231
		x"e8",	--3232
		x"e8",	--3233
		x"e8",	--3234
		x"e8",	--3235
		x"31",	--3236
		x"33",	--3237
		x"35",	--3238
		x"37",	--3239
		x"39",	--3240
		x"62",	--3241
		x"64",	--3242
		x"66",	--3243
		x"00",	--3244
		x"00",	--3245
		x"00",	--3246
		x"00",	--3247
		x"00",	--3248
		x"01",	--3249
		x"02",	--3250
		x"03",	--3251
		x"03",	--3252
		x"04",	--3253
		x"04",	--3254
		x"04",	--3255
		x"04",	--3256
		x"05",	--3257
		x"05",	--3258
		x"05",	--3259
		x"05",	--3260
		x"05",	--3261
		x"05",	--3262
		x"05",	--3263
		x"05",	--3264
		x"06",	--3265
		x"06",	--3266
		x"06",	--3267
		x"06",	--3268
		x"06",	--3269
		x"06",	--3270
		x"06",	--3271
		x"06",	--3272
		x"06",	--3273
		x"06",	--3274
		x"06",	--3275
		x"06",	--3276
		x"06",	--3277
		x"06",	--3278
		x"06",	--3279
		x"06",	--3280
		x"07",	--3281
		x"07",	--3282
		x"07",	--3283
		x"07",	--3284
		x"07",	--3285
		x"07",	--3286
		x"07",	--3287
		x"07",	--3288
		x"07",	--3289
		x"07",	--3290
		x"07",	--3291
		x"07",	--3292
		x"07",	--3293
		x"07",	--3294
		x"07",	--3295
		x"07",	--3296
		x"07",	--3297
		x"07",	--3298
		x"07",	--3299
		x"07",	--3300
		x"07",	--3301
		x"07",	--3302
		x"07",	--3303
		x"07",	--3304
		x"07",	--3305
		x"07",	--3306
		x"07",	--3307
		x"07",	--3308
		x"07",	--3309
		x"07",	--3310
		x"07",	--3311
		x"07",	--3312
		x"08",	--3313
		x"08",	--3314
		x"08",	--3315
		x"08",	--3316
		x"08",	--3317
		x"08",	--3318
		x"08",	--3319
		x"08",	--3320
		x"08",	--3321
		x"08",	--3322
		x"08",	--3323
		x"08",	--3324
		x"08",	--3325
		x"08",	--3326
		x"08",	--3327
		x"08",	--3328
		x"08",	--3329
		x"08",	--3330
		x"08",	--3331
		x"08",	--3332
		x"08",	--3333
		x"08",	--3334
		x"08",	--3335
		x"08",	--3336
		x"08",	--3337
		x"08",	--3338
		x"08",	--3339
		x"08",	--3340
		x"08",	--3341
		x"08",	--3342
		x"08",	--3343
		x"08",	--3344
		x"08",	--3345
		x"08",	--3346
		x"08",	--3347
		x"08",	--3348
		x"08",	--3349
		x"08",	--3350
		x"08",	--3351
		x"08",	--3352
		x"08",	--3353
		x"08",	--3354
		x"08",	--3355
		x"08",	--3356
		x"08",	--3357
		x"08",	--3358
		x"08",	--3359
		x"08",	--3360
		x"08",	--3361
		x"08",	--3362
		x"08",	--3363
		x"08",	--3364
		x"08",	--3365
		x"08",	--3366
		x"08",	--3367
		x"08",	--3368
		x"08",	--3369
		x"08",	--3370
		x"08",	--3371
		x"08",	--3372
		x"08",	--3373
		x"08",	--3374
		x"08",	--3375
		x"08",	--3376
		x"ff",	--3377
		x"ff",	--3378
		x"ff",	--3379
		x"ff",	--3380
		x"ff",	--3381
		x"ff",	--3382
		x"ff",	--3383
		x"ff",	--3384
		x"ff",	--3385
		x"ff",	--3386
		x"ff",	--3387
		x"ff",	--3388
		x"ff",	--3389
		x"ff",	--3390
		x"ff",	--3391
		x"ff",	--3392
		x"ff",	--3393
		x"ff",	--3394
		x"ff",	--3395
		x"ff",	--3396
		x"ff",	--3397
		x"ff",	--3398
		x"ff",	--3399
		x"ff",	--3400
		x"ff",	--3401
		x"ff",	--3402
		x"ff",	--3403
		x"ff",	--3404
		x"ff",	--3405
		x"ff",	--3406
		x"ff",	--3407
		x"ff",	--3408
		x"ff",	--3409
		x"ff",	--3410
		x"ff",	--3411
		x"ff",	--3412
		x"ff",	--3413
		x"ff",	--3414
		x"ff",	--3415
		x"ff",	--3416
		x"ff",	--3417
		x"ff",	--3418
		x"ff",	--3419
		x"ff",	--3420
		x"ff",	--3421
		x"ff",	--3422
		x"ff",	--3423
		x"ff",	--3424
		x"ff",	--3425
		x"ff",	--3426
		x"ff",	--3427
		x"ff",	--3428
		x"ff",	--3429
		x"ff",	--3430
		x"ff",	--3431
		x"ff",	--3432
		x"ff",	--3433
		x"ff",	--3434
		x"ff",	--3435
		x"ff",	--3436
		x"ff",	--3437
		x"ff",	--3438
		x"ff",	--3439
		x"ff",	--3440
		x"ff",	--3441
		x"ff",	--3442
		x"ff",	--3443
		x"ff",	--3444
		x"ff",	--3445
		x"ff",	--3446
		x"ff",	--3447
		x"ff",	--3448
		x"ff",	--3449
		x"ff",	--3450
		x"ff",	--3451
		x"ff",	--3452
		x"ff",	--3453
		x"ff",	--3454
		x"ff",	--3455
		x"ff",	--3456
		x"ff",	--3457
		x"ff",	--3458
		x"ff",	--3459
		x"ff",	--3460
		x"ff",	--3461
		x"ff",	--3462
		x"ff",	--3463
		x"ff",	--3464
		x"ff",	--3465
		x"ff",	--3466
		x"ff",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"e9",	--4087
		x"e1",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
