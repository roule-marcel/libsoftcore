library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"24",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"0a",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"24",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"2e",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"1a",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"24",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"0a",	--29
		x"f9",	--30
		x"31",	--31
		x"a6",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"98",	--44
		x"b0",	--45
		x"4a",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"46",	--50
		x"b0",	--51
		x"5c",	--52
		x"21",	--53
		x"3d",	--54
		x"63",	--55
		x"3e",	--56
		x"12",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"7a",	--61
		x"3d",	--62
		x"74",	--63
		x"3e",	--64
		x"82",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"7a",	--69
		x"3d",	--70
		x"7a",	--71
		x"3e",	--72
		x"f6",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"7a",	--77
		x"3d",	--78
		x"7f",	--79
		x"3e",	--80
		x"46",	--81
		x"7f",	--82
		x"70",	--83
		x"b0",	--84
		x"7a",	--85
		x"3d",	--86
		x"83",	--87
		x"3e",	--88
		x"66",	--89
		x"7f",	--90
		x"65",	--91
		x"b0",	--92
		x"7a",	--93
		x"3d",	--94
		x"8b",	--95
		x"3e",	--96
		x"ce",	--97
		x"7f",	--98
		x"73",	--99
		x"b0",	--100
		x"7a",	--101
		x"3d",	--102
		x"9c",	--103
		x"3e",	--104
		x"d2",	--105
		x"7f",	--106
		x"63",	--107
		x"b0",	--108
		x"7a",	--109
		x"3d",	--110
		x"b0",	--111
		x"3e",	--112
		x"d6",	--113
		x"7f",	--114
		x"62",	--115
		x"b0",	--116
		x"7a",	--117
		x"0e",	--118
		x"0f",	--119
		x"b0",	--120
		x"10",	--121
		x"2c",	--122
		x"3d",	--123
		x"20",	--124
		x"3e",	--125
		x"80",	--126
		x"0f",	--127
		x"3f",	--128
		x"0e",	--129
		x"b0",	--130
		x"20",	--131
		x"0f",	--132
		x"3f",	--133
		x"0e",	--134
		x"b0",	--135
		x"68",	--136
		x"2c",	--137
		x"3d",	--138
		x"20",	--139
		x"3e",	--140
		x"88",	--141
		x"0f",	--142
		x"2f",	--143
		x"b0",	--144
		x"20",	--145
		x"0f",	--146
		x"2f",	--147
		x"b0",	--148
		x"68",	--149
		x"0e",	--150
		x"2e",	--151
		x"0f",	--152
		x"3f",	--153
		x"0e",	--154
		x"b0",	--155
		x"3c",	--156
		x"3e",	--157
		x"98",	--158
		x"0f",	--159
		x"2f",	--160
		x"b0",	--161
		x"6e",	--162
		x"3e",	--163
		x"9c",	--164
		x"0f",	--165
		x"b0",	--166
		x"6e",	--167
		x"0e",	--168
		x"0f",	--169
		x"2f",	--170
		x"b0",	--171
		x"5c",	--172
		x"b0",	--173
		x"46",	--174
		x"3e",	--175
		x"ff",	--176
		x"3f",	--177
		x"fc",	--178
		x"b0",	--179
		x"56",	--180
		x"0d",	--181
		x"3e",	--182
		x"e8",	--183
		x"b0",	--184
		x"9a",	--185
		x"0c",	--186
		x"0d",	--187
		x"1e",	--188
		x"0f",	--189
		x"3f",	--190
		x"24",	--191
		x"b0",	--192
		x"04",	--193
		x"0c",	--194
		x"0d",	--195
		x"1e",	--196
		x"0f",	--197
		x"3f",	--198
		x"18",	--199
		x"b0",	--200
		x"04",	--201
		x"0e",	--202
		x"3e",	--203
		x"18",	--204
		x"0f",	--205
		x"3f",	--206
		x"24",	--207
		x"b0",	--208
		x"cc",	--209
		x"f2",	--210
		x"80",	--211
		x"19",	--212
		x"32",	--213
		x"0b",	--214
		x"b0",	--215
		x"b6",	--216
		x"0f",	--217
		x"fc",	--218
		x"b0",	--219
		x"de",	--220
		x"7f",	--221
		x"15",	--222
		x"7f",	--223
		x"0d",	--224
		x"1b",	--225
		x"30",	--226
		x"bb",	--227
		x"b0",	--228
		x"5c",	--229
		x"21",	--230
		x"3f",	--231
		x"30",	--232
		x"0f",	--233
		x"0b",	--234
		x"cb",	--235
		x"00",	--236
		x"0e",	--237
		x"5f",	--238
		x"30",	--239
		x"b0",	--240
		x"ae",	--241
		x"0b",	--242
		x"e3",	--243
		x"0b",	--244
		x"e1",	--245
		x"3b",	--246
		x"30",	--247
		x"be",	--248
		x"b0",	--249
		x"5c",	--250
		x"21",	--251
		x"da",	--252
		x"3b",	--253
		x"28",	--254
		x"d7",	--255
		x"82",	--256
		x"0c",	--257
		x"0c",	--258
		x"4e",	--259
		x"8e",	--260
		x"0e",	--261
		x"30",	--262
		x"c2",	--263
		x"81",	--264
		x"5c",	--265
		x"b0",	--266
		x"5c",	--267
		x"21",	--268
		x"1f",	--269
		x"58",	--270
		x"3e",	--271
		x"30",	--272
		x"0e",	--273
		x"0e",	--274
		x"ce",	--275
		x"00",	--276
		x"1b",	--277
		x"c0",	--278
		x"30",	--279
		x"94",	--280
		x"8f",	--281
		x"00",	--282
		x"8f",	--283
		x"02",	--284
		x"8f",	--285
		x"04",	--286
		x"8f",	--287
		x"06",	--288
		x"8f",	--289
		x"08",	--290
		x"8f",	--291
		x"0a",	--292
		x"30",	--293
		x"8f",	--294
		x"06",	--295
		x"8f",	--296
		x"08",	--297
		x"8f",	--298
		x"0a",	--299
		x"30",	--300
		x"8f",	--301
		x"00",	--302
		x"30",	--303
		x"8f",	--304
		x"02",	--305
		x"30",	--306
		x"8f",	--307
		x"04",	--308
		x"30",	--309
		x"8f",	--310
		x"06",	--311
		x"30",	--312
		x"1d",	--313
		x"06",	--314
		x"0d",	--315
		x"0e",	--316
		x"1d",	--317
		x"08",	--318
		x"8f",	--319
		x"08",	--320
		x"02",	--321
		x"32",	--322
		x"03",	--323
		x"82",	--324
		x"32",	--325
		x"a2",	--326
		x"38",	--327
		x"1c",	--328
		x"3a",	--329
		x"32",	--330
		x"02",	--331
		x"32",	--332
		x"03",	--333
		x"82",	--334
		x"32",	--335
		x"92",	--336
		x"02",	--337
		x"38",	--338
		x"1d",	--339
		x"3a",	--340
		x"32",	--341
		x"0d",	--342
		x"1e",	--343
		x"0a",	--344
		x"02",	--345
		x"32",	--346
		x"03",	--347
		x"82",	--348
		x"32",	--349
		x"92",	--350
		x"04",	--351
		x"38",	--352
		x"1f",	--353
		x"3a",	--354
		x"32",	--355
		x"0f",	--356
		x"30",	--357
		x"30",	--358
		x"0f",	--359
		x"30",	--360
		x"0f",	--361
		x"30",	--362
		x"b2",	--363
		x"00",	--364
		x"92",	--365
		x"b2",	--366
		x"30",	--367
		x"94",	--368
		x"b2",	--369
		x"41",	--370
		x"96",	--371
		x"30",	--372
		x"9c",	--373
		x"b0",	--374
		x"5c",	--375
		x"92",	--376
		x"90",	--377
		x"b1",	--378
		x"ba",	--379
		x"00",	--380
		x"b0",	--381
		x"5c",	--382
		x"21",	--383
		x"0f",	--384
		x"30",	--385
		x"b0",	--386
		x"32",	--387
		x"30",	--388
		x"0b",	--389
		x"0a",	--390
		x"0a",	--391
		x"3b",	--392
		x"00",	--393
		x"0d",	--394
		x"0e",	--395
		x"1f",	--396
		x"1e",	--397
		x"b0",	--398
		x"bc",	--399
		x"0d",	--400
		x"0e",	--401
		x"1f",	--402
		x"1c",	--403
		x"b0",	--404
		x"bc",	--405
		x"30",	--406
		x"d3",	--407
		x"b0",	--408
		x"5c",	--409
		x"21",	--410
		x"3a",	--411
		x"3b",	--412
		x"30",	--413
		x"82",	--414
		x"1e",	--415
		x"82",	--416
		x"1c",	--417
		x"30",	--418
		x"0b",	--419
		x"0a",	--420
		x"21",	--421
		x"0a",	--422
		x"0b",	--423
		x"b2",	--424
		x"00",	--425
		x"47",	--426
		x"3a",	--427
		x"03",	--428
		x"4c",	--429
		x"37",	--430
		x"0e",	--431
		x"1f",	--432
		x"02",	--433
		x"b0",	--434
		x"52",	--435
		x"0a",	--436
		x"0e",	--437
		x"1f",	--438
		x"04",	--439
		x"b0",	--440
		x"52",	--441
		x"0b",	--442
		x"0f",	--443
		x"0a",	--444
		x"30",	--445
		x"20",	--446
		x"b0",	--447
		x"5c",	--448
		x"31",	--449
		x"06",	--450
		x"0e",	--451
		x"0f",	--452
		x"b0",	--453
		x"d0",	--454
		x"0c",	--455
		x"3d",	--456
		x"c8",	--457
		x"b0",	--458
		x"a0",	--459
		x"0d",	--460
		x"0e",	--461
		x"1f",	--462
		x"1e",	--463
		x"b0",	--464
		x"bc",	--465
		x"0e",	--466
		x"0f",	--467
		x"b0",	--468
		x"d0",	--469
		x"0c",	--470
		x"3d",	--471
		x"c8",	--472
		x"b0",	--473
		x"a0",	--474
		x"0d",	--475
		x"0e",	--476
		x"1f",	--477
		x"1c",	--478
		x"b0",	--479
		x"bc",	--480
		x"0f",	--481
		x"21",	--482
		x"3a",	--483
		x"3b",	--484
		x"30",	--485
		x"0e",	--486
		x"1f",	--487
		x"06",	--488
		x"b0",	--489
		x"52",	--490
		x"1d",	--491
		x"0e",	--492
		x"1f",	--493
		x"00",	--494
		x"b0",	--495
		x"9a",	--496
		x"bd",	--497
		x"0e",	--498
		x"3f",	--499
		x"0a",	--500
		x"b0",	--501
		x"56",	--502
		x"82",	--503
		x"00",	--504
		x"b1",	--505
		x"30",	--506
		x"da",	--507
		x"b0",	--508
		x"5c",	--509
		x"b1",	--510
		x"f4",	--511
		x"00",	--512
		x"b0",	--513
		x"5c",	--514
		x"a1",	--515
		x"00",	--516
		x"30",	--517
		x"05",	--518
		x"b0",	--519
		x"5c",	--520
		x"21",	--521
		x"3f",	--522
		x"d6",	--523
		x"0b",	--524
		x"0a",	--525
		x"1f",	--526
		x"22",	--527
		x"b0",	--528
		x"76",	--529
		x"0a",	--530
		x"0b",	--531
		x"1f",	--532
		x"20",	--533
		x"b0",	--534
		x"76",	--535
		x"0b",	--536
		x"0a",	--537
		x"0f",	--538
		x"0e",	--539
		x"30",	--540
		x"28",	--541
		x"30",	--542
		x"24",	--543
		x"b0",	--544
		x"28",	--545
		x"31",	--546
		x"0c",	--547
		x"30",	--548
		x"24",	--549
		x"30",	--550
		x"30",	--551
		x"b0",	--552
		x"5c",	--553
		x"21",	--554
		x"3a",	--555
		x"3b",	--556
		x"30",	--557
		x"82",	--558
		x"20",	--559
		x"82",	--560
		x"22",	--561
		x"30",	--562
		x"0b",	--563
		x"0a",	--564
		x"09",	--565
		x"21",	--566
		x"0a",	--567
		x"0b",	--568
		x"81",	--569
		x"00",	--570
		x"1f",	--571
		x"1a",	--572
		x"b2",	--573
		x"02",	--574
		x"36",	--575
		x"92",	--576
		x"0a",	--577
		x"0e",	--578
		x"1f",	--579
		x"02",	--580
		x"b0",	--581
		x"52",	--582
		x"09",	--583
		x"3a",	--584
		x"03",	--585
		x"1b",	--586
		x"0d",	--587
		x"0e",	--588
		x"1f",	--589
		x"02",	--590
		x"b0",	--591
		x"9a",	--592
		x"0f",	--593
		x"21",	--594
		x"39",	--595
		x"3a",	--596
		x"3b",	--597
		x"30",	--598
		x"82",	--599
		x"0a",	--600
		x"13",	--601
		x"82",	--602
		x"0a",	--603
		x"1f",	--604
		x"02",	--605
		x"b0",	--606
		x"c2",	--607
		x"0f",	--608
		x"21",	--609
		x"39",	--610
		x"3a",	--611
		x"3b",	--612
		x"30",	--613
		x"0e",	--614
		x"1f",	--615
		x"04",	--616
		x"b0",	--617
		x"52",	--618
		x"0d",	--619
		x"df",	--620
		x"0f",	--621
		x"b0",	--622
		x"18",	--623
		x"0f",	--624
		x"21",	--625
		x"39",	--626
		x"3a",	--627
		x"3b",	--628
		x"30",	--629
		x"0e",	--630
		x"3f",	--631
		x"18",	--632
		x"b0",	--633
		x"56",	--634
		x"82",	--635
		x"02",	--636
		x"c2",	--637
		x"5e",	--638
		x"19",	--639
		x"4e",	--640
		x"0f",	--641
		x"03",	--642
		x"c2",	--643
		x"19",	--644
		x"30",	--645
		x"c2",	--646
		x"19",	--647
		x"30",	--648
		x"1f",	--649
		x"82",	--650
		x"0c",	--651
		x"01",	--652
		x"0f",	--653
		x"82",	--654
		x"0c",	--655
		x"0f",	--656
		x"30",	--657
		x"1e",	--658
		x"0e",	--659
		x"3e",	--660
		x"06",	--661
		x"0f",	--662
		x"0f",	--663
		x"10",	--664
		x"36",	--665
		x"c2",	--666
		x"19",	--667
		x"3e",	--668
		x"07",	--669
		x"03",	--670
		x"82",	--671
		x"0e",	--672
		x"30",	--673
		x"1e",	--674
		x"82",	--675
		x"0e",	--676
		x"30",	--677
		x"f2",	--678
		x"0e",	--679
		x"19",	--680
		x"f2",	--681
		x"f2",	--682
		x"0a",	--683
		x"19",	--684
		x"ee",	--685
		x"e2",	--686
		x"19",	--687
		x"eb",	--688
		x"f2",	--689
		x"0d",	--690
		x"19",	--691
		x"e7",	--692
		x"f2",	--693
		x"09",	--694
		x"19",	--695
		x"e3",	--696
		x"f2",	--697
		x"03",	--698
		x"19",	--699
		x"df",	--700
		x"f2",	--701
		x"07",	--702
		x"19",	--703
		x"db",	--704
		x"0b",	--705
		x"0a",	--706
		x"21",	--707
		x"0a",	--708
		x"0b",	--709
		x"30",	--710
		x"c6",	--711
		x"b0",	--712
		x"5c",	--713
		x"21",	--714
		x"3a",	--715
		x"03",	--716
		x"1b",	--717
		x"0e",	--718
		x"1f",	--719
		x"02",	--720
		x"b0",	--721
		x"52",	--722
		x"0a",	--723
		x"0e",	--724
		x"1f",	--725
		x"04",	--726
		x"b0",	--727
		x"52",	--728
		x"0b",	--729
		x"0f",	--730
		x"0a",	--731
		x"30",	--732
		x"0e",	--733
		x"b0",	--734
		x"5c",	--735
		x"31",	--736
		x"06",	--737
		x"8a",	--738
		x"00",	--739
		x"0f",	--740
		x"21",	--741
		x"3a",	--742
		x"3b",	--743
		x"30",	--744
		x"30",	--745
		x"ce",	--746
		x"b0",	--747
		x"5c",	--748
		x"b1",	--749
		x"e8",	--750
		x"00",	--751
		x"b0",	--752
		x"5c",	--753
		x"a1",	--754
		x"00",	--755
		x"30",	--756
		x"f9",	--757
		x"b0",	--758
		x"5c",	--759
		x"21",	--760
		x"3f",	--761
		x"ea",	--762
		x"0b",	--763
		x"21",	--764
		x"0b",	--765
		x"1f",	--766
		x"17",	--767
		x"16",	--768
		x"30",	--769
		x"29",	--770
		x"b0",	--771
		x"5c",	--772
		x"21",	--773
		x"0e",	--774
		x"1f",	--775
		x"02",	--776
		x"b0",	--777
		x"52",	--778
		x"2f",	--779
		x"0f",	--780
		x"30",	--781
		x"0e",	--782
		x"b0",	--783
		x"5c",	--784
		x"31",	--785
		x"06",	--786
		x"0f",	--787
		x"21",	--788
		x"3b",	--789
		x"30",	--790
		x"30",	--791
		x"ce",	--792
		x"b0",	--793
		x"5c",	--794
		x"b1",	--795
		x"e8",	--796
		x"00",	--797
		x"b0",	--798
		x"5c",	--799
		x"a1",	--800
		x"00",	--801
		x"30",	--802
		x"1a",	--803
		x"b0",	--804
		x"5c",	--805
		x"21",	--806
		x"3f",	--807
		x"eb",	--808
		x"0b",	--809
		x"0a",	--810
		x"8e",	--811
		x"00",	--812
		x"6d",	--813
		x"4d",	--814
		x"5e",	--815
		x"1f",	--816
		x"0a",	--817
		x"0c",	--818
		x"0f",	--819
		x"7b",	--820
		x"0a",	--821
		x"2b",	--822
		x"0c",	--823
		x"0c",	--824
		x"0c",	--825
		x"0c",	--826
		x"8d",	--827
		x"0c",	--828
		x"3c",	--829
		x"d0",	--830
		x"1a",	--831
		x"7d",	--832
		x"4d",	--833
		x"17",	--834
		x"7d",	--835
		x"78",	--836
		x"1a",	--837
		x"4b",	--838
		x"7b",	--839
		x"d0",	--840
		x"0a",	--841
		x"e9",	--842
		x"7b",	--843
		x"0a",	--844
		x"34",	--845
		x"0c",	--846
		x"0b",	--847
		x"0b",	--848
		x"0b",	--849
		x"0c",	--850
		x"8d",	--851
		x"0c",	--852
		x"3c",	--853
		x"d0",	--854
		x"7d",	--855
		x"4d",	--856
		x"e9",	--857
		x"9e",	--858
		x"00",	--859
		x"0f",	--860
		x"3a",	--861
		x"3b",	--862
		x"30",	--863
		x"1a",	--864
		x"de",	--865
		x"4b",	--866
		x"7b",	--867
		x"9f",	--868
		x"7b",	--869
		x"06",	--870
		x"0a",	--871
		x"0c",	--872
		x"0c",	--873
		x"0c",	--874
		x"0c",	--875
		x"8d",	--876
		x"0c",	--877
		x"3c",	--878
		x"a9",	--879
		x"1a",	--880
		x"ce",	--881
		x"4b",	--882
		x"7b",	--883
		x"bf",	--884
		x"7b",	--885
		x"06",	--886
		x"0a",	--887
		x"0c",	--888
		x"0c",	--889
		x"0c",	--890
		x"0c",	--891
		x"8d",	--892
		x"0c",	--893
		x"3c",	--894
		x"c9",	--895
		x"1a",	--896
		x"be",	--897
		x"8d",	--898
		x"0d",	--899
		x"30",	--900
		x"30",	--901
		x"b0",	--902
		x"5c",	--903
		x"21",	--904
		x"0c",	--905
		x"0f",	--906
		x"3a",	--907
		x"3b",	--908
		x"30",	--909
		x"0c",	--910
		x"ca",	--911
		x"0b",	--912
		x"0a",	--913
		x"0b",	--914
		x"0a",	--915
		x"8f",	--916
		x"00",	--917
		x"8f",	--918
		x"02",	--919
		x"8f",	--920
		x"04",	--921
		x"0c",	--922
		x"0d",	--923
		x"3e",	--924
		x"00",	--925
		x"3f",	--926
		x"6e",	--927
		x"b0",	--928
		x"36",	--929
		x"8b",	--930
		x"02",	--931
		x"02",	--932
		x"32",	--933
		x"03",	--934
		x"82",	--935
		x"32",	--936
		x"b2",	--937
		x"18",	--938
		x"38",	--939
		x"9b",	--940
		x"3a",	--941
		x"06",	--942
		x"32",	--943
		x"0f",	--944
		x"3a",	--945
		x"3b",	--946
		x"30",	--947
		x"0b",	--948
		x"09",	--949
		x"08",	--950
		x"8f",	--951
		x"06",	--952
		x"bf",	--953
		x"00",	--954
		x"08",	--955
		x"2b",	--956
		x"1e",	--957
		x"02",	--958
		x"0f",	--959
		x"b0",	--960
		x"d0",	--961
		x"0c",	--962
		x"3d",	--963
		x"00",	--964
		x"b0",	--965
		x"7c",	--966
		x"08",	--967
		x"09",	--968
		x"1e",	--969
		x"06",	--970
		x"0f",	--971
		x"b0",	--972
		x"d0",	--973
		x"0c",	--974
		x"0d",	--975
		x"0e",	--976
		x"0f",	--977
		x"b0",	--978
		x"2c",	--979
		x"b0",	--980
		x"0c",	--981
		x"8b",	--982
		x"04",	--983
		x"9b",	--984
		x"00",	--985
		x"38",	--986
		x"39",	--987
		x"3b",	--988
		x"30",	--989
		x"0b",	--990
		x"0a",	--991
		x"09",	--992
		x"0a",	--993
		x"0b",	--994
		x"8f",	--995
		x"06",	--996
		x"8f",	--997
		x"08",	--998
		x"29",	--999
		x"1e",	--1000
		x"02",	--1001
		x"0f",	--1002
		x"b0",	--1003
		x"d0",	--1004
		x"0c",	--1005
		x"0d",	--1006
		x"0e",	--1007
		x"0f",	--1008
		x"b0",	--1009
		x"7c",	--1010
		x"0a",	--1011
		x"0b",	--1012
		x"1e",	--1013
		x"06",	--1014
		x"0f",	--1015
		x"b0",	--1016
		x"d0",	--1017
		x"0c",	--1018
		x"0d",	--1019
		x"0e",	--1020
		x"0f",	--1021
		x"b0",	--1022
		x"2c",	--1023
		x"b0",	--1024
		x"0c",	--1025
		x"89",	--1026
		x"04",	--1027
		x"39",	--1028
		x"3a",	--1029
		x"3b",	--1030
		x"30",	--1031
		x"0b",	--1032
		x"0a",	--1033
		x"92",	--1034
		x"10",	--1035
		x"14",	--1036
		x"3b",	--1037
		x"68",	--1038
		x"0a",	--1039
		x"2b",	--1040
		x"5f",	--1041
		x"fc",	--1042
		x"8f",	--1043
		x"0f",	--1044
		x"30",	--1045
		x"45",	--1046
		x"b0",	--1047
		x"5c",	--1048
		x"31",	--1049
		x"06",	--1050
		x"1a",	--1051
		x"3b",	--1052
		x"06",	--1053
		x"1a",	--1054
		x"10",	--1055
		x"ef",	--1056
		x"0f",	--1057
		x"3a",	--1058
		x"3b",	--1059
		x"30",	--1060
		x"1e",	--1061
		x"10",	--1062
		x"3e",	--1063
		x"20",	--1064
		x"12",	--1065
		x"0f",	--1066
		x"0f",	--1067
		x"0f",	--1068
		x"0f",	--1069
		x"3f",	--1070
		x"64",	--1071
		x"ff",	--1072
		x"68",	--1073
		x"00",	--1074
		x"bf",	--1075
		x"10",	--1076
		x"02",	--1077
		x"bf",	--1078
		x"04",	--1079
		x"04",	--1080
		x"1e",	--1081
		x"82",	--1082
		x"10",	--1083
		x"30",	--1084
		x"0b",	--1085
		x"1b",	--1086
		x"10",	--1087
		x"3b",	--1088
		x"20",	--1089
		x"12",	--1090
		x"0c",	--1091
		x"0c",	--1092
		x"0c",	--1093
		x"0c",	--1094
		x"3c",	--1095
		x"64",	--1096
		x"cc",	--1097
		x"00",	--1098
		x"8c",	--1099
		x"02",	--1100
		x"8c",	--1101
		x"04",	--1102
		x"1b",	--1103
		x"82",	--1104
		x"10",	--1105
		x"0f",	--1106
		x"3b",	--1107
		x"30",	--1108
		x"3f",	--1109
		x"fc",	--1110
		x"0b",	--1111
		x"31",	--1112
		x"f0",	--1113
		x"1b",	--1114
		x"10",	--1115
		x"1b",	--1116
		x"0f",	--1117
		x"5f",	--1118
		x"64",	--1119
		x"16",	--1120
		x"3d",	--1121
		x"6a",	--1122
		x"0c",	--1123
		x"05",	--1124
		x"3d",	--1125
		x"06",	--1126
		x"cd",	--1127
		x"fa",	--1128
		x"0e",	--1129
		x"1c",	--1130
		x"0c",	--1131
		x"f8",	--1132
		x"30",	--1133
		x"4d",	--1134
		x"b0",	--1135
		x"5c",	--1136
		x"21",	--1137
		x"3f",	--1138
		x"31",	--1139
		x"10",	--1140
		x"3b",	--1141
		x"30",	--1142
		x"0c",	--1143
		x"81",	--1144
		x"00",	--1145
		x"6d",	--1146
		x"4d",	--1147
		x"24",	--1148
		x"1e",	--1149
		x"1f",	--1150
		x"06",	--1151
		x"6d",	--1152
		x"4d",	--1153
		x"11",	--1154
		x"1e",	--1155
		x"3f",	--1156
		x"0e",	--1157
		x"7d",	--1158
		x"20",	--1159
		x"f7",	--1160
		x"ce",	--1161
		x"ff",	--1162
		x"0d",	--1163
		x"0d",	--1164
		x"0d",	--1165
		x"8d",	--1166
		x"00",	--1167
		x"1f",	--1168
		x"6d",	--1169
		x"4d",	--1170
		x"ef",	--1171
		x"0e",	--1172
		x"0e",	--1173
		x"0c",	--1174
		x"0c",	--1175
		x"3c",	--1176
		x"64",	--1177
		x"0e",	--1178
		x"9c",	--1179
		x"02",	--1180
		x"31",	--1181
		x"10",	--1182
		x"3b",	--1183
		x"30",	--1184
		x"1f",	--1185
		x"f1",	--1186
		x"b2",	--1187
		x"d2",	--1188
		x"60",	--1189
		x"b2",	--1190
		x"b8",	--1191
		x"72",	--1192
		x"0f",	--1193
		x"30",	--1194
		x"0b",	--1195
		x"0b",	--1196
		x"1f",	--1197
		x"12",	--1198
		x"3f",	--1199
		x"20",	--1200
		x"19",	--1201
		x"0c",	--1202
		x"0c",	--1203
		x"0d",	--1204
		x"0d",	--1205
		x"0d",	--1206
		x"0d",	--1207
		x"0d",	--1208
		x"3d",	--1209
		x"24",	--1210
		x"8d",	--1211
		x"00",	--1212
		x"8d",	--1213
		x"02",	--1214
		x"8d",	--1215
		x"08",	--1216
		x"8d",	--1217
		x"0a",	--1218
		x"8d",	--1219
		x"0c",	--1220
		x"0e",	--1221
		x"1e",	--1222
		x"82",	--1223
		x"12",	--1224
		x"3b",	--1225
		x"30",	--1226
		x"3f",	--1227
		x"fc",	--1228
		x"0f",	--1229
		x"0c",	--1230
		x"0c",	--1231
		x"0c",	--1232
		x"0c",	--1233
		x"0c",	--1234
		x"3c",	--1235
		x"24",	--1236
		x"8c",	--1237
		x"02",	--1238
		x"8c",	--1239
		x"04",	--1240
		x"8c",	--1241
		x"06",	--1242
		x"8c",	--1243
		x"08",	--1244
		x"9c",	--1245
		x"00",	--1246
		x"0f",	--1247
		x"30",	--1248
		x"0f",	--1249
		x"0e",	--1250
		x"0e",	--1251
		x"0e",	--1252
		x"0e",	--1253
		x"0e",	--1254
		x"8e",	--1255
		x"24",	--1256
		x"0f",	--1257
		x"30",	--1258
		x"0f",	--1259
		x"0e",	--1260
		x"0d",	--1261
		x"0c",	--1262
		x"0b",	--1263
		x"0a",	--1264
		x"09",	--1265
		x"08",	--1266
		x"07",	--1267
		x"92",	--1268
		x"12",	--1269
		x"33",	--1270
		x"3a",	--1271
		x"24",	--1272
		x"0b",	--1273
		x"2b",	--1274
		x"08",	--1275
		x"38",	--1276
		x"07",	--1277
		x"37",	--1278
		x"06",	--1279
		x"09",	--1280
		x"0f",	--1281
		x"1f",	--1282
		x"8b",	--1283
		x"00",	--1284
		x"19",	--1285
		x"3a",	--1286
		x"0e",	--1287
		x"3b",	--1288
		x"0e",	--1289
		x"38",	--1290
		x"0e",	--1291
		x"37",	--1292
		x"0e",	--1293
		x"19",	--1294
		x"12",	--1295
		x"19",	--1296
		x"8a",	--1297
		x"00",	--1298
		x"f1",	--1299
		x"2f",	--1300
		x"1f",	--1301
		x"02",	--1302
		x"ea",	--1303
		x"8b",	--1304
		x"00",	--1305
		x"1f",	--1306
		x"0a",	--1307
		x"9b",	--1308
		x"08",	--1309
		x"88",	--1310
		x"00",	--1311
		x"e4",	--1312
		x"2f",	--1313
		x"1f",	--1314
		x"87",	--1315
		x"00",	--1316
		x"2f",	--1317
		x"de",	--1318
		x"8a",	--1319
		x"00",	--1320
		x"db",	--1321
		x"b2",	--1322
		x"fe",	--1323
		x"60",	--1324
		x"37",	--1325
		x"38",	--1326
		x"39",	--1327
		x"3a",	--1328
		x"3b",	--1329
		x"3c",	--1330
		x"3d",	--1331
		x"3e",	--1332
		x"3f",	--1333
		x"00",	--1334
		x"8f",	--1335
		x"00",	--1336
		x"0f",	--1337
		x"30",	--1338
		x"2f",	--1339
		x"2e",	--1340
		x"1f",	--1341
		x"02",	--1342
		x"30",	--1343
		x"5e",	--1344
		x"81",	--1345
		x"3e",	--1346
		x"fc",	--1347
		x"c2",	--1348
		x"84",	--1349
		x"0f",	--1350
		x"30",	--1351
		x"3f",	--1352
		x"0f",	--1353
		x"5f",	--1354
		x"0c",	--1355
		x"8f",	--1356
		x"b0",	--1357
		x"80",	--1358
		x"30",	--1359
		x"0b",	--1360
		x"0b",	--1361
		x"0e",	--1362
		x"0e",	--1363
		x"0e",	--1364
		x"0e",	--1365
		x"0e",	--1366
		x"0f",	--1367
		x"b0",	--1368
		x"90",	--1369
		x"0f",	--1370
		x"b0",	--1371
		x"90",	--1372
		x"3b",	--1373
		x"30",	--1374
		x"0b",	--1375
		x"0a",	--1376
		x"0a",	--1377
		x"3b",	--1378
		x"07",	--1379
		x"0e",	--1380
		x"4d",	--1381
		x"7d",	--1382
		x"0f",	--1383
		x"03",	--1384
		x"0e",	--1385
		x"7d",	--1386
		x"fd",	--1387
		x"1e",	--1388
		x"0a",	--1389
		x"3f",	--1390
		x"31",	--1391
		x"b0",	--1392
		x"80",	--1393
		x"3b",	--1394
		x"3b",	--1395
		x"ef",	--1396
		x"3a",	--1397
		x"3b",	--1398
		x"30",	--1399
		x"3f",	--1400
		x"30",	--1401
		x"f5",	--1402
		x"0b",	--1403
		x"0b",	--1404
		x"0e",	--1405
		x"8e",	--1406
		x"8e",	--1407
		x"0f",	--1408
		x"b0",	--1409
		x"a0",	--1410
		x"0f",	--1411
		x"b0",	--1412
		x"a0",	--1413
		x"3b",	--1414
		x"30",	--1415
		x"0b",	--1416
		x"0a",	--1417
		x"0a",	--1418
		x"0b",	--1419
		x"0d",	--1420
		x"8d",	--1421
		x"8d",	--1422
		x"0f",	--1423
		x"b0",	--1424
		x"a0",	--1425
		x"0f",	--1426
		x"b0",	--1427
		x"a0",	--1428
		x"0c",	--1429
		x"0d",	--1430
		x"8d",	--1431
		x"8c",	--1432
		x"4d",	--1433
		x"0d",	--1434
		x"0f",	--1435
		x"b0",	--1436
		x"a0",	--1437
		x"0f",	--1438
		x"b0",	--1439
		x"a0",	--1440
		x"3a",	--1441
		x"3b",	--1442
		x"30",	--1443
		x"0b",	--1444
		x"0a",	--1445
		x"09",	--1446
		x"0a",	--1447
		x"0e",	--1448
		x"19",	--1449
		x"09",	--1450
		x"39",	--1451
		x"0b",	--1452
		x"0d",	--1453
		x"0d",	--1454
		x"6f",	--1455
		x"8f",	--1456
		x"b0",	--1457
		x"a0",	--1458
		x"0b",	--1459
		x"0e",	--1460
		x"1b",	--1461
		x"3b",	--1462
		x"07",	--1463
		x"05",	--1464
		x"3f",	--1465
		x"20",	--1466
		x"b0",	--1467
		x"80",	--1468
		x"ef",	--1469
		x"3f",	--1470
		x"3a",	--1471
		x"b0",	--1472
		x"80",	--1473
		x"ea",	--1474
		x"39",	--1475
		x"3a",	--1476
		x"3b",	--1477
		x"30",	--1478
		x"0b",	--1479
		x"0a",	--1480
		x"09",	--1481
		x"0a",	--1482
		x"0e",	--1483
		x"17",	--1484
		x"09",	--1485
		x"39",	--1486
		x"0b",	--1487
		x"6f",	--1488
		x"8f",	--1489
		x"b0",	--1490
		x"90",	--1491
		x"0b",	--1492
		x"0e",	--1493
		x"1b",	--1494
		x"3b",	--1495
		x"07",	--1496
		x"f6",	--1497
		x"3f",	--1498
		x"20",	--1499
		x"b0",	--1500
		x"80",	--1501
		x"6f",	--1502
		x"8f",	--1503
		x"b0",	--1504
		x"90",	--1505
		x"0b",	--1506
		x"f2",	--1507
		x"39",	--1508
		x"3a",	--1509
		x"3b",	--1510
		x"30",	--1511
		x"0b",	--1512
		x"0a",	--1513
		x"09",	--1514
		x"31",	--1515
		x"ec",	--1516
		x"0b",	--1517
		x"0f",	--1518
		x"34",	--1519
		x"3b",	--1520
		x"0a",	--1521
		x"38",	--1522
		x"09",	--1523
		x"0a",	--1524
		x"0a",	--1525
		x"3e",	--1526
		x"0a",	--1527
		x"0f",	--1528
		x"b0",	--1529
		x"ee",	--1530
		x"7f",	--1531
		x"30",	--1532
		x"ca",	--1533
		x"00",	--1534
		x"19",	--1535
		x"3e",	--1536
		x"0a",	--1537
		x"0f",	--1538
		x"b0",	--1539
		x"bc",	--1540
		x"0b",	--1541
		x"3f",	--1542
		x"0a",	--1543
		x"eb",	--1544
		x"0a",	--1545
		x"1a",	--1546
		x"09",	--1547
		x"3e",	--1548
		x"0a",	--1549
		x"0f",	--1550
		x"b0",	--1551
		x"ee",	--1552
		x"7f",	--1553
		x"30",	--1554
		x"c9",	--1555
		x"00",	--1556
		x"3a",	--1557
		x"0f",	--1558
		x"0f",	--1559
		x"6f",	--1560
		x"8f",	--1561
		x"b0",	--1562
		x"80",	--1563
		x"0a",	--1564
		x"f7",	--1565
		x"31",	--1566
		x"14",	--1567
		x"39",	--1568
		x"3a",	--1569
		x"3b",	--1570
		x"30",	--1571
		x"3f",	--1572
		x"2d",	--1573
		x"b0",	--1574
		x"80",	--1575
		x"3b",	--1576
		x"1b",	--1577
		x"c5",	--1578
		x"1a",	--1579
		x"09",	--1580
		x"dd",	--1581
		x"0b",	--1582
		x"0a",	--1583
		x"09",	--1584
		x"0b",	--1585
		x"3b",	--1586
		x"39",	--1587
		x"6f",	--1588
		x"4f",	--1589
		x"0b",	--1590
		x"1a",	--1591
		x"8f",	--1592
		x"b0",	--1593
		x"80",	--1594
		x"0a",	--1595
		x"09",	--1596
		x"19",	--1597
		x"5f",	--1598
		x"01",	--1599
		x"4f",	--1600
		x"10",	--1601
		x"7f",	--1602
		x"25",	--1603
		x"f3",	--1604
		x"0a",	--1605
		x"1a",	--1606
		x"5f",	--1607
		x"01",	--1608
		x"7f",	--1609
		x"db",	--1610
		x"7f",	--1611
		x"54",	--1612
		x"ee",	--1613
		x"4f",	--1614
		x"0f",	--1615
		x"10",	--1616
		x"64",	--1617
		x"39",	--1618
		x"3a",	--1619
		x"3b",	--1620
		x"30",	--1621
		x"09",	--1622
		x"29",	--1623
		x"1e",	--1624
		x"02",	--1625
		x"2f",	--1626
		x"b0",	--1627
		x"48",	--1628
		x"0b",	--1629
		x"dd",	--1630
		x"09",	--1631
		x"29",	--1632
		x"2f",	--1633
		x"b0",	--1634
		x"f6",	--1635
		x"0b",	--1636
		x"d6",	--1637
		x"0f",	--1638
		x"2b",	--1639
		x"29",	--1640
		x"6f",	--1641
		x"4f",	--1642
		x"d0",	--1643
		x"19",	--1644
		x"8f",	--1645
		x"b0",	--1646
		x"80",	--1647
		x"7f",	--1648
		x"4f",	--1649
		x"fa",	--1650
		x"c8",	--1651
		x"09",	--1652
		x"29",	--1653
		x"1e",	--1654
		x"02",	--1655
		x"2f",	--1656
		x"b0",	--1657
		x"8e",	--1658
		x"0b",	--1659
		x"bf",	--1660
		x"09",	--1661
		x"29",	--1662
		x"2e",	--1663
		x"0f",	--1664
		x"8f",	--1665
		x"8f",	--1666
		x"8f",	--1667
		x"8f",	--1668
		x"b0",	--1669
		x"10",	--1670
		x"0b",	--1671
		x"b3",	--1672
		x"09",	--1673
		x"29",	--1674
		x"2f",	--1675
		x"b0",	--1676
		x"d0",	--1677
		x"0b",	--1678
		x"ac",	--1679
		x"09",	--1680
		x"29",	--1681
		x"2f",	--1682
		x"b0",	--1683
		x"80",	--1684
		x"0b",	--1685
		x"a5",	--1686
		x"09",	--1687
		x"29",	--1688
		x"2f",	--1689
		x"b0",	--1690
		x"a0",	--1691
		x"0b",	--1692
		x"9e",	--1693
		x"09",	--1694
		x"29",	--1695
		x"2f",	--1696
		x"b0",	--1697
		x"be",	--1698
		x"0b",	--1699
		x"97",	--1700
		x"3f",	--1701
		x"25",	--1702
		x"b0",	--1703
		x"80",	--1704
		x"92",	--1705
		x"0f",	--1706
		x"0e",	--1707
		x"1f",	--1708
		x"14",	--1709
		x"df",	--1710
		x"85",	--1711
		x"e4",	--1712
		x"1f",	--1713
		x"14",	--1714
		x"3f",	--1715
		x"3f",	--1716
		x"13",	--1717
		x"92",	--1718
		x"14",	--1719
		x"1e",	--1720
		x"14",	--1721
		x"1f",	--1722
		x"16",	--1723
		x"0e",	--1724
		x"02",	--1725
		x"92",	--1726
		x"16",	--1727
		x"f2",	--1728
		x"10",	--1729
		x"81",	--1730
		x"3e",	--1731
		x"3f",	--1732
		x"b1",	--1733
		x"f0",	--1734
		x"00",	--1735
		x"00",	--1736
		x"82",	--1737
		x"14",	--1738
		x"ec",	--1739
		x"0c",	--1740
		x"0d",	--1741
		x"3e",	--1742
		x"00",	--1743
		x"3f",	--1744
		x"6e",	--1745
		x"b0",	--1746
		x"f6",	--1747
		x"3e",	--1748
		x"82",	--1749
		x"82",	--1750
		x"f2",	--1751
		x"11",	--1752
		x"80",	--1753
		x"30",	--1754
		x"1e",	--1755
		x"14",	--1756
		x"1f",	--1757
		x"16",	--1758
		x"0e",	--1759
		x"05",	--1760
		x"1f",	--1761
		x"14",	--1762
		x"1f",	--1763
		x"16",	--1764
		x"30",	--1765
		x"1d",	--1766
		x"14",	--1767
		x"1e",	--1768
		x"16",	--1769
		x"3f",	--1770
		x"40",	--1771
		x"0f",	--1772
		x"0f",	--1773
		x"30",	--1774
		x"1f",	--1775
		x"16",	--1776
		x"5f",	--1777
		x"e4",	--1778
		x"1d",	--1779
		x"16",	--1780
		x"1e",	--1781
		x"14",	--1782
		x"0d",	--1783
		x"0b",	--1784
		x"1e",	--1785
		x"16",	--1786
		x"3e",	--1787
		x"3f",	--1788
		x"03",	--1789
		x"82",	--1790
		x"16",	--1791
		x"30",	--1792
		x"92",	--1793
		x"16",	--1794
		x"30",	--1795
		x"4f",	--1796
		x"30",	--1797
		x"0b",	--1798
		x"0a",	--1799
		x"0a",	--1800
		x"0b",	--1801
		x"0c",	--1802
		x"3d",	--1803
		x"00",	--1804
		x"b0",	--1805
		x"f0",	--1806
		x"0f",	--1807
		x"07",	--1808
		x"0e",	--1809
		x"0f",	--1810
		x"b0",	--1811
		x"40",	--1812
		x"3a",	--1813
		x"3b",	--1814
		x"30",	--1815
		x"0c",	--1816
		x"3d",	--1817
		x"00",	--1818
		x"0e",	--1819
		x"0f",	--1820
		x"b0",	--1821
		x"2c",	--1822
		x"b0",	--1823
		x"40",	--1824
		x"0e",	--1825
		x"3f",	--1826
		x"00",	--1827
		x"3a",	--1828
		x"3b",	--1829
		x"30",	--1830
		x"0b",	--1831
		x"0a",	--1832
		x"09",	--1833
		x"08",	--1834
		x"07",	--1835
		x"06",	--1836
		x"05",	--1837
		x"04",	--1838
		x"31",	--1839
		x"fa",	--1840
		x"08",	--1841
		x"6b",	--1842
		x"6b",	--1843
		x"67",	--1844
		x"6c",	--1845
		x"6c",	--1846
		x"e9",	--1847
		x"6b",	--1848
		x"02",	--1849
		x"30",	--1850
		x"ce",	--1851
		x"6c",	--1852
		x"e3",	--1853
		x"6c",	--1854
		x"bb",	--1855
		x"6b",	--1856
		x"df",	--1857
		x"91",	--1858
		x"02",	--1859
		x"00",	--1860
		x"1b",	--1861
		x"02",	--1862
		x"14",	--1863
		x"04",	--1864
		x"15",	--1865
		x"06",	--1866
		x"16",	--1867
		x"04",	--1868
		x"17",	--1869
		x"06",	--1870
		x"2c",	--1871
		x"0c",	--1872
		x"09",	--1873
		x"0c",	--1874
		x"bf",	--1875
		x"39",	--1876
		x"20",	--1877
		x"50",	--1878
		x"1c",	--1879
		x"d7",	--1880
		x"81",	--1881
		x"02",	--1882
		x"81",	--1883
		x"04",	--1884
		x"4c",	--1885
		x"7c",	--1886
		x"1f",	--1887
		x"0b",	--1888
		x"0a",	--1889
		x"0b",	--1890
		x"12",	--1891
		x"0b",	--1892
		x"0a",	--1893
		x"7c",	--1894
		x"fb",	--1895
		x"81",	--1896
		x"02",	--1897
		x"81",	--1898
		x"04",	--1899
		x"1c",	--1900
		x"0d",	--1901
		x"79",	--1902
		x"1f",	--1903
		x"04",	--1904
		x"0c",	--1905
		x"0d",	--1906
		x"79",	--1907
		x"fc",	--1908
		x"3c",	--1909
		x"3d",	--1910
		x"0c",	--1911
		x"0d",	--1912
		x"1a",	--1913
		x"0b",	--1914
		x"0c",	--1915
		x"02",	--1916
		x"0d",	--1917
		x"e5",	--1918
		x"16",	--1919
		x"02",	--1920
		x"17",	--1921
		x"04",	--1922
		x"06",	--1923
		x"07",	--1924
		x"5f",	--1925
		x"01",	--1926
		x"5f",	--1927
		x"01",	--1928
		x"28",	--1929
		x"c8",	--1930
		x"01",	--1931
		x"a8",	--1932
		x"02",	--1933
		x"0e",	--1934
		x"0f",	--1935
		x"0e",	--1936
		x"0f",	--1937
		x"88",	--1938
		x"04",	--1939
		x"88",	--1940
		x"06",	--1941
		x"f8",	--1942
		x"03",	--1943
		x"00",	--1944
		x"0f",	--1945
		x"4d",	--1946
		x"0f",	--1947
		x"31",	--1948
		x"06",	--1949
		x"34",	--1950
		x"35",	--1951
		x"36",	--1952
		x"37",	--1953
		x"38",	--1954
		x"39",	--1955
		x"3a",	--1956
		x"3b",	--1957
		x"30",	--1958
		x"2b",	--1959
		x"67",	--1960
		x"81",	--1961
		x"00",	--1962
		x"04",	--1963
		x"05",	--1964
		x"5f",	--1965
		x"01",	--1966
		x"5f",	--1967
		x"01",	--1968
		x"d8",	--1969
		x"4f",	--1970
		x"68",	--1971
		x"0e",	--1972
		x"0f",	--1973
		x"0e",	--1974
		x"0f",	--1975
		x"0f",	--1976
		x"69",	--1977
		x"c8",	--1978
		x"01",	--1979
		x"a8",	--1980
		x"02",	--1981
		x"88",	--1982
		x"04",	--1983
		x"88",	--1984
		x"06",	--1985
		x"0c",	--1986
		x"0d",	--1987
		x"3c",	--1988
		x"3d",	--1989
		x"3d",	--1990
		x"ff",	--1991
		x"05",	--1992
		x"3d",	--1993
		x"00",	--1994
		x"17",	--1995
		x"3c",	--1996
		x"15",	--1997
		x"1b",	--1998
		x"02",	--1999
		x"3b",	--2000
		x"0e",	--2001
		x"0f",	--2002
		x"0a",	--2003
		x"3b",	--2004
		x"0c",	--2005
		x"0d",	--2006
		x"3c",	--2007
		x"3d",	--2008
		x"3d",	--2009
		x"ff",	--2010
		x"f5",	--2011
		x"3c",	--2012
		x"88",	--2013
		x"04",	--2014
		x"88",	--2015
		x"06",	--2016
		x"88",	--2017
		x"02",	--2018
		x"f8",	--2019
		x"03",	--2020
		x"00",	--2021
		x"0f",	--2022
		x"b3",	--2023
		x"0c",	--2024
		x"0d",	--2025
		x"1c",	--2026
		x"0d",	--2027
		x"12",	--2028
		x"0f",	--2029
		x"0e",	--2030
		x"0a",	--2031
		x"0b",	--2032
		x"0a",	--2033
		x"0b",	--2034
		x"88",	--2035
		x"04",	--2036
		x"88",	--2037
		x"06",	--2038
		x"98",	--2039
		x"02",	--2040
		x"0f",	--2041
		x"a1",	--2042
		x"6b",	--2043
		x"9f",	--2044
		x"ad",	--2045
		x"00",	--2046
		x"9d",	--2047
		x"02",	--2048
		x"02",	--2049
		x"9d",	--2050
		x"04",	--2051
		x"04",	--2052
		x"9d",	--2053
		x"06",	--2054
		x"06",	--2055
		x"5e",	--2056
		x"01",	--2057
		x"5e",	--2058
		x"01",	--2059
		x"cd",	--2060
		x"01",	--2061
		x"0f",	--2062
		x"8c",	--2063
		x"06",	--2064
		x"07",	--2065
		x"9a",	--2066
		x"39",	--2067
		x"19",	--2068
		x"39",	--2069
		x"20",	--2070
		x"8f",	--2071
		x"3e",	--2072
		x"3c",	--2073
		x"b6",	--2074
		x"c1",	--2075
		x"0e",	--2076
		x"0f",	--2077
		x"0e",	--2078
		x"0f",	--2079
		x"97",	--2080
		x"0f",	--2081
		x"79",	--2082
		x"d8",	--2083
		x"01",	--2084
		x"a8",	--2085
		x"02",	--2086
		x"3e",	--2087
		x"3f",	--2088
		x"1e",	--2089
		x"0f",	--2090
		x"88",	--2091
		x"04",	--2092
		x"88",	--2093
		x"06",	--2094
		x"92",	--2095
		x"0c",	--2096
		x"7b",	--2097
		x"81",	--2098
		x"00",	--2099
		x"81",	--2100
		x"02",	--2101
		x"81",	--2102
		x"04",	--2103
		x"4d",	--2104
		x"7d",	--2105
		x"1f",	--2106
		x"0c",	--2107
		x"4b",	--2108
		x"0c",	--2109
		x"0d",	--2110
		x"12",	--2111
		x"0d",	--2112
		x"0c",	--2113
		x"7b",	--2114
		x"fb",	--2115
		x"81",	--2116
		x"02",	--2117
		x"81",	--2118
		x"04",	--2119
		x"1c",	--2120
		x"0d",	--2121
		x"79",	--2122
		x"1f",	--2123
		x"04",	--2124
		x"0c",	--2125
		x"0d",	--2126
		x"79",	--2127
		x"fc",	--2128
		x"3c",	--2129
		x"3d",	--2130
		x"0c",	--2131
		x"0d",	--2132
		x"1a",	--2133
		x"0b",	--2134
		x"0c",	--2135
		x"04",	--2136
		x"0d",	--2137
		x"02",	--2138
		x"0a",	--2139
		x"0b",	--2140
		x"14",	--2141
		x"02",	--2142
		x"15",	--2143
		x"04",	--2144
		x"04",	--2145
		x"05",	--2146
		x"49",	--2147
		x"0a",	--2148
		x"0b",	--2149
		x"18",	--2150
		x"6c",	--2151
		x"33",	--2152
		x"df",	--2153
		x"01",	--2154
		x"01",	--2155
		x"2f",	--2156
		x"3f",	--2157
		x"1e",	--2158
		x"2c",	--2159
		x"31",	--2160
		x"e0",	--2161
		x"81",	--2162
		x"04",	--2163
		x"81",	--2164
		x"06",	--2165
		x"81",	--2166
		x"00",	--2167
		x"81",	--2168
		x"02",	--2169
		x"0e",	--2170
		x"3e",	--2171
		x"18",	--2172
		x"0f",	--2173
		x"2f",	--2174
		x"b0",	--2175
		x"02",	--2176
		x"0e",	--2177
		x"3e",	--2178
		x"10",	--2179
		x"0f",	--2180
		x"b0",	--2181
		x"02",	--2182
		x"0d",	--2183
		x"3d",	--2184
		x"0e",	--2185
		x"3e",	--2186
		x"10",	--2187
		x"0f",	--2188
		x"3f",	--2189
		x"18",	--2190
		x"b0",	--2191
		x"4e",	--2192
		x"b0",	--2193
		x"24",	--2194
		x"31",	--2195
		x"20",	--2196
		x"30",	--2197
		x"31",	--2198
		x"e0",	--2199
		x"81",	--2200
		x"04",	--2201
		x"81",	--2202
		x"06",	--2203
		x"81",	--2204
		x"00",	--2205
		x"81",	--2206
		x"02",	--2207
		x"0e",	--2208
		x"3e",	--2209
		x"18",	--2210
		x"0f",	--2211
		x"2f",	--2212
		x"b0",	--2213
		x"02",	--2214
		x"0e",	--2215
		x"3e",	--2216
		x"10",	--2217
		x"0f",	--2218
		x"b0",	--2219
		x"02",	--2220
		x"d1",	--2221
		x"11",	--2222
		x"0d",	--2223
		x"3d",	--2224
		x"0e",	--2225
		x"3e",	--2226
		x"10",	--2227
		x"0f",	--2228
		x"3f",	--2229
		x"18",	--2230
		x"b0",	--2231
		x"4e",	--2232
		x"b0",	--2233
		x"24",	--2234
		x"31",	--2235
		x"20",	--2236
		x"30",	--2237
		x"0b",	--2238
		x"0a",	--2239
		x"09",	--2240
		x"08",	--2241
		x"07",	--2242
		x"06",	--2243
		x"05",	--2244
		x"04",	--2245
		x"31",	--2246
		x"dc",	--2247
		x"81",	--2248
		x"04",	--2249
		x"81",	--2250
		x"06",	--2251
		x"81",	--2252
		x"00",	--2253
		x"81",	--2254
		x"02",	--2255
		x"0e",	--2256
		x"3e",	--2257
		x"18",	--2258
		x"0f",	--2259
		x"2f",	--2260
		x"b0",	--2261
		x"02",	--2262
		x"0e",	--2263
		x"3e",	--2264
		x"10",	--2265
		x"0f",	--2266
		x"b0",	--2267
		x"02",	--2268
		x"5f",	--2269
		x"18",	--2270
		x"6f",	--2271
		x"b6",	--2272
		x"5e",	--2273
		x"10",	--2274
		x"6e",	--2275
		x"d9",	--2276
		x"6f",	--2277
		x"ae",	--2278
		x"6e",	--2279
		x"e2",	--2280
		x"6f",	--2281
		x"ac",	--2282
		x"6e",	--2283
		x"d1",	--2284
		x"14",	--2285
		x"1c",	--2286
		x"15",	--2287
		x"1e",	--2288
		x"18",	--2289
		x"14",	--2290
		x"19",	--2291
		x"16",	--2292
		x"3c",	--2293
		x"20",	--2294
		x"0e",	--2295
		x"0f",	--2296
		x"06",	--2297
		x"07",	--2298
		x"81",	--2299
		x"20",	--2300
		x"81",	--2301
		x"22",	--2302
		x"0a",	--2303
		x"0b",	--2304
		x"81",	--2305
		x"20",	--2306
		x"08",	--2307
		x"08",	--2308
		x"09",	--2309
		x"12",	--2310
		x"05",	--2311
		x"04",	--2312
		x"b1",	--2313
		x"20",	--2314
		x"19",	--2315
		x"14",	--2316
		x"0d",	--2317
		x"0a",	--2318
		x"0b",	--2319
		x"0e",	--2320
		x"0f",	--2321
		x"1c",	--2322
		x"0d",	--2323
		x"0b",	--2324
		x"03",	--2325
		x"0b",	--2326
		x"0c",	--2327
		x"0d",	--2328
		x"0e",	--2329
		x"0f",	--2330
		x"06",	--2331
		x"07",	--2332
		x"09",	--2333
		x"e5",	--2334
		x"16",	--2335
		x"07",	--2336
		x"e2",	--2337
		x"0a",	--2338
		x"f5",	--2339
		x"f2",	--2340
		x"81",	--2341
		x"20",	--2342
		x"81",	--2343
		x"22",	--2344
		x"0c",	--2345
		x"1a",	--2346
		x"1a",	--2347
		x"1a",	--2348
		x"12",	--2349
		x"06",	--2350
		x"26",	--2351
		x"81",	--2352
		x"0a",	--2353
		x"5d",	--2354
		x"d1",	--2355
		x"11",	--2356
		x"19",	--2357
		x"83",	--2358
		x"c1",	--2359
		x"09",	--2360
		x"0c",	--2361
		x"3c",	--2362
		x"3f",	--2363
		x"00",	--2364
		x"18",	--2365
		x"1d",	--2366
		x"0a",	--2367
		x"3d",	--2368
		x"1a",	--2369
		x"20",	--2370
		x"1b",	--2371
		x"22",	--2372
		x"0c",	--2373
		x"0e",	--2374
		x"0f",	--2375
		x"0b",	--2376
		x"2a",	--2377
		x"0a",	--2378
		x"0b",	--2379
		x"3d",	--2380
		x"3f",	--2381
		x"00",	--2382
		x"f5",	--2383
		x"81",	--2384
		x"20",	--2385
		x"81",	--2386
		x"22",	--2387
		x"81",	--2388
		x"0a",	--2389
		x"0c",	--2390
		x"0d",	--2391
		x"3c",	--2392
		x"7f",	--2393
		x"0d",	--2394
		x"3c",	--2395
		x"40",	--2396
		x"44",	--2397
		x"81",	--2398
		x"0c",	--2399
		x"81",	--2400
		x"0e",	--2401
		x"f1",	--2402
		x"03",	--2403
		x"08",	--2404
		x"0f",	--2405
		x"3f",	--2406
		x"b0",	--2407
		x"24",	--2408
		x"31",	--2409
		x"24",	--2410
		x"34",	--2411
		x"35",	--2412
		x"36",	--2413
		x"37",	--2414
		x"38",	--2415
		x"39",	--2416
		x"3a",	--2417
		x"3b",	--2418
		x"30",	--2419
		x"1e",	--2420
		x"0f",	--2421
		x"d3",	--2422
		x"3a",	--2423
		x"03",	--2424
		x"08",	--2425
		x"1e",	--2426
		x"10",	--2427
		x"1c",	--2428
		x"20",	--2429
		x"1d",	--2430
		x"22",	--2431
		x"12",	--2432
		x"0d",	--2433
		x"0c",	--2434
		x"06",	--2435
		x"07",	--2436
		x"06",	--2437
		x"37",	--2438
		x"00",	--2439
		x"81",	--2440
		x"20",	--2441
		x"81",	--2442
		x"22",	--2443
		x"12",	--2444
		x"0f",	--2445
		x"0e",	--2446
		x"1a",	--2447
		x"0f",	--2448
		x"e7",	--2449
		x"81",	--2450
		x"0a",	--2451
		x"a6",	--2452
		x"6e",	--2453
		x"36",	--2454
		x"5f",	--2455
		x"d1",	--2456
		x"11",	--2457
		x"19",	--2458
		x"20",	--2459
		x"c1",	--2460
		x"19",	--2461
		x"0f",	--2462
		x"3f",	--2463
		x"18",	--2464
		x"c5",	--2465
		x"0d",	--2466
		x"ba",	--2467
		x"0c",	--2468
		x"0d",	--2469
		x"3c",	--2470
		x"80",	--2471
		x"0d",	--2472
		x"0c",	--2473
		x"b3",	--2474
		x"0d",	--2475
		x"b1",	--2476
		x"81",	--2477
		x"20",	--2478
		x"03",	--2479
		x"81",	--2480
		x"22",	--2481
		x"ab",	--2482
		x"3e",	--2483
		x"40",	--2484
		x"0f",	--2485
		x"3e",	--2486
		x"80",	--2487
		x"3f",	--2488
		x"a4",	--2489
		x"4d",	--2490
		x"7b",	--2491
		x"4f",	--2492
		x"de",	--2493
		x"5f",	--2494
		x"d1",	--2495
		x"11",	--2496
		x"19",	--2497
		x"06",	--2498
		x"c1",	--2499
		x"11",	--2500
		x"0f",	--2501
		x"3f",	--2502
		x"10",	--2503
		x"9e",	--2504
		x"4f",	--2505
		x"f8",	--2506
		x"6f",	--2507
		x"f1",	--2508
		x"3f",	--2509
		x"1e",	--2510
		x"97",	--2511
		x"0b",	--2512
		x"0a",	--2513
		x"09",	--2514
		x"08",	--2515
		x"07",	--2516
		x"31",	--2517
		x"e8",	--2518
		x"81",	--2519
		x"04",	--2520
		x"81",	--2521
		x"06",	--2522
		x"81",	--2523
		x"00",	--2524
		x"81",	--2525
		x"02",	--2526
		x"0e",	--2527
		x"3e",	--2528
		x"10",	--2529
		x"0f",	--2530
		x"2f",	--2531
		x"b0",	--2532
		x"02",	--2533
		x"0e",	--2534
		x"3e",	--2535
		x"0f",	--2536
		x"b0",	--2537
		x"02",	--2538
		x"5f",	--2539
		x"10",	--2540
		x"6f",	--2541
		x"5d",	--2542
		x"5e",	--2543
		x"08",	--2544
		x"6e",	--2545
		x"82",	--2546
		x"d1",	--2547
		x"09",	--2548
		x"11",	--2549
		x"6f",	--2550
		x"58",	--2551
		x"6f",	--2552
		x"56",	--2553
		x"6e",	--2554
		x"6f",	--2555
		x"6e",	--2556
		x"4c",	--2557
		x"1d",	--2558
		x"12",	--2559
		x"1d",	--2560
		x"0a",	--2561
		x"81",	--2562
		x"12",	--2563
		x"1e",	--2564
		x"14",	--2565
		x"1f",	--2566
		x"16",	--2567
		x"18",	--2568
		x"0c",	--2569
		x"19",	--2570
		x"0e",	--2571
		x"0f",	--2572
		x"1e",	--2573
		x"0e",	--2574
		x"0f",	--2575
		x"3d",	--2576
		x"81",	--2577
		x"12",	--2578
		x"37",	--2579
		x"1f",	--2580
		x"0c",	--2581
		x"3d",	--2582
		x"00",	--2583
		x"0a",	--2584
		x"0b",	--2585
		x"0b",	--2586
		x"0a",	--2587
		x"0b",	--2588
		x"0e",	--2589
		x"0f",	--2590
		x"12",	--2591
		x"0d",	--2592
		x"0c",	--2593
		x"0e",	--2594
		x"0f",	--2595
		x"37",	--2596
		x"0b",	--2597
		x"0f",	--2598
		x"f7",	--2599
		x"f2",	--2600
		x"0e",	--2601
		x"f4",	--2602
		x"ef",	--2603
		x"09",	--2604
		x"e5",	--2605
		x"0e",	--2606
		x"e3",	--2607
		x"dd",	--2608
		x"0c",	--2609
		x"0d",	--2610
		x"3c",	--2611
		x"7f",	--2612
		x"0d",	--2613
		x"3c",	--2614
		x"40",	--2615
		x"1c",	--2616
		x"81",	--2617
		x"14",	--2618
		x"81",	--2619
		x"16",	--2620
		x"0f",	--2621
		x"3f",	--2622
		x"10",	--2623
		x"b0",	--2624
		x"24",	--2625
		x"31",	--2626
		x"18",	--2627
		x"37",	--2628
		x"38",	--2629
		x"39",	--2630
		x"3a",	--2631
		x"3b",	--2632
		x"30",	--2633
		x"e1",	--2634
		x"10",	--2635
		x"0f",	--2636
		x"3f",	--2637
		x"10",	--2638
		x"f0",	--2639
		x"4f",	--2640
		x"fa",	--2641
		x"3f",	--2642
		x"1e",	--2643
		x"eb",	--2644
		x"0d",	--2645
		x"e2",	--2646
		x"0c",	--2647
		x"0d",	--2648
		x"3c",	--2649
		x"80",	--2650
		x"0d",	--2651
		x"0c",	--2652
		x"db",	--2653
		x"0d",	--2654
		x"d9",	--2655
		x"0e",	--2656
		x"02",	--2657
		x"0f",	--2658
		x"d5",	--2659
		x"3a",	--2660
		x"40",	--2661
		x"0b",	--2662
		x"3a",	--2663
		x"80",	--2664
		x"3b",	--2665
		x"ce",	--2666
		x"81",	--2667
		x"14",	--2668
		x"81",	--2669
		x"16",	--2670
		x"81",	--2671
		x"12",	--2672
		x"0f",	--2673
		x"3f",	--2674
		x"10",	--2675
		x"cb",	--2676
		x"0f",	--2677
		x"3f",	--2678
		x"c8",	--2679
		x"31",	--2680
		x"e8",	--2681
		x"81",	--2682
		x"04",	--2683
		x"81",	--2684
		x"06",	--2685
		x"81",	--2686
		x"00",	--2687
		x"81",	--2688
		x"02",	--2689
		x"0e",	--2690
		x"3e",	--2691
		x"10",	--2692
		x"0f",	--2693
		x"2f",	--2694
		x"b0",	--2695
		x"02",	--2696
		x"0e",	--2697
		x"3e",	--2698
		x"0f",	--2699
		x"b0",	--2700
		x"02",	--2701
		x"e1",	--2702
		x"10",	--2703
		x"0d",	--2704
		x"e1",	--2705
		x"08",	--2706
		x"0a",	--2707
		x"0e",	--2708
		x"3e",	--2709
		x"0f",	--2710
		x"3f",	--2711
		x"10",	--2712
		x"b0",	--2713
		x"26",	--2714
		x"31",	--2715
		x"18",	--2716
		x"30",	--2717
		x"3f",	--2718
		x"fb",	--2719
		x"31",	--2720
		x"f4",	--2721
		x"81",	--2722
		x"00",	--2723
		x"81",	--2724
		x"02",	--2725
		x"0e",	--2726
		x"2e",	--2727
		x"0f",	--2728
		x"b0",	--2729
		x"02",	--2730
		x"5f",	--2731
		x"04",	--2732
		x"6f",	--2733
		x"28",	--2734
		x"27",	--2735
		x"6f",	--2736
		x"07",	--2737
		x"1d",	--2738
		x"06",	--2739
		x"0d",	--2740
		x"21",	--2741
		x"3d",	--2742
		x"1f",	--2743
		x"09",	--2744
		x"c1",	--2745
		x"05",	--2746
		x"26",	--2747
		x"3e",	--2748
		x"3f",	--2749
		x"ff",	--2750
		x"31",	--2751
		x"0c",	--2752
		x"30",	--2753
		x"1e",	--2754
		x"08",	--2755
		x"1f",	--2756
		x"0a",	--2757
		x"3c",	--2758
		x"1e",	--2759
		x"4c",	--2760
		x"4d",	--2761
		x"7d",	--2762
		x"1f",	--2763
		x"0f",	--2764
		x"c1",	--2765
		x"05",	--2766
		x"ef",	--2767
		x"3e",	--2768
		x"3f",	--2769
		x"1e",	--2770
		x"0f",	--2771
		x"31",	--2772
		x"0c",	--2773
		x"30",	--2774
		x"0e",	--2775
		x"0f",	--2776
		x"31",	--2777
		x"0c",	--2778
		x"30",	--2779
		x"12",	--2780
		x"0f",	--2781
		x"0e",	--2782
		x"7d",	--2783
		x"fb",	--2784
		x"eb",	--2785
		x"0e",	--2786
		x"3f",	--2787
		x"00",	--2788
		x"31",	--2789
		x"0c",	--2790
		x"30",	--2791
		x"0b",	--2792
		x"0a",	--2793
		x"09",	--2794
		x"08",	--2795
		x"31",	--2796
		x"0a",	--2797
		x"0b",	--2798
		x"c1",	--2799
		x"01",	--2800
		x"0e",	--2801
		x"0d",	--2802
		x"0b",	--2803
		x"0b",	--2804
		x"e1",	--2805
		x"00",	--2806
		x"0f",	--2807
		x"b0",	--2808
		x"24",	--2809
		x"31",	--2810
		x"38",	--2811
		x"39",	--2812
		x"3a",	--2813
		x"3b",	--2814
		x"30",	--2815
		x"f1",	--2816
		x"03",	--2817
		x"00",	--2818
		x"b1",	--2819
		x"1e",	--2820
		x"02",	--2821
		x"81",	--2822
		x"04",	--2823
		x"81",	--2824
		x"06",	--2825
		x"0e",	--2826
		x"0f",	--2827
		x"b0",	--2828
		x"b2",	--2829
		x"3f",	--2830
		x"0f",	--2831
		x"18",	--2832
		x"e5",	--2833
		x"81",	--2834
		x"04",	--2835
		x"81",	--2836
		x"06",	--2837
		x"4e",	--2838
		x"7e",	--2839
		x"1f",	--2840
		x"06",	--2841
		x"3e",	--2842
		x"1e",	--2843
		x"0e",	--2844
		x"81",	--2845
		x"02",	--2846
		x"d7",	--2847
		x"91",	--2848
		x"04",	--2849
		x"04",	--2850
		x"91",	--2851
		x"06",	--2852
		x"06",	--2853
		x"7e",	--2854
		x"f8",	--2855
		x"f1",	--2856
		x"0e",	--2857
		x"3e",	--2858
		x"1e",	--2859
		x"1c",	--2860
		x"0d",	--2861
		x"48",	--2862
		x"78",	--2863
		x"1f",	--2864
		x"04",	--2865
		x"0c",	--2866
		x"0d",	--2867
		x"78",	--2868
		x"fc",	--2869
		x"3c",	--2870
		x"3d",	--2871
		x"0c",	--2872
		x"0d",	--2873
		x"18",	--2874
		x"09",	--2875
		x"0c",	--2876
		x"04",	--2877
		x"0d",	--2878
		x"02",	--2879
		x"08",	--2880
		x"09",	--2881
		x"7e",	--2882
		x"1f",	--2883
		x"0e",	--2884
		x"0d",	--2885
		x"0e",	--2886
		x"0d",	--2887
		x"0e",	--2888
		x"81",	--2889
		x"04",	--2890
		x"81",	--2891
		x"06",	--2892
		x"3e",	--2893
		x"1e",	--2894
		x"0e",	--2895
		x"81",	--2896
		x"02",	--2897
		x"a4",	--2898
		x"12",	--2899
		x"0b",	--2900
		x"0a",	--2901
		x"7e",	--2902
		x"fb",	--2903
		x"ec",	--2904
		x"0b",	--2905
		x"0a",	--2906
		x"09",	--2907
		x"1f",	--2908
		x"17",	--2909
		x"3e",	--2910
		x"00",	--2911
		x"2c",	--2912
		x"3a",	--2913
		x"18",	--2914
		x"0b",	--2915
		x"39",	--2916
		x"0c",	--2917
		x"0d",	--2918
		x"4f",	--2919
		x"4f",	--2920
		x"17",	--2921
		x"3c",	--2922
		x"26",	--2923
		x"6e",	--2924
		x"0f",	--2925
		x"0a",	--2926
		x"0b",	--2927
		x"0f",	--2928
		x"39",	--2929
		x"3a",	--2930
		x"3b",	--2931
		x"30",	--2932
		x"3f",	--2933
		x"00",	--2934
		x"0f",	--2935
		x"3a",	--2936
		x"0b",	--2937
		x"39",	--2938
		x"18",	--2939
		x"0c",	--2940
		x"0d",	--2941
		x"4f",	--2942
		x"4f",	--2943
		x"e9",	--2944
		x"12",	--2945
		x"0d",	--2946
		x"0c",	--2947
		x"7f",	--2948
		x"fb",	--2949
		x"e3",	--2950
		x"3a",	--2951
		x"10",	--2952
		x"0b",	--2953
		x"39",	--2954
		x"10",	--2955
		x"ef",	--2956
		x"3a",	--2957
		x"20",	--2958
		x"0b",	--2959
		x"09",	--2960
		x"ea",	--2961
		x"0b",	--2962
		x"0a",	--2963
		x"09",	--2964
		x"08",	--2965
		x"07",	--2966
		x"0d",	--2967
		x"1e",	--2968
		x"04",	--2969
		x"1f",	--2970
		x"06",	--2971
		x"5a",	--2972
		x"01",	--2973
		x"6c",	--2974
		x"6c",	--2975
		x"70",	--2976
		x"6c",	--2977
		x"6a",	--2978
		x"6c",	--2979
		x"36",	--2980
		x"0e",	--2981
		x"32",	--2982
		x"1b",	--2983
		x"02",	--2984
		x"3b",	--2985
		x"82",	--2986
		x"6d",	--2987
		x"3b",	--2988
		x"80",	--2989
		x"5e",	--2990
		x"0c",	--2991
		x"0d",	--2992
		x"3c",	--2993
		x"7f",	--2994
		x"0d",	--2995
		x"3c",	--2996
		x"40",	--2997
		x"40",	--2998
		x"3e",	--2999
		x"3f",	--3000
		x"0f",	--3001
		x"0f",	--3002
		x"4a",	--3003
		x"0d",	--3004
		x"3d",	--3005
		x"7f",	--3006
		x"12",	--3007
		x"0f",	--3008
		x"0e",	--3009
		x"12",	--3010
		x"0f",	--3011
		x"0e",	--3012
		x"12",	--3013
		x"0f",	--3014
		x"0e",	--3015
		x"12",	--3016
		x"0f",	--3017
		x"0e",	--3018
		x"12",	--3019
		x"0f",	--3020
		x"0e",	--3021
		x"12",	--3022
		x"0f",	--3023
		x"0e",	--3024
		x"12",	--3025
		x"0f",	--3026
		x"0e",	--3027
		x"3e",	--3028
		x"3f",	--3029
		x"7f",	--3030
		x"4d",	--3031
		x"05",	--3032
		x"0f",	--3033
		x"cc",	--3034
		x"4d",	--3035
		x"0e",	--3036
		x"0f",	--3037
		x"4d",	--3038
		x"0d",	--3039
		x"0d",	--3040
		x"0d",	--3041
		x"0d",	--3042
		x"0d",	--3043
		x"0d",	--3044
		x"0d",	--3045
		x"0c",	--3046
		x"3c",	--3047
		x"7f",	--3048
		x"0c",	--3049
		x"4f",	--3050
		x"0f",	--3051
		x"0f",	--3052
		x"0f",	--3053
		x"0d",	--3054
		x"0d",	--3055
		x"0f",	--3056
		x"37",	--3057
		x"38",	--3058
		x"39",	--3059
		x"3a",	--3060
		x"3b",	--3061
		x"30",	--3062
		x"0d",	--3063
		x"be",	--3064
		x"0c",	--3065
		x"0d",	--3066
		x"3c",	--3067
		x"80",	--3068
		x"0d",	--3069
		x"0c",	--3070
		x"02",	--3071
		x"0d",	--3072
		x"b8",	--3073
		x"3e",	--3074
		x"40",	--3075
		x"0f",	--3076
		x"b4",	--3077
		x"12",	--3078
		x"0f",	--3079
		x"0e",	--3080
		x"0d",	--3081
		x"3d",	--3082
		x"80",	--3083
		x"b2",	--3084
		x"7d",	--3085
		x"0e",	--3086
		x"0f",	--3087
		x"cd",	--3088
		x"0e",	--3089
		x"3f",	--3090
		x"10",	--3091
		x"3e",	--3092
		x"3f",	--3093
		x"7f",	--3094
		x"7d",	--3095
		x"c5",	--3096
		x"37",	--3097
		x"82",	--3098
		x"07",	--3099
		x"37",	--3100
		x"1a",	--3101
		x"4f",	--3102
		x"0c",	--3103
		x"0d",	--3104
		x"4b",	--3105
		x"7b",	--3106
		x"1f",	--3107
		x"05",	--3108
		x"12",	--3109
		x"0d",	--3110
		x"0c",	--3111
		x"7b",	--3112
		x"fb",	--3113
		x"18",	--3114
		x"09",	--3115
		x"77",	--3116
		x"1f",	--3117
		x"04",	--3118
		x"08",	--3119
		x"09",	--3120
		x"77",	--3121
		x"fc",	--3122
		x"38",	--3123
		x"39",	--3124
		x"08",	--3125
		x"09",	--3126
		x"1e",	--3127
		x"0f",	--3128
		x"08",	--3129
		x"04",	--3130
		x"09",	--3131
		x"02",	--3132
		x"0e",	--3133
		x"0f",	--3134
		x"08",	--3135
		x"09",	--3136
		x"08",	--3137
		x"09",	--3138
		x"0e",	--3139
		x"0f",	--3140
		x"3e",	--3141
		x"7f",	--3142
		x"0f",	--3143
		x"3e",	--3144
		x"40",	--3145
		x"26",	--3146
		x"38",	--3147
		x"3f",	--3148
		x"09",	--3149
		x"0e",	--3150
		x"0f",	--3151
		x"12",	--3152
		x"0f",	--3153
		x"0e",	--3154
		x"12",	--3155
		x"0f",	--3156
		x"0e",	--3157
		x"12",	--3158
		x"0f",	--3159
		x"0e",	--3160
		x"12",	--3161
		x"0f",	--3162
		x"0e",	--3163
		x"12",	--3164
		x"0f",	--3165
		x"0e",	--3166
		x"12",	--3167
		x"0f",	--3168
		x"0e",	--3169
		x"12",	--3170
		x"0f",	--3171
		x"0e",	--3172
		x"3e",	--3173
		x"3f",	--3174
		x"7f",	--3175
		x"5d",	--3176
		x"39",	--3177
		x"00",	--3178
		x"72",	--3179
		x"4d",	--3180
		x"70",	--3181
		x"08",	--3182
		x"09",	--3183
		x"da",	--3184
		x"0f",	--3185
		x"d8",	--3186
		x"0e",	--3187
		x"0f",	--3188
		x"3e",	--3189
		x"80",	--3190
		x"0f",	--3191
		x"0e",	--3192
		x"04",	--3193
		x"38",	--3194
		x"40",	--3195
		x"09",	--3196
		x"d0",	--3197
		x"0f",	--3198
		x"ce",	--3199
		x"f9",	--3200
		x"0b",	--3201
		x"0a",	--3202
		x"2a",	--3203
		x"5b",	--3204
		x"02",	--3205
		x"3b",	--3206
		x"7f",	--3207
		x"1d",	--3208
		x"02",	--3209
		x"12",	--3210
		x"0d",	--3211
		x"12",	--3212
		x"0d",	--3213
		x"12",	--3214
		x"0d",	--3215
		x"12",	--3216
		x"0d",	--3217
		x"12",	--3218
		x"0d",	--3219
		x"12",	--3220
		x"0d",	--3221
		x"12",	--3222
		x"0d",	--3223
		x"4d",	--3224
		x"5f",	--3225
		x"03",	--3226
		x"3f",	--3227
		x"80",	--3228
		x"0f",	--3229
		x"0f",	--3230
		x"ce",	--3231
		x"01",	--3232
		x"0d",	--3233
		x"2d",	--3234
		x"0a",	--3235
		x"51",	--3236
		x"be",	--3237
		x"82",	--3238
		x"02",	--3239
		x"0c",	--3240
		x"0d",	--3241
		x"0c",	--3242
		x"0d",	--3243
		x"0c",	--3244
		x"0d",	--3245
		x"0c",	--3246
		x"0d",	--3247
		x"0c",	--3248
		x"0d",	--3249
		x"0c",	--3250
		x"0d",	--3251
		x"0c",	--3252
		x"0d",	--3253
		x"0c",	--3254
		x"0d",	--3255
		x"fe",	--3256
		x"03",	--3257
		x"00",	--3258
		x"3d",	--3259
		x"00",	--3260
		x"0b",	--3261
		x"3f",	--3262
		x"81",	--3263
		x"0c",	--3264
		x"0d",	--3265
		x"0a",	--3266
		x"3f",	--3267
		x"3d",	--3268
		x"00",	--3269
		x"f9",	--3270
		x"8e",	--3271
		x"02",	--3272
		x"8e",	--3273
		x"04",	--3274
		x"8e",	--3275
		x"06",	--3276
		x"3a",	--3277
		x"3b",	--3278
		x"30",	--3279
		x"3d",	--3280
		x"ff",	--3281
		x"2a",	--3282
		x"3d",	--3283
		x"81",	--3284
		x"8e",	--3285
		x"02",	--3286
		x"fe",	--3287
		x"03",	--3288
		x"00",	--3289
		x"0c",	--3290
		x"0d",	--3291
		x"0c",	--3292
		x"0d",	--3293
		x"0c",	--3294
		x"0d",	--3295
		x"0c",	--3296
		x"0d",	--3297
		x"0c",	--3298
		x"0d",	--3299
		x"0c",	--3300
		x"0d",	--3301
		x"0c",	--3302
		x"0d",	--3303
		x"0c",	--3304
		x"0d",	--3305
		x"0a",	--3306
		x"0b",	--3307
		x"0a",	--3308
		x"3b",	--3309
		x"00",	--3310
		x"8e",	--3311
		x"04",	--3312
		x"8e",	--3313
		x"06",	--3314
		x"3a",	--3315
		x"3b",	--3316
		x"30",	--3317
		x"0b",	--3318
		x"ad",	--3319
		x"ee",	--3320
		x"00",	--3321
		x"3a",	--3322
		x"3b",	--3323
		x"30",	--3324
		x"0a",	--3325
		x"0c",	--3326
		x"0c",	--3327
		x"0d",	--3328
		x"0c",	--3329
		x"3d",	--3330
		x"10",	--3331
		x"0c",	--3332
		x"02",	--3333
		x"0d",	--3334
		x"08",	--3335
		x"de",	--3336
		x"00",	--3337
		x"e4",	--3338
		x"0b",	--3339
		x"f2",	--3340
		x"ee",	--3341
		x"00",	--3342
		x"e3",	--3343
		x"ce",	--3344
		x"00",	--3345
		x"dc",	--3346
		x"0b",	--3347
		x"6d",	--3348
		x"6d",	--3349
		x"12",	--3350
		x"6c",	--3351
		x"6c",	--3352
		x"0f",	--3353
		x"6d",	--3354
		x"41",	--3355
		x"6c",	--3356
		x"11",	--3357
		x"6d",	--3358
		x"0d",	--3359
		x"6c",	--3360
		x"14",	--3361
		x"5d",	--3362
		x"01",	--3363
		x"5d",	--3364
		x"01",	--3365
		x"14",	--3366
		x"4d",	--3367
		x"09",	--3368
		x"1e",	--3369
		x"0f",	--3370
		x"3b",	--3371
		x"30",	--3372
		x"6c",	--3373
		x"28",	--3374
		x"ce",	--3375
		x"01",	--3376
		x"f7",	--3377
		x"3e",	--3378
		x"0f",	--3379
		x"3b",	--3380
		x"30",	--3381
		x"cf",	--3382
		x"01",	--3383
		x"f0",	--3384
		x"3e",	--3385
		x"f8",	--3386
		x"1b",	--3387
		x"02",	--3388
		x"1c",	--3389
		x"02",	--3390
		x"0c",	--3391
		x"e6",	--3392
		x"0b",	--3393
		x"16",	--3394
		x"1b",	--3395
		x"04",	--3396
		x"1f",	--3397
		x"06",	--3398
		x"1c",	--3399
		x"04",	--3400
		x"1e",	--3401
		x"06",	--3402
		x"0e",	--3403
		x"da",	--3404
		x"0f",	--3405
		x"02",	--3406
		x"0c",	--3407
		x"d6",	--3408
		x"0f",	--3409
		x"06",	--3410
		x"0e",	--3411
		x"02",	--3412
		x"0b",	--3413
		x"02",	--3414
		x"0e",	--3415
		x"d1",	--3416
		x"4d",	--3417
		x"ce",	--3418
		x"3e",	--3419
		x"d6",	--3420
		x"6c",	--3421
		x"d7",	--3422
		x"5e",	--3423
		x"01",	--3424
		x"5f",	--3425
		x"01",	--3426
		x"0e",	--3427
		x"c5",	--3428
		x"1e",	--3429
		x"1a",	--3430
		x"1e",	--3431
		x"0b",	--3432
		x"1d",	--3433
		x"18",	--3434
		x"cd",	--3435
		x"00",	--3436
		x"1d",	--3437
		x"82",	--3438
		x"18",	--3439
		x"3e",	--3440
		x"82",	--3441
		x"1a",	--3442
		x"30",	--3443
		x"3f",	--3444
		x"30",	--3445
		x"0b",	--3446
		x"0a",	--3447
		x"21",	--3448
		x"81",	--3449
		x"00",	--3450
		x"1a",	--3451
		x"18",	--3452
		x"1b",	--3453
		x"1a",	--3454
		x"0d",	--3455
		x"0e",	--3456
		x"3f",	--3457
		x"ca",	--3458
		x"b0",	--3459
		x"1e",	--3460
		x"0f",	--3461
		x"05",	--3462
		x"0e",	--3463
		x"0e",	--3464
		x"ce",	--3465
		x"ff",	--3466
		x"04",	--3467
		x"1e",	--3468
		x"18",	--3469
		x"ce",	--3470
		x"00",	--3471
		x"21",	--3472
		x"3a",	--3473
		x"3b",	--3474
		x"30",	--3475
		x"92",	--3476
		x"02",	--3477
		x"18",	--3478
		x"b2",	--3479
		x"ff",	--3480
		x"1a",	--3481
		x"0e",	--3482
		x"3e",	--3483
		x"06",	--3484
		x"1f",	--3485
		x"04",	--3486
		x"b0",	--3487
		x"ec",	--3488
		x"30",	--3489
		x"92",	--3490
		x"02",	--3491
		x"18",	--3492
		x"92",	--3493
		x"04",	--3494
		x"1a",	--3495
		x"0e",	--3496
		x"3e",	--3497
		x"1f",	--3498
		x"06",	--3499
		x"b0",	--3500
		x"ec",	--3501
		x"30",	--3502
		x"0c",	--3503
		x"82",	--3504
		x"18",	--3505
		x"b2",	--3506
		x"ff",	--3507
		x"1a",	--3508
		x"0e",	--3509
		x"0f",	--3510
		x"b0",	--3511
		x"ec",	--3512
		x"30",	--3513
		x"82",	--3514
		x"18",	--3515
		x"82",	--3516
		x"1a",	--3517
		x"0e",	--3518
		x"0f",	--3519
		x"b0",	--3520
		x"ec",	--3521
		x"30",	--3522
		x"0b",	--3523
		x"0a",	--3524
		x"09",	--3525
		x"08",	--3526
		x"07",	--3527
		x"06",	--3528
		x"05",	--3529
		x"04",	--3530
		x"31",	--3531
		x"08",	--3532
		x"81",	--3533
		x"04",	--3534
		x"09",	--3535
		x"1f",	--3536
		x"1a",	--3537
		x"1d",	--3538
		x"1c",	--3539
		x"4c",	--3540
		x"04",	--3541
		x"84",	--3542
		x"45",	--3543
		x"4e",	--3544
		x"7e",	--3545
		x"40",	--3546
		x"11",	--3547
		x"f1",	--3548
		x"30",	--3549
		x"00",	--3550
		x"0e",	--3551
		x"8e",	--3552
		x"5e",	--3553
		x"03",	--3554
		x"7e",	--3555
		x"58",	--3556
		x"02",	--3557
		x"7e",	--3558
		x"78",	--3559
		x"c1",	--3560
		x"01",	--3561
		x"0c",	--3562
		x"2c",	--3563
		x"0f",	--3564
		x"7e",	--3565
		x"20",	--3566
		x"04",	--3567
		x"f1",	--3568
		x"30",	--3569
		x"00",	--3570
		x"04",	--3571
		x"4c",	--3572
		x"05",	--3573
		x"c1",	--3574
		x"00",	--3575
		x"0c",	--3576
		x"1c",	--3577
		x"01",	--3578
		x"0c",	--3579
		x"0a",	--3580
		x"8c",	--3581
		x"8c",	--3582
		x"8c",	--3583
		x"8c",	--3584
		x"0b",	--3585
		x"06",	--3586
		x"0c",	--3587
		x"8c",	--3588
		x"8c",	--3589
		x"8c",	--3590
		x"8c",	--3591
		x"07",	--3592
		x"0a",	--3593
		x"0b",	--3594
		x"0e",	--3595
		x"8e",	--3596
		x"c1",	--3597
		x"02",	--3598
		x"6e",	--3599
		x"02",	--3600
		x"07",	--3601
		x"01",	--3602
		x"37",	--3603
		x"4f",	--3604
		x"7f",	--3605
		x"10",	--3606
		x"3c",	--3607
		x"1d",	--3608
		x"04",	--3609
		x"3d",	--3610
		x"1d",	--3611
		x"cd",	--3612
		x"00",	--3613
		x"fc",	--3614
		x"1d",	--3615
		x"04",	--3616
		x"09",	--3617
		x"02",	--3618
		x"09",	--3619
		x"01",	--3620
		x"09",	--3621
		x"e1",	--3622
		x"02",	--3623
		x"05",	--3624
		x"09",	--3625
		x"02",	--3626
		x"09",	--3627
		x"01",	--3628
		x"09",	--3629
		x"05",	--3630
		x"07",	--3631
		x"01",	--3632
		x"05",	--3633
		x"4f",	--3634
		x"0d",	--3635
		x"f1",	--3636
		x"20",	--3637
		x"06",	--3638
		x"06",	--3639
		x"0b",	--3640
		x"0e",	--3641
		x"0f",	--3642
		x"0f",	--3643
		x"6f",	--3644
		x"8f",	--3645
		x"16",	--3646
		x"88",	--3647
		x"01",	--3648
		x"06",	--3649
		x"06",	--3650
		x"f6",	--3651
		x"0b",	--3652
		x"f1",	--3653
		x"30",	--3654
		x"06",	--3655
		x"05",	--3656
		x"05",	--3657
		x"5f",	--3658
		x"06",	--3659
		x"8f",	--3660
		x"88",	--3661
		x"1b",	--3662
		x"0f",	--3663
		x"0f",	--3664
		x"0f",	--3665
		x"f7",	--3666
		x"0a",	--3667
		x"06",	--3668
		x"0b",	--3669
		x"07",	--3670
		x"1b",	--3671
		x"0f",	--3672
		x"0f",	--3673
		x"6f",	--3674
		x"8f",	--3675
		x"16",	--3676
		x"88",	--3677
		x"06",	--3678
		x"f7",	--3679
		x"e1",	--3680
		x"02",	--3681
		x"02",	--3682
		x"4a",	--3683
		x"08",	--3684
		x"1a",	--3685
		x"04",	--3686
		x"0a",	--3687
		x"0d",	--3688
		x"3f",	--3689
		x"30",	--3690
		x"88",	--3691
		x"7a",	--3692
		x"4a",	--3693
		x"fa",	--3694
		x"44",	--3695
		x"0b",	--3696
		x"f3",	--3697
		x"37",	--3698
		x"8f",	--3699
		x"88",	--3700
		x"1b",	--3701
		x"0f",	--3702
		x"0f",	--3703
		x"6f",	--3704
		x"4f",	--3705
		x"07",	--3706
		x"07",	--3707
		x"f5",	--3708
		x"04",	--3709
		x"3f",	--3710
		x"20",	--3711
		x"88",	--3712
		x"1b",	--3713
		x"0b",	--3714
		x"fa",	--3715
		x"0f",	--3716
		x"31",	--3717
		x"34",	--3718
		x"35",	--3719
		x"36",	--3720
		x"37",	--3721
		x"38",	--3722
		x"39",	--3723
		x"3a",	--3724
		x"3b",	--3725
		x"30",	--3726
		x"0b",	--3727
		x"0a",	--3728
		x"09",	--3729
		x"08",	--3730
		x"07",	--3731
		x"06",	--3732
		x"05",	--3733
		x"04",	--3734
		x"31",	--3735
		x"b6",	--3736
		x"81",	--3737
		x"3a",	--3738
		x"06",	--3739
		x"05",	--3740
		x"81",	--3741
		x"3e",	--3742
		x"c1",	--3743
		x"2f",	--3744
		x"c1",	--3745
		x"2b",	--3746
		x"c1",	--3747
		x"2e",	--3748
		x"c1",	--3749
		x"2a",	--3750
		x"81",	--3751
		x"30",	--3752
		x"81",	--3753
		x"26",	--3754
		x"07",	--3755
		x"81",	--3756
		x"2c",	--3757
		x"0e",	--3758
		x"3e",	--3759
		x"1c",	--3760
		x"81",	--3761
		x"1c",	--3762
		x"30",	--3763
		x"98",	--3764
		x"0f",	--3765
		x"1f",	--3766
		x"81",	--3767
		x"40",	--3768
		x"07",	--3769
		x"1e",	--3770
		x"7e",	--3771
		x"25",	--3772
		x"13",	--3773
		x"81",	--3774
		x"00",	--3775
		x"81",	--3776
		x"02",	--3777
		x"81",	--3778
		x"3e",	--3779
		x"c1",	--3780
		x"2f",	--3781
		x"c1",	--3782
		x"2b",	--3783
		x"c1",	--3784
		x"2e",	--3785
		x"c1",	--3786
		x"2a",	--3787
		x"81",	--3788
		x"30",	--3789
		x"30",	--3790
		x"8e",	--3791
		x"05",	--3792
		x"8e",	--3793
		x"0f",	--3794
		x"91",	--3795
		x"3c",	--3796
		x"91",	--3797
		x"2c",	--3798
		x"30",	--3799
		x"74",	--3800
		x"7e",	--3801
		x"63",	--3802
		x"c5",	--3803
		x"7e",	--3804
		x"64",	--3805
		x"27",	--3806
		x"7e",	--3807
		x"30",	--3808
		x"94",	--3809
		x"7e",	--3810
		x"31",	--3811
		x"1a",	--3812
		x"7e",	--3813
		x"2a",	--3814
		x"77",	--3815
		x"7e",	--3816
		x"2b",	--3817
		x"0a",	--3818
		x"7e",	--3819
		x"23",	--3820
		x"42",	--3821
		x"7e",	--3822
		x"25",	--3823
		x"e0",	--3824
		x"7e",	--3825
		x"20",	--3826
		x"32",	--3827
		x"56",	--3828
		x"7e",	--3829
		x"2d",	--3830
		x"49",	--3831
		x"7e",	--3832
		x"2e",	--3833
		x"5b",	--3834
		x"7e",	--3835
		x"2b",	--3836
		x"28",	--3837
		x"47",	--3838
		x"7e",	--3839
		x"3a",	--3840
		x"8c",	--3841
		x"7e",	--3842
		x"58",	--3843
		x"21",	--3844
		x"e9",	--3845
		x"7e",	--3846
		x"6f",	--3847
		x"24",	--3848
		x"7e",	--3849
		x"70",	--3850
		x"0a",	--3851
		x"7e",	--3852
		x"69",	--3853
		x"e3",	--3854
		x"7e",	--3855
		x"6c",	--3856
		x"22",	--3857
		x"7e",	--3858
		x"64",	--3859
		x"11",	--3860
		x"dc",	--3861
		x"7e",	--3862
		x"73",	--3863
		x"98",	--3864
		x"7e",	--3865
		x"74",	--3866
		x"04",	--3867
		x"7e",	--3868
		x"70",	--3869
		x"07",	--3870
		x"b8",	--3871
		x"7e",	--3872
		x"75",	--3873
		x"d1",	--3874
		x"7e",	--3875
		x"78",	--3876
		x"d2",	--3877
		x"19",	--3878
		x"3e",	--3879
		x"18",	--3880
		x"2c",	--3881
		x"08",	--3882
		x"30",	--3883
		x"62",	--3884
		x"b1",	--3885
		x"28",	--3886
		x"cb",	--3887
		x"f1",	--3888
		x"00",	--3889
		x"30",	--3890
		x"92",	--3891
		x"69",	--3892
		x"59",	--3893
		x"6e",	--3894
		x"04",	--3895
		x"7e",	--3896
		x"fe",	--3897
		x"6e",	--3898
		x"01",	--3899
		x"5e",	--3900
		x"c1",	--3901
		x"00",	--3902
		x"30",	--3903
		x"92",	--3904
		x"f1",	--3905
		x"10",	--3906
		x"00",	--3907
		x"30",	--3908
		x"92",	--3909
		x"f1",	--3910
		x"2b",	--3911
		x"02",	--3912
		x"30",	--3913
		x"92",	--3914
		x"f1",	--3915
		x"2b",	--3916
		x"02",	--3917
		x"02",	--3918
		x"30",	--3919
		x"92",	--3920
		x"f1",	--3921
		x"20",	--3922
		x"02",	--3923
		x"30",	--3924
		x"92",	--3925
		x"c1",	--3926
		x"2a",	--3927
		x"02",	--3928
		x"30",	--3929
		x"78",	--3930
		x"d1",	--3931
		x"2e",	--3932
		x"30",	--3933
		x"92",	--3934
		x"0e",	--3935
		x"2e",	--3936
		x"2a",	--3937
		x"0a",	--3938
		x"03",	--3939
		x"81",	--3940
		x"26",	--3941
		x"0d",	--3942
		x"c1",	--3943
		x"2e",	--3944
		x"02",	--3945
		x"30",	--3946
		x"88",	--3947
		x"f1",	--3948
		x"10",	--3949
		x"00",	--3950
		x"3a",	--3951
		x"81",	--3952
		x"26",	--3953
		x"91",	--3954
		x"26",	--3955
		x"05",	--3956
		x"27",	--3957
		x"81",	--3958
		x"26",	--3959
		x"15",	--3960
		x"c1",	--3961
		x"2e",	--3962
		x"12",	--3963
		x"69",	--3964
		x"79",	--3965
		x"10",	--3966
		x"5e",	--3967
		x"01",	--3968
		x"4e",	--3969
		x"4e",	--3970
		x"0e",	--3971
		x"0e",	--3972
		x"4e",	--3973
		x"6a",	--3974
		x"7a",	--3975
		x"7f",	--3976
		x"4a",	--3977
		x"c1",	--3978
		x"00",	--3979
		x"30",	--3980
		x"92",	--3981
		x"1a",	--3982
		x"26",	--3983
		x"0a",	--3984
		x"0c",	--3985
		x"0c",	--3986
		x"0c",	--3987
		x"0a",	--3988
		x"81",	--3989
		x"26",	--3990
		x"b1",	--3991
		x"d0",	--3992
		x"26",	--3993
		x"8e",	--3994
		x"81",	--3995
		x"26",	--3996
		x"d1",	--3997
		x"2a",	--3998
		x"30",	--3999
		x"92",	--4000
		x"07",	--4001
		x"27",	--4002
		x"6e",	--4003
		x"c1",	--4004
		x"2e",	--4005
		x"03",	--4006
		x"c1",	--4007
		x"2a",	--4008
		x"26",	--4009
		x"c1",	--4010
		x"04",	--4011
		x"c1",	--4012
		x"05",	--4013
		x"0e",	--4014
		x"2e",	--4015
		x"03",	--4016
		x"07",	--4017
		x"27",	--4018
		x"2e",	--4019
		x"c1",	--4020
		x"2e",	--4021
		x"07",	--4022
		x"e1",	--4023
		x"01",	--4024
		x"1f",	--4025
		x"26",	--4026
		x"c1",	--4027
		x"03",	--4028
		x"06",	--4029
		x"c1",	--4030
		x"2a",	--4031
		x"03",	--4032
		x"91",	--4033
		x"26",	--4034
		x"30",	--4035
		x"0e",	--4036
		x"02",	--4037
		x"3e",	--4038
		x"26",	--4039
		x"11",	--4040
		x"04",	--4041
		x"11",	--4042
		x"04",	--4043
		x"1d",	--4044
		x"34",	--4045
		x"1f",	--4046
		x"3e",	--4047
		x"b0",	--4048
		x"86",	--4049
		x"21",	--4050
		x"81",	--4051
		x"2c",	--4052
		x"05",	--4053
		x"30",	--4054
		x"74",	--4055
		x"07",	--4056
		x"27",	--4057
		x"29",	--4058
		x"81",	--4059
		x"1e",	--4060
		x"5e",	--4061
		x"09",	--4062
		x"01",	--4063
		x"4e",	--4064
		x"4e",	--4065
		x"4e",	--4066
		x"4e",	--4067
		x"6a",	--4068
		x"7a",	--4069
		x"f7",	--4070
		x"4a",	--4071
		x"c1",	--4072
		x"00",	--4073
		x"05",	--4074
		x"b1",	--4075
		x"10",	--4076
		x"28",	--4077
		x"53",	--4078
		x"d1",	--4079
		x"01",	--4080
		x"06",	--4081
		x"e1",	--4082
		x"00",	--4083
		x"b1",	--4084
		x"0a",	--4085
		x"28",	--4086
		x"03",	--4087
		x"b1",	--4088
		x"10",	--4089
		x"28",	--4090
		x"6b",	--4091
		x"6b",	--4092
		x"24",	--4093
		x"0c",	--4094
		x"3c",	--4095
		x"28",	--4096
		x"17",	--4097
		x"02",	--4098
		x"16",	--4099
		x"04",	--4100
		x"1b",	--4101
		x"06",	--4102
		x"81",	--4103
		x"1e",	--4104
		x"81",	--4105
		x"20",	--4106
		x"81",	--4107
		x"22",	--4108
		x"81",	--4109
		x"24",	--4110
		x"d1",	--4111
		x"2b",	--4112
		x"08",	--4113
		x"06",	--4114
		x"07",	--4115
		x"04",	--4116
		x"06",	--4117
		x"02",	--4118
		x"0b",	--4119
		x"02",	--4120
		x"c1",	--4121
		x"2b",	--4122
		x"0b",	--4123
		x"0b",	--4124
		x"0b",	--4125
		x"c1",	--4126
		x"2f",	--4127
		x"05",	--4128
		x"20",	--4129
		x"5b",	--4130
		x"07",	--4131
		x"0d",	--4132
		x"27",	--4133
		x"28",	--4134
		x"1b",	--4135
		x"02",	--4136
		x"81",	--4137
		x"1e",	--4138
		x"81",	--4139
		x"20",	--4140
		x"d1",	--4141
		x"2b",	--4142
		x"08",	--4143
		x"09",	--4144
		x"06",	--4145
		x"27",	--4146
		x"2b",	--4147
		x"81",	--4148
		x"1e",	--4149
		x"d1",	--4150
		x"2b",	--4151
		x"0b",	--4152
		x"02",	--4153
		x"c1",	--4154
		x"2b",	--4155
		x"0b",	--4156
		x"0b",	--4157
		x"0b",	--4158
		x"c1",	--4159
		x"2f",	--4160
		x"05",	--4161
		x"f1",	--4162
		x"00",	--4163
		x"12",	--4164
		x"c1",	--4165
		x"2b",	--4166
		x"0f",	--4167
		x"68",	--4168
		x"b1",	--4169
		x"10",	--4170
		x"28",	--4171
		x"03",	--4172
		x"78",	--4173
		x"40",	--4174
		x"05",	--4175
		x"b1",	--4176
		x"28",	--4177
		x"04",	--4178
		x"78",	--4179
		x"20",	--4180
		x"c1",	--4181
		x"00",	--4182
		x"68",	--4183
		x"68",	--4184
		x"30",	--4185
		x"c1",	--4186
		x"2f",	--4187
		x"2d",	--4188
		x"f1",	--4189
		x"2d",	--4190
		x"02",	--4191
		x"68",	--4192
		x"11",	--4193
		x"b1",	--4194
		x"1e",	--4195
		x"b1",	--4196
		x"20",	--4197
		x"b1",	--4198
		x"22",	--4199
		x"b1",	--4200
		x"24",	--4201
		x"91",	--4202
		x"1e",	--4203
		x"81",	--4204
		x"20",	--4205
		x"81",	--4206
		x"22",	--4207
		x"81",	--4208
		x"24",	--4209
		x"17",	--4210
		x"58",	--4211
		x"0f",	--4212
		x"1a",	--4213
		x"1e",	--4214
		x"1b",	--4215
		x"20",	--4216
		x"3a",	--4217
		x"3b",	--4218
		x"0e",	--4219
		x"0f",	--4220
		x"1e",	--4221
		x"0f",	--4222
		x"81",	--4223
		x"1e",	--4224
		x"81",	--4225
		x"20",	--4226
		x"06",	--4227
		x"1a",	--4228
		x"1e",	--4229
		x"3a",	--4230
		x"1a",	--4231
		x"81",	--4232
		x"1e",	--4233
		x"c1",	--4234
		x"1b",	--4235
		x"68",	--4236
		x"6a",	--4237
		x"16",	--4238
		x"1e",	--4239
		x"91",	--4240
		x"20",	--4241
		x"3c",	--4242
		x"18",	--4243
		x"22",	--4244
		x"14",	--4245
		x"24",	--4246
		x"07",	--4247
		x"37",	--4248
		x"1a",	--4249
		x"09",	--4250
		x"91",	--4251
		x"28",	--4252
		x"32",	--4253
		x"1b",	--4254
		x"28",	--4255
		x"8b",	--4256
		x"8b",	--4257
		x"8b",	--4258
		x"8b",	--4259
		x"81",	--4260
		x"34",	--4261
		x"81",	--4262
		x"36",	--4263
		x"81",	--4264
		x"38",	--4265
		x"11",	--4266
		x"3a",	--4267
		x"11",	--4268
		x"3a",	--4269
		x"11",	--4270
		x"3a",	--4271
		x"11",	--4272
		x"3a",	--4273
		x"0c",	--4274
		x"1d",	--4275
		x"44",	--4276
		x"0e",	--4277
		x"0f",	--4278
		x"b0",	--4279
		x"28",	--4280
		x"31",	--4281
		x"0b",	--4282
		x"3c",	--4283
		x"0a",	--4284
		x"05",	--4285
		x"7b",	--4286
		x"30",	--4287
		x"c7",	--4288
		x"00",	--4289
		x"0c",	--4290
		x"4b",	--4291
		x"d1",	--4292
		x"01",	--4293
		x"03",	--4294
		x"7a",	--4295
		x"37",	--4296
		x"02",	--4297
		x"7a",	--4298
		x"57",	--4299
		x"4a",	--4300
		x"c7",	--4301
		x"00",	--4302
		x"06",	--4303
		x"36",	--4304
		x"11",	--4305
		x"3a",	--4306
		x"11",	--4307
		x"3a",	--4308
		x"11",	--4309
		x"3a",	--4310
		x"11",	--4311
		x"3a",	--4312
		x"0c",	--4313
		x"1d",	--4314
		x"44",	--4315
		x"0e",	--4316
		x"0f",	--4317
		x"b0",	--4318
		x"02",	--4319
		x"31",	--4320
		x"09",	--4321
		x"81",	--4322
		x"3c",	--4323
		x"08",	--4324
		x"04",	--4325
		x"37",	--4326
		x"0c",	--4327
		x"b2",	--4328
		x"0d",	--4329
		x"b0",	--4330
		x"0e",	--4331
		x"ae",	--4332
		x"0f",	--4333
		x"ac",	--4334
		x"81",	--4335
		x"1e",	--4336
		x"81",	--4337
		x"20",	--4338
		x"81",	--4339
		x"22",	--4340
		x"81",	--4341
		x"24",	--4342
		x"6c",	--4343
		x"58",	--4344
		x"3e",	--4345
		x"14",	--4346
		x"1e",	--4347
		x"17",	--4348
		x"20",	--4349
		x"08",	--4350
		x"38",	--4351
		x"1a",	--4352
		x"19",	--4353
		x"28",	--4354
		x"89",	--4355
		x"89",	--4356
		x"89",	--4357
		x"89",	--4358
		x"1c",	--4359
		x"28",	--4360
		x"0d",	--4361
		x"0e",	--4362
		x"0f",	--4363
		x"b0",	--4364
		x"2c",	--4365
		x"0b",	--4366
		x"3e",	--4367
		x"0a",	--4368
		x"05",	--4369
		x"7b",	--4370
		x"30",	--4371
		x"c8",	--4372
		x"00",	--4373
		x"0c",	--4374
		x"4b",	--4375
		x"d1",	--4376
		x"01",	--4377
		x"03",	--4378
		x"7a",	--4379
		x"37",	--4380
		x"02",	--4381
		x"7a",	--4382
		x"57",	--4383
		x"4a",	--4384
		x"c8",	--4385
		x"00",	--4386
		x"06",	--4387
		x"36",	--4388
		x"1c",	--4389
		x"28",	--4390
		x"0d",	--4391
		x"0e",	--4392
		x"0f",	--4393
		x"b0",	--4394
		x"f6",	--4395
		x"04",	--4396
		x"07",	--4397
		x"38",	--4398
		x"0e",	--4399
		x"d0",	--4400
		x"0f",	--4401
		x"ce",	--4402
		x"81",	--4403
		x"1e",	--4404
		x"81",	--4405
		x"20",	--4406
		x"2c",	--4407
		x"17",	--4408
		x"1e",	--4409
		x"08",	--4410
		x"38",	--4411
		x"1a",	--4412
		x"1e",	--4413
		x"28",	--4414
		x"0f",	--4415
		x"b0",	--4416
		x"9c",	--4417
		x"0d",	--4418
		x"3f",	--4419
		x"0a",	--4420
		x"05",	--4421
		x"7d",	--4422
		x"30",	--4423
		x"c8",	--4424
		x"00",	--4425
		x"0c",	--4426
		x"4d",	--4427
		x"d1",	--4428
		x"01",	--4429
		x"03",	--4430
		x"7c",	--4431
		x"37",	--4432
		x"02",	--4433
		x"7c",	--4434
		x"57",	--4435
		x"4c",	--4436
		x"c8",	--4437
		x"00",	--4438
		x"06",	--4439
		x"36",	--4440
		x"1e",	--4441
		x"28",	--4442
		x"0f",	--4443
		x"b0",	--4444
		x"82",	--4445
		x"07",	--4446
		x"38",	--4447
		x"0f",	--4448
		x"db",	--4449
		x"81",	--4450
		x"1e",	--4451
		x"b1",	--4452
		x"0a",	--4453
		x"28",	--4454
		x"02",	--4455
		x"c1",	--4456
		x"02",	--4457
		x"c1",	--4458
		x"2e",	--4459
		x"2a",	--4460
		x"0f",	--4461
		x"3f",	--4462
		x"1c",	--4463
		x"81",	--4464
		x"42",	--4465
		x"1a",	--4466
		x"1c",	--4467
		x"8a",	--4468
		x"8a",	--4469
		x"8a",	--4470
		x"8a",	--4471
		x"81",	--4472
		x"44",	--4473
		x"81",	--4474
		x"46",	--4475
		x"0a",	--4476
		x"8a",	--4477
		x"8a",	--4478
		x"8a",	--4479
		x"8a",	--4480
		x"81",	--4481
		x"48",	--4482
		x"1c",	--4483
		x"42",	--4484
		x"1d",	--4485
		x"44",	--4486
		x"1c",	--4487
		x"46",	--4488
		x"1d",	--4489
		x"48",	--4490
		x"2c",	--4491
		x"1c",	--4492
		x"26",	--4493
		x"0e",	--4494
		x"e1",	--4495
		x"01",	--4496
		x"5e",	--4497
		x"26",	--4498
		x"4e",	--4499
		x"c1",	--4500
		x"03",	--4501
		x"06",	--4502
		x"c1",	--4503
		x"2a",	--4504
		x"03",	--4505
		x"91",	--4506
		x"26",	--4507
		x"30",	--4508
		x"11",	--4509
		x"04",	--4510
		x"11",	--4511
		x"04",	--4512
		x"1d",	--4513
		x"34",	--4514
		x"0e",	--4515
		x"1e",	--4516
		x"1f",	--4517
		x"3e",	--4518
		x"b0",	--4519
		x"86",	--4520
		x"21",	--4521
		x"81",	--4522
		x"2c",	--4523
		x"0d",	--4524
		x"7f",	--4525
		x"8f",	--4526
		x"91",	--4527
		x"3c",	--4528
		x"0e",	--4529
		x"0e",	--4530
		x"19",	--4531
		x"40",	--4532
		x"f7",	--4533
		x"81",	--4534
		x"3e",	--4535
		x"81",	--4536
		x"2c",	--4537
		x"07",	--4538
		x"0e",	--4539
		x"91",	--4540
		x"26",	--4541
		x"30",	--4542
		x"d1",	--4543
		x"2e",	--4544
		x"c1",	--4545
		x"2a",	--4546
		x"03",	--4547
		x"05",	--4548
		x"d1",	--4549
		x"2a",	--4550
		x"81",	--4551
		x"26",	--4552
		x"17",	--4553
		x"16",	--4554
		x"40",	--4555
		x"6e",	--4556
		x"4e",	--4557
		x"02",	--4558
		x"30",	--4559
		x"6a",	--4560
		x"1f",	--4561
		x"2c",	--4562
		x"31",	--4563
		x"4a",	--4564
		x"34",	--4565
		x"35",	--4566
		x"36",	--4567
		x"37",	--4568
		x"38",	--4569
		x"39",	--4570
		x"3a",	--4571
		x"3b",	--4572
		x"30",	--4573
		x"0d",	--4574
		x"0f",	--4575
		x"04",	--4576
		x"3d",	--4577
		x"03",	--4578
		x"3f",	--4579
		x"1f",	--4580
		x"0e",	--4581
		x"03",	--4582
		x"5d",	--4583
		x"3e",	--4584
		x"1e",	--4585
		x"0d",	--4586
		x"b0",	--4587
		x"82",	--4588
		x"3d",	--4589
		x"6d",	--4590
		x"02",	--4591
		x"3e",	--4592
		x"1e",	--4593
		x"5d",	--4594
		x"02",	--4595
		x"3f",	--4596
		x"1f",	--4597
		x"30",	--4598
		x"b0",	--4599
		x"bc",	--4600
		x"0f",	--4601
		x"30",	--4602
		x"0b",	--4603
		x"0a",	--4604
		x"09",	--4605
		x"79",	--4606
		x"20",	--4607
		x"0a",	--4608
		x"0b",	--4609
		x"0c",	--4610
		x"0d",	--4611
		x"0e",	--4612
		x"0f",	--4613
		x"0c",	--4614
		x"0d",	--4615
		x"0d",	--4616
		x"06",	--4617
		x"02",	--4618
		x"0c",	--4619
		x"03",	--4620
		x"0c",	--4621
		x"0d",	--4622
		x"1e",	--4623
		x"19",	--4624
		x"f2",	--4625
		x"39",	--4626
		x"3a",	--4627
		x"3b",	--4628
		x"30",	--4629
		x"b0",	--4630
		x"f6",	--4631
		x"0e",	--4632
		x"0f",	--4633
		x"30",	--4634
		x"0b",	--4635
		x"0b",	--4636
		x"0f",	--4637
		x"06",	--4638
		x"3b",	--4639
		x"03",	--4640
		x"3e",	--4641
		x"3f",	--4642
		x"1e",	--4643
		x"0f",	--4644
		x"0d",	--4645
		x"05",	--4646
		x"5b",	--4647
		x"3c",	--4648
		x"3d",	--4649
		x"1c",	--4650
		x"0d",	--4651
		x"b0",	--4652
		x"f6",	--4653
		x"6b",	--4654
		x"04",	--4655
		x"3c",	--4656
		x"3d",	--4657
		x"1c",	--4658
		x"0d",	--4659
		x"5b",	--4660
		x"04",	--4661
		x"3e",	--4662
		x"3f",	--4663
		x"1e",	--4664
		x"0f",	--4665
		x"3b",	--4666
		x"30",	--4667
		x"b0",	--4668
		x"36",	--4669
		x"0e",	--4670
		x"0f",	--4671
		x"30",	--4672
		x"7c",	--4673
		x"10",	--4674
		x"0d",	--4675
		x"0e",	--4676
		x"0f",	--4677
		x"0e",	--4678
		x"0e",	--4679
		x"02",	--4680
		x"0e",	--4681
		x"1f",	--4682
		x"1c",	--4683
		x"f8",	--4684
		x"30",	--4685
		x"b0",	--4686
		x"82",	--4687
		x"0f",	--4688
		x"30",	--4689
		x"07",	--4690
		x"06",	--4691
		x"05",	--4692
		x"04",	--4693
		x"30",	--4694
		x"40",	--4695
		x"04",	--4696
		x"05",	--4697
		x"06",	--4698
		x"07",	--4699
		x"08",	--4700
		x"09",	--4701
		x"0a",	--4702
		x"0b",	--4703
		x"0c",	--4704
		x"0d",	--4705
		x"0e",	--4706
		x"0f",	--4707
		x"08",	--4708
		x"09",	--4709
		x"0a",	--4710
		x"0b",	--4711
		x"0b",	--4712
		x"0e",	--4713
		x"08",	--4714
		x"0a",	--4715
		x"0b",	--4716
		x"05",	--4717
		x"09",	--4718
		x"08",	--4719
		x"02",	--4720
		x"08",	--4721
		x"05",	--4722
		x"08",	--4723
		x"09",	--4724
		x"0a",	--4725
		x"0b",	--4726
		x"1c",	--4727
		x"91",	--4728
		x"00",	--4729
		x"e5",	--4730
		x"21",	--4731
		x"34",	--4732
		x"35",	--4733
		x"36",	--4734
		x"37",	--4735
		x"30",	--4736
		x"0b",	--4737
		x"0a",	--4738
		x"09",	--4739
		x"08",	--4740
		x"18",	--4741
		x"0a",	--4742
		x"19",	--4743
		x"0c",	--4744
		x"1a",	--4745
		x"0e",	--4746
		x"1b",	--4747
		x"10",	--4748
		x"b0",	--4749
		x"a4",	--4750
		x"38",	--4751
		x"39",	--4752
		x"3a",	--4753
		x"3b",	--4754
		x"30",	--4755
		x"0b",	--4756
		x"0a",	--4757
		x"09",	--4758
		x"08",	--4759
		x"18",	--4760
		x"0a",	--4761
		x"19",	--4762
		x"0c",	--4763
		x"1a",	--4764
		x"0e",	--4765
		x"1b",	--4766
		x"10",	--4767
		x"b0",	--4768
		x"a4",	--4769
		x"0c",	--4770
		x"0d",	--4771
		x"0e",	--4772
		x"0f",	--4773
		x"38",	--4774
		x"39",	--4775
		x"3a",	--4776
		x"3b",	--4777
		x"30",	--4778
		x"0b",	--4779
		x"0a",	--4780
		x"09",	--4781
		x"08",	--4782
		x"07",	--4783
		x"18",	--4784
		x"0c",	--4785
		x"19",	--4786
		x"0e",	--4787
		x"1a",	--4788
		x"10",	--4789
		x"1b",	--4790
		x"12",	--4791
		x"b0",	--4792
		x"a4",	--4793
		x"17",	--4794
		x"14",	--4795
		x"87",	--4796
		x"00",	--4797
		x"87",	--4798
		x"02",	--4799
		x"87",	--4800
		x"04",	--4801
		x"87",	--4802
		x"06",	--4803
		x"37",	--4804
		x"38",	--4805
		x"39",	--4806
		x"3a",	--4807
		x"3b",	--4808
		x"30",	--4809
		x"00",	--4810
		x"32",	--4811
		x"f0",	--4812
		x"fd",	--4813
		x"57",	--4814
		x"69",	--4815
		x"69",	--4816
		x"67",	--4817
		x"66",	--4818
		x"72",	--4819
		x"61",	--4820
		x"6e",	--4821
		x"77",	--4822
		x"2e",	--4823
		x"69",	--4824
		x"20",	--4825
		x"69",	--4826
		x"65",	--4827
		x"0a",	--4828
		x"57",	--4829
		x"20",	--4830
		x"68",	--4831
		x"75",	--4832
		x"64",	--4833
		x"6e",	--4834
		x"74",	--4835
		x"73",	--4836
		x"65",	--4837
		x"74",	--4838
		x"61",	--4839
		x"0d",	--4840
		x"00",	--4841
		x"74",	--4842
		x"70",	--4843
		x"0a",	--4844
		x"65",	--4845
		x"72",	--4846
		x"72",	--4847
		x"20",	--4848
		x"69",	--4849
		x"73",	--4850
		x"6e",	--4851
		x"20",	--4852
		x"72",	--4853
		x"75",	--4854
		x"65",	--4855
		x"74",	--4856
		x"0a",	--4857
		x"63",	--4858
		x"72",	--4859
		x"65",	--4860
		x"74",	--4861
		x"75",	--4862
		x"61",	--4863
		x"65",	--4864
		x"0d",	--4865
		x"00",	--4866
		x"25",	--4867
		x"20",	--4868
		x"45",	--4869
		x"54",	--4870
		x"52",	--4871
		x"47",	--4872
		x"54",	--4873
		x"3c",	--4874
		x"49",	--4875
		x"45",	--4876
		x"55",	--4877
		x"3e",	--4878
		x"0a",	--4879
		x"25",	--4880
		x"20",	--4881
		x"64",	--4882
		x"0a",	--4883
		x"25",	--4884
		x"64",	--4885
		x"25",	--4886
		x"64",	--4887
		x"25",	--4888
		x"0d",	--4889
		x"00",	--4890
		x"34",	--4891
		x"5c",	--4892
		x"62",	--4893
		x"6a",	--4894
		x"72",	--4895
		x"7a",	--4896
		x"4c",	--4897
		x"54",	--4898
		x"0d",	--4899
		x"3d",	--4900
		x"3d",	--4901
		x"3d",	--4902
		x"20",	--4903
		x"61",	--4904
		x"63",	--4905
		x"6c",	--4906
		x"4d",	--4907
		x"55",	--4908
		x"3d",	--4909
		x"3d",	--4910
		x"3d",	--4911
		x"0d",	--4912
		x"00",	--4913
		x"6e",	--4914
		x"65",	--4915
		x"61",	--4916
		x"74",	--4917
		x"76",	--4918
		x"20",	--4919
		x"6f",	--4920
		x"65",	--4921
		x"77",	--4922
		x"69",	--4923
		x"65",	--4924
		x"72",	--4925
		x"61",	--4926
		x"00",	--4927
		x"77",	--4928
		x"00",	--4929
		x"6e",	--4930
		x"6f",	--4931
		x"65",	--4932
		x"00",	--4933
		x"70",	--4934
		x"65",	--4935
		x"20",	--4936
		x"6f",	--4937
		x"74",	--4938
		x"6f",	--4939
		x"6c",	--4940
		x"72",	--4941
		x"73",	--4942
		x"65",	--4943
		x"64",	--4944
		x"63",	--4945
		x"6e",	--4946
		x"69",	--4947
		x"75",	--4948
		x"61",	--4949
		x"69",	--4950
		x"6e",	--4951
		x"62",	--4952
		x"6f",	--4953
		x"6c",	--4954
		x"61",	--4955
		x"65",	--4956
		x"00",	--4957
		x"0a",	--4958
		x"08",	--4959
		x"08",	--4960
		x"25",	--4961
		x"00",	--4962
		x"77",	--4963
		x"69",	--4964
		x"65",	--4965
		x"0d",	--4966
		x"65",	--4967
		x"72",	--4968
		x"72",	--4969
		x"20",	--4970
		x"69",	--4971
		x"73",	--4972
		x"6e",	--4973
		x"20",	--4974
		x"72",	--4975
		x"75",	--4976
		x"65",	--4977
		x"74",	--4978
		x"0a",	--4979
		x"63",	--4980
		x"72",	--4981
		x"65",	--4982
		x"74",	--4983
		x"75",	--4984
		x"61",	--4985
		x"65",	--4986
		x"0d",	--4987
		x"00",	--4988
		x"25",	--4989
		x"20",	--4990
		x"45",	--4991
		x"49",	--4992
		x"54",	--4993
		x"52",	--4994
		x"56",	--4995
		x"4c",	--4996
		x"45",	--4997
		x"0a",	--4998
		x"72",	--4999
		x"25",	--5000
		x"20",	--5001
		x"3d",	--5002
		x"64",	--5003
		x"0a",	--5004
		x"09",	--5005
		x"73",	--5006
		x"52",	--5007
		x"47",	--5008
		x"53",	--5009
		x"45",	--5010
		x"0d",	--5011
		x"00",	--5012
		x"65",	--5013
		x"64",	--5014
		x"0d",	--5015
		x"25",	--5016
		x"20",	--5017
		x"73",	--5018
		x"6e",	--5019
		x"74",	--5020
		x"61",	--5021
		x"6e",	--5022
		x"6d",	--5023
		x"65",	--5024
		x"0d",	--5025
		x"00",	--5026
		x"63",	--5027
		x"25",	--5028
		x"0d",	--5029
		x"00",	--5030
		x"63",	--5031
		x"20",	--5032
		x"6f",	--5033
		x"73",	--5034
		x"63",	--5035
		x"20",	--5036
		x"6f",	--5037
		x"6d",	--5038
		x"6e",	--5039
		x"0d",	--5040
		x"00",	--5041
		x"4a",	--5042
		x"78",	--5043
		x"78",	--5044
		x"78",	--5045
		x"78",	--5046
		x"78",	--5047
		x"78",	--5048
		x"78",	--5049
		x"78",	--5050
		x"78",	--5051
		x"78",	--5052
		x"78",	--5053
		x"78",	--5054
		x"78",	--5055
		x"78",	--5056
		x"78",	--5057
		x"78",	--5058
		x"78",	--5059
		x"78",	--5060
		x"78",	--5061
		x"78",	--5062
		x"78",	--5063
		x"78",	--5064
		x"78",	--5065
		x"78",	--5066
		x"78",	--5067
		x"78",	--5068
		x"78",	--5069
		x"78",	--5070
		x"3c",	--5071
		x"78",	--5072
		x"78",	--5073
		x"78",	--5074
		x"78",	--5075
		x"78",	--5076
		x"78",	--5077
		x"78",	--5078
		x"78",	--5079
		x"78",	--5080
		x"78",	--5081
		x"78",	--5082
		x"78",	--5083
		x"78",	--5084
		x"78",	--5085
		x"78",	--5086
		x"78",	--5087
		x"78",	--5088
		x"78",	--5089
		x"78",	--5090
		x"78",	--5091
		x"78",	--5092
		x"78",	--5093
		x"78",	--5094
		x"78",	--5095
		x"78",	--5096
		x"78",	--5097
		x"78",	--5098
		x"78",	--5099
		x"78",	--5100
		x"78",	--5101
		x"78",	--5102
		x"2e",	--5103
		x"20",	--5104
		x"12",	--5105
		x"78",	--5106
		x"78",	--5107
		x"78",	--5108
		x"78",	--5109
		x"78",	--5110
		x"78",	--5111
		x"78",	--5112
		x"fa",	--5113
		x"78",	--5114
		x"e8",	--5115
		x"78",	--5116
		x"78",	--5117
		x"78",	--5118
		x"78",	--5119
		x"cc",	--5120
		x"78",	--5121
		x"78",	--5122
		x"78",	--5123
		x"be",	--5124
		x"ac",	--5125
		x"30",	--5126
		x"32",	--5127
		x"34",	--5128
		x"36",	--5129
		x"38",	--5130
		x"61",	--5131
		x"63",	--5132
		x"65",	--5133
		x"00",	--5134
		x"00",	--5135
		x"00",	--5136
		x"00",	--5137
		x"00",	--5138
		x"00",	--5139
		x"02",	--5140
		x"03",	--5141
		x"03",	--5142
		x"04",	--5143
		x"04",	--5144
		x"04",	--5145
		x"04",	--5146
		x"05",	--5147
		x"05",	--5148
		x"05",	--5149
		x"05",	--5150
		x"05",	--5151
		x"05",	--5152
		x"05",	--5153
		x"05",	--5154
		x"06",	--5155
		x"06",	--5156
		x"06",	--5157
		x"06",	--5158
		x"06",	--5159
		x"06",	--5160
		x"06",	--5161
		x"06",	--5162
		x"06",	--5163
		x"06",	--5164
		x"06",	--5165
		x"06",	--5166
		x"06",	--5167
		x"06",	--5168
		x"06",	--5169
		x"06",	--5170
		x"07",	--5171
		x"07",	--5172
		x"07",	--5173
		x"07",	--5174
		x"07",	--5175
		x"07",	--5176
		x"07",	--5177
		x"07",	--5178
		x"07",	--5179
		x"07",	--5180
		x"07",	--5181
		x"07",	--5182
		x"07",	--5183
		x"07",	--5184
		x"07",	--5185
		x"07",	--5186
		x"07",	--5187
		x"07",	--5188
		x"07",	--5189
		x"07",	--5190
		x"07",	--5191
		x"07",	--5192
		x"07",	--5193
		x"07",	--5194
		x"07",	--5195
		x"07",	--5196
		x"07",	--5197
		x"07",	--5198
		x"07",	--5199
		x"07",	--5200
		x"07",	--5201
		x"07",	--5202
		x"08",	--5203
		x"08",	--5204
		x"08",	--5205
		x"08",	--5206
		x"08",	--5207
		x"08",	--5208
		x"08",	--5209
		x"08",	--5210
		x"08",	--5211
		x"08",	--5212
		x"08",	--5213
		x"08",	--5214
		x"08",	--5215
		x"08",	--5216
		x"08",	--5217
		x"08",	--5218
		x"08",	--5219
		x"08",	--5220
		x"08",	--5221
		x"08",	--5222
		x"08",	--5223
		x"08",	--5224
		x"08",	--5225
		x"08",	--5226
		x"08",	--5227
		x"08",	--5228
		x"08",	--5229
		x"08",	--5230
		x"08",	--5231
		x"08",	--5232
		x"08",	--5233
		x"08",	--5234
		x"08",	--5235
		x"08",	--5236
		x"08",	--5237
		x"08",	--5238
		x"08",	--5239
		x"08",	--5240
		x"08",	--5241
		x"08",	--5242
		x"08",	--5243
		x"08",	--5244
		x"08",	--5245
		x"08",	--5246
		x"08",	--5247
		x"08",	--5248
		x"08",	--5249
		x"08",	--5250
		x"08",	--5251
		x"08",	--5252
		x"08",	--5253
		x"08",	--5254
		x"08",	--5255
		x"08",	--5256
		x"08",	--5257
		x"08",	--5258
		x"08",	--5259
		x"08",	--5260
		x"08",	--5261
		x"08",	--5262
		x"08",	--5263
		x"08",	--5264
		x"08",	--5265
		x"08",	--5266
		x"28",	--5267
		x"75",	--5268
		x"6c",	--5269
		x"00",	--5270
		x"ff",	--5271
		x"ff",	--5272
		x"68",	--5273
		x"6c",	--5274
		x"00",	--5275
		x"ff",	--5276
		x"ff",	--5277
		x"ff",	--5278
		x"ff",	--5279
		x"ff",	--5280
		x"ff",	--5281
		x"ff",	--5282
		x"ff",	--5283
		x"ff",	--5284
		x"ff",	--5285
		x"ff",	--5286
		x"ff",	--5287
		x"ff",	--5288
		x"ff",	--5289
		x"ff",	--5290
		x"ff",	--5291
		x"ff",	--5292
		x"ff",	--5293
		x"ff",	--5294
		x"ff",	--5295
		x"ff",	--5296
		x"ff",	--5297
		x"ff",	--5298
		x"ff",	--5299
		x"ff",	--5300
		x"ff",	--5301
		x"ff",	--5302
		x"ff",	--5303
		x"ff",	--5304
		x"ff",	--5305
		x"ff",	--5306
		x"ff",	--5307
		x"ff",	--5308
		x"ff",	--5309
		x"ff",	--5310
		x"ff",	--5311
		x"ff",	--5312
		x"ff",	--5313
		x"ff",	--5314
		x"ff",	--5315
		x"ff",	--5316
		x"ff",	--5317
		x"ff",	--5318
		x"ff",	--5319
		x"ff",	--5320
		x"ff",	--5321
		x"ff",	--5322
		x"ff",	--5323
		x"ff",	--5324
		x"ff",	--5325
		x"ff",	--5326
		x"ff",	--5327
		x"ff",	--5328
		x"ff",	--5329
		x"ff",	--5330
		x"ff",	--5331
		x"ff",	--5332
		x"ff",	--5333
		x"ff",	--5334
		x"ff",	--5335
		x"ff",	--5336
		x"ff",	--5337
		x"ff",	--5338
		x"ff",	--5339
		x"ff",	--5340
		x"ff",	--5341
		x"ff",	--5342
		x"ff",	--5343
		x"ff",	--5344
		x"ff",	--5345
		x"ff",	--5346
		x"ff",	--5347
		x"ff",	--5348
		x"ff",	--5349
		x"ff",	--5350
		x"ff",	--5351
		x"ff",	--5352
		x"ff",	--5353
		x"ff",	--5354
		x"ff",	--5355
		x"ff",	--5356
		x"ff",	--5357
		x"ff",	--5358
		x"ff",	--5359
		x"ff",	--5360
		x"ff",	--5361
		x"ff",	--5362
		x"ff",	--5363
		x"ff",	--5364
		x"ff",	--5365
		x"ff",	--5366
		x"ff",	--5367
		x"ff",	--5368
		x"ff",	--5369
		x"ff",	--5370
		x"ff",	--5371
		x"ff",	--5372
		x"ff",	--5373
		x"ff",	--5374
		x"ff",	--5375
		x"ff",	--5376
		x"ff",	--5377
		x"ff",	--5378
		x"ff",	--5379
		x"ff",	--5380
		x"ff",	--5381
		x"ff",	--5382
		x"ff",	--5383
		x"ff",	--5384
		x"ff",	--5385
		x"ff",	--5386
		x"ff",	--5387
		x"ff",	--5388
		x"ff",	--5389
		x"ff",	--5390
		x"ff",	--5391
		x"ff",	--5392
		x"ff",	--5393
		x"ff",	--5394
		x"ff",	--5395
		x"ff",	--5396
		x"ff",	--5397
		x"ff",	--5398
		x"ff",	--5399
		x"ff",	--5400
		x"ff",	--5401
		x"ff",	--5402
		x"ff",	--5403
		x"ff",	--5404
		x"ff",	--5405
		x"ff",	--5406
		x"ff",	--5407
		x"ff",	--5408
		x"ff",	--5409
		x"ff",	--5410
		x"ff",	--5411
		x"ff",	--5412
		x"ff",	--5413
		x"ff",	--5414
		x"ff",	--5415
		x"ff",	--5416
		x"ff",	--5417
		x"ff",	--5418
		x"ff",	--5419
		x"ff",	--5420
		x"ff",	--5421
		x"ff",	--5422
		x"ff",	--5423
		x"ff",	--5424
		x"ff",	--5425
		x"ff",	--5426
		x"ff",	--5427
		x"ff",	--5428
		x"ff",	--5429
		x"ff",	--5430
		x"ff",	--5431
		x"ff",	--5432
		x"ff",	--5433
		x"ff",	--5434
		x"ff",	--5435
		x"ff",	--5436
		x"ff",	--5437
		x"ff",	--5438
		x"ff",	--5439
		x"ff",	--5440
		x"ff",	--5441
		x"ff",	--5442
		x"ff",	--5443
		x"ff",	--5444
		x"ff",	--5445
		x"ff",	--5446
		x"ff",	--5447
		x"ff",	--5448
		x"ff",	--5449
		x"ff",	--5450
		x"ff",	--5451
		x"ff",	--5452
		x"ff",	--5453
		x"ff",	--5454
		x"ff",	--5455
		x"ff",	--5456
		x"ff",	--5457
		x"ff",	--5458
		x"ff",	--5459
		x"ff",	--5460
		x"ff",	--5461
		x"ff",	--5462
		x"ff",	--5463
		x"ff",	--5464
		x"ff",	--5465
		x"ff",	--5466
		x"ff",	--5467
		x"ff",	--5468
		x"ff",	--5469
		x"ff",	--5470
		x"ff",	--5471
		x"ff",	--5472
		x"ff",	--5473
		x"ff",	--5474
		x"ff",	--5475
		x"ff",	--5476
		x"ff",	--5477
		x"ff",	--5478
		x"ff",	--5479
		x"ff",	--5480
		x"ff",	--5481
		x"ff",	--5482
		x"ff",	--5483
		x"ff",	--5484
		x"ff",	--5485
		x"ff",	--5486
		x"ff",	--5487
		x"ff",	--5488
		x"ff",	--5489
		x"ff",	--5490
		x"ff",	--5491
		x"ff",	--5492
		x"ff",	--5493
		x"ff",	--5494
		x"ff",	--5495
		x"ff",	--5496
		x"ff",	--5497
		x"ff",	--5498
		x"ff",	--5499
		x"ff",	--5500
		x"ff",	--5501
		x"ff",	--5502
		x"ff",	--5503
		x"ff",	--5504
		x"ff",	--5505
		x"ff",	--5506
		x"ff",	--5507
		x"ff",	--5508
		x"ff",	--5509
		x"ff",	--5510
		x"ff",	--5511
		x"ff",	--5512
		x"ff",	--5513
		x"ff",	--5514
		x"ff",	--5515
		x"ff",	--5516
		x"ff",	--5517
		x"ff",	--5518
		x"ff",	--5519
		x"ff",	--5520
		x"ff",	--5521
		x"ff",	--5522
		x"ff",	--5523
		x"ff",	--5524
		x"ff",	--5525
		x"ff",	--5526
		x"ff",	--5527
		x"ff",	--5528
		x"ff",	--5529
		x"ff",	--5530
		x"ff",	--5531
		x"ff",	--5532
		x"ff",	--5533
		x"ff",	--5534
		x"ff",	--5535
		x"ff",	--5536
		x"ff",	--5537
		x"ff",	--5538
		x"ff",	--5539
		x"ff",	--5540
		x"ff",	--5541
		x"ff",	--5542
		x"ff",	--5543
		x"ff",	--5544
		x"ff",	--5545
		x"ff",	--5546
		x"ff",	--5547
		x"ff",	--5548
		x"ff",	--5549
		x"ff",	--5550
		x"ff",	--5551
		x"ff",	--5552
		x"ff",	--5553
		x"ff",	--5554
		x"ff",	--5555
		x"ff",	--5556
		x"ff",	--5557
		x"ff",	--5558
		x"ff",	--5559
		x"ff",	--5560
		x"ff",	--5561
		x"ff",	--5562
		x"ff",	--5563
		x"ff",	--5564
		x"ff",	--5565
		x"ff",	--5566
		x"ff",	--5567
		x"ff",	--5568
		x"ff",	--5569
		x"ff",	--5570
		x"ff",	--5571
		x"ff",	--5572
		x"ff",	--5573
		x"ff",	--5574
		x"ff",	--5575
		x"ff",	--5576
		x"ff",	--5577
		x"ff",	--5578
		x"ff",	--5579
		x"ff",	--5580
		x"ff",	--5581
		x"ff",	--5582
		x"ff",	--5583
		x"ff",	--5584
		x"ff",	--5585
		x"ff",	--5586
		x"ff",	--5587
		x"ff",	--5588
		x"ff",	--5589
		x"ff",	--5590
		x"ff",	--5591
		x"ff",	--5592
		x"ff",	--5593
		x"ff",	--5594
		x"ff",	--5595
		x"ff",	--5596
		x"ff",	--5597
		x"ff",	--5598
		x"ff",	--5599
		x"ff",	--5600
		x"ff",	--5601
		x"ff",	--5602
		x"ff",	--5603
		x"ff",	--5604
		x"ff",	--5605
		x"ff",	--5606
		x"ff",	--5607
		x"ff",	--5608
		x"ff",	--5609
		x"ff",	--5610
		x"ff",	--5611
		x"ff",	--5612
		x"ff",	--5613
		x"ff",	--5614
		x"ff",	--5615
		x"ff",	--5616
		x"ff",	--5617
		x"ff",	--5618
		x"ff",	--5619
		x"ff",	--5620
		x"ff",	--5621
		x"ff",	--5622
		x"ff",	--5623
		x"ff",	--5624
		x"ff",	--5625
		x"ff",	--5626
		x"ff",	--5627
		x"ff",	--5628
		x"ff",	--5629
		x"ff",	--5630
		x"ff",	--5631
		x"ff",	--5632
		x"ff",	--5633
		x"ff",	--5634
		x"ff",	--5635
		x"ff",	--5636
		x"ff",	--5637
		x"ff",	--5638
		x"ff",	--5639
		x"ff",	--5640
		x"ff",	--5641
		x"ff",	--5642
		x"ff",	--5643
		x"ff",	--5644
		x"ff",	--5645
		x"ff",	--5646
		x"ff",	--5647
		x"ff",	--5648
		x"ff",	--5649
		x"ff",	--5650
		x"ff",	--5651
		x"ff",	--5652
		x"ff",	--5653
		x"ff",	--5654
		x"ff",	--5655
		x"ff",	--5656
		x"ff",	--5657
		x"ff",	--5658
		x"ff",	--5659
		x"ff",	--5660
		x"ff",	--5661
		x"ff",	--5662
		x"ff",	--5663
		x"ff",	--5664
		x"ff",	--5665
		x"ff",	--5666
		x"ff",	--5667
		x"ff",	--5668
		x"ff",	--5669
		x"ff",	--5670
		x"ff",	--5671
		x"ff",	--5672
		x"ff",	--5673
		x"ff",	--5674
		x"ff",	--5675
		x"ff",	--5676
		x"ff",	--5677
		x"ff",	--5678
		x"ff",	--5679
		x"ff",	--5680
		x"ff",	--5681
		x"ff",	--5682
		x"ff",	--5683
		x"ff",	--5684
		x"ff",	--5685
		x"ff",	--5686
		x"ff",	--5687
		x"ff",	--5688
		x"ff",	--5689
		x"ff",	--5690
		x"ff",	--5691
		x"ff",	--5692
		x"ff",	--5693
		x"ff",	--5694
		x"ff",	--5695
		x"ff",	--5696
		x"ff",	--5697
		x"ff",	--5698
		x"ff",	--5699
		x"ff",	--5700
		x"ff",	--5701
		x"ff",	--5702
		x"ff",	--5703
		x"ff",	--5704
		x"ff",	--5705
		x"ff",	--5706
		x"ff",	--5707
		x"ff",	--5708
		x"ff",	--5709
		x"ff",	--5710
		x"ff",	--5711
		x"ff",	--5712
		x"ff",	--5713
		x"ff",	--5714
		x"ff",	--5715
		x"ff",	--5716
		x"ff",	--5717
		x"ff",	--5718
		x"ff",	--5719
		x"ff",	--5720
		x"ff",	--5721
		x"ff",	--5722
		x"ff",	--5723
		x"ff",	--5724
		x"ff",	--5725
		x"ff",	--5726
		x"ff",	--5727
		x"ff",	--5728
		x"ff",	--5729
		x"ff",	--5730
		x"ff",	--5731
		x"ff",	--5732
		x"ff",	--5733
		x"ff",	--5734
		x"ff",	--5735
		x"ff",	--5736
		x"ff",	--5737
		x"ff",	--5738
		x"ff",	--5739
		x"ff",	--5740
		x"ff",	--5741
		x"ff",	--5742
		x"ff",	--5743
		x"ff",	--5744
		x"ff",	--5745
		x"ff",	--5746
		x"ff",	--5747
		x"ff",	--5748
		x"ff",	--5749
		x"ff",	--5750
		x"ff",	--5751
		x"ff",	--5752
		x"ff",	--5753
		x"ff",	--5754
		x"ff",	--5755
		x"ff",	--5756
		x"ff",	--5757
		x"ff",	--5758
		x"ff",	--5759
		x"ff",	--5760
		x"ff",	--5761
		x"ff",	--5762
		x"ff",	--5763
		x"ff",	--5764
		x"ff",	--5765
		x"ff",	--5766
		x"ff",	--5767
		x"ff",	--5768
		x"ff",	--5769
		x"ff",	--5770
		x"ff",	--5771
		x"ff",	--5772
		x"ff",	--5773
		x"ff",	--5774
		x"ff",	--5775
		x"ff",	--5776
		x"ff",	--5777
		x"ff",	--5778
		x"ff",	--5779
		x"ff",	--5780
		x"ff",	--5781
		x"ff",	--5782
		x"ff",	--5783
		x"ff",	--5784
		x"ff",	--5785
		x"ff",	--5786
		x"ff",	--5787
		x"ff",	--5788
		x"ff",	--5789
		x"ff",	--5790
		x"ff",	--5791
		x"ff",	--5792
		x"ff",	--5793
		x"ff",	--5794
		x"ff",	--5795
		x"ff",	--5796
		x"ff",	--5797
		x"ff",	--5798
		x"ff",	--5799
		x"ff",	--5800
		x"ff",	--5801
		x"ff",	--5802
		x"ff",	--5803
		x"ff",	--5804
		x"ff",	--5805
		x"ff",	--5806
		x"ff",	--5807
		x"ff",	--5808
		x"ff",	--5809
		x"ff",	--5810
		x"ff",	--5811
		x"ff",	--5812
		x"ff",	--5813
		x"ff",	--5814
		x"ff",	--5815
		x"ff",	--5816
		x"ff",	--5817
		x"ff",	--5818
		x"ff",	--5819
		x"ff",	--5820
		x"ff",	--5821
		x"ff",	--5822
		x"ff",	--5823
		x"ff",	--5824
		x"ff",	--5825
		x"ff",	--5826
		x"ff",	--5827
		x"ff",	--5828
		x"ff",	--5829
		x"ff",	--5830
		x"ff",	--5831
		x"ff",	--5832
		x"ff",	--5833
		x"ff",	--5834
		x"ff",	--5835
		x"ff",	--5836
		x"ff",	--5837
		x"ff",	--5838
		x"ff",	--5839
		x"ff",	--5840
		x"ff",	--5841
		x"ff",	--5842
		x"ff",	--5843
		x"ff",	--5844
		x"ff",	--5845
		x"ff",	--5846
		x"ff",	--5847
		x"ff",	--5848
		x"ff",	--5849
		x"ff",	--5850
		x"ff",	--5851
		x"ff",	--5852
		x"ff",	--5853
		x"ff",	--5854
		x"ff",	--5855
		x"ff",	--5856
		x"ff",	--5857
		x"ff",	--5858
		x"ff",	--5859
		x"ff",	--5860
		x"ff",	--5861
		x"ff",	--5862
		x"ff",	--5863
		x"ff",	--5864
		x"ff",	--5865
		x"ff",	--5866
		x"ff",	--5867
		x"ff",	--5868
		x"ff",	--5869
		x"ff",	--5870
		x"ff",	--5871
		x"ff",	--5872
		x"ff",	--5873
		x"ff",	--5874
		x"ff",	--5875
		x"ff",	--5876
		x"ff",	--5877
		x"ff",	--5878
		x"ff",	--5879
		x"ff",	--5880
		x"ff",	--5881
		x"ff",	--5882
		x"ff",	--5883
		x"ff",	--5884
		x"ff",	--5885
		x"ff",	--5886
		x"ff",	--5887
		x"ff",	--5888
		x"ff",	--5889
		x"ff",	--5890
		x"ff",	--5891
		x"ff",	--5892
		x"ff",	--5893
		x"ff",	--5894
		x"ff",	--5895
		x"ff",	--5896
		x"ff",	--5897
		x"ff",	--5898
		x"ff",	--5899
		x"ff",	--5900
		x"ff",	--5901
		x"ff",	--5902
		x"ff",	--5903
		x"ff",	--5904
		x"ff",	--5905
		x"ff",	--5906
		x"ff",	--5907
		x"ff",	--5908
		x"ff",	--5909
		x"ff",	--5910
		x"ff",	--5911
		x"ff",	--5912
		x"ff",	--5913
		x"ff",	--5914
		x"ff",	--5915
		x"ff",	--5916
		x"ff",	--5917
		x"ff",	--5918
		x"ff",	--5919
		x"ff",	--5920
		x"ff",	--5921
		x"ff",	--5922
		x"ff",	--5923
		x"ff",	--5924
		x"ff",	--5925
		x"ff",	--5926
		x"ff",	--5927
		x"ff",	--5928
		x"ff",	--5929
		x"ff",	--5930
		x"ff",	--5931
		x"ff",	--5932
		x"ff",	--5933
		x"ff",	--5934
		x"ff",	--5935
		x"ff",	--5936
		x"ff",	--5937
		x"ff",	--5938
		x"ff",	--5939
		x"ff",	--5940
		x"ff",	--5941
		x"ff",	--5942
		x"ff",	--5943
		x"ff",	--5944
		x"ff",	--5945
		x"ff",	--5946
		x"ff",	--5947
		x"ff",	--5948
		x"ff",	--5949
		x"ff",	--5950
		x"ff",	--5951
		x"ff",	--5952
		x"ff",	--5953
		x"ff",	--5954
		x"ff",	--5955
		x"ff",	--5956
		x"ff",	--5957
		x"ff",	--5958
		x"ff",	--5959
		x"ff",	--5960
		x"ff",	--5961
		x"ff",	--5962
		x"ff",	--5963
		x"ff",	--5964
		x"ff",	--5965
		x"ff",	--5966
		x"ff",	--5967
		x"ff",	--5968
		x"ff",	--5969
		x"ff",	--5970
		x"ff",	--5971
		x"ff",	--5972
		x"ff",	--5973
		x"ff",	--5974
		x"ff",	--5975
		x"ff",	--5976
		x"ff",	--5977
		x"ff",	--5978
		x"ff",	--5979
		x"ff",	--5980
		x"ff",	--5981
		x"ff",	--5982
		x"ff",	--5983
		x"ff",	--5984
		x"ff",	--5985
		x"ff",	--5986
		x"ff",	--5987
		x"ff",	--5988
		x"ff",	--5989
		x"ff",	--5990
		x"ff",	--5991
		x"ff",	--5992
		x"ff",	--5993
		x"ff",	--5994
		x"ff",	--5995
		x"ff",	--5996
		x"ff",	--5997
		x"ff",	--5998
		x"ff",	--5999
		x"ff",	--6000
		x"ff",	--6001
		x"ff",	--6002
		x"ff",	--6003
		x"ff",	--6004
		x"ff",	--6005
		x"ff",	--6006
		x"ff",	--6007
		x"ff",	--6008
		x"ff",	--6009
		x"ff",	--6010
		x"ff",	--6011
		x"ff",	--6012
		x"ff",	--6013
		x"ff",	--6014
		x"ff",	--6015
		x"ff",	--6016
		x"ff",	--6017
		x"ff",	--6018
		x"ff",	--6019
		x"ff",	--6020
		x"ff",	--6021
		x"ff",	--6022
		x"ff",	--6023
		x"ff",	--6024
		x"ff",	--6025
		x"ff",	--6026
		x"ff",	--6027
		x"ff",	--6028
		x"ff",	--6029
		x"ff",	--6030
		x"ff",	--6031
		x"ff",	--6032
		x"ff",	--6033
		x"ff",	--6034
		x"ff",	--6035
		x"ff",	--6036
		x"ff",	--6037
		x"ff",	--6038
		x"ff",	--6039
		x"ff",	--6040
		x"ff",	--6041
		x"ff",	--6042
		x"ff",	--6043
		x"ff",	--6044
		x"ff",	--6045
		x"ff",	--6046
		x"ff",	--6047
		x"ff",	--6048
		x"ff",	--6049
		x"ff",	--6050
		x"ff",	--6051
		x"ff",	--6052
		x"ff",	--6053
		x"ff",	--6054
		x"ff",	--6055
		x"ff",	--6056
		x"ff",	--6057
		x"ff",	--6058
		x"ff",	--6059
		x"ff",	--6060
		x"ff",	--6061
		x"ff",	--6062
		x"ff",	--6063
		x"ff",	--6064
		x"ff",	--6065
		x"ff",	--6066
		x"ff",	--6067
		x"ff",	--6068
		x"ff",	--6069
		x"ff",	--6070
		x"ff",	--6071
		x"ff",	--6072
		x"ff",	--6073
		x"ff",	--6074
		x"ff",	--6075
		x"ff",	--6076
		x"ff",	--6077
		x"ff",	--6078
		x"ff",	--6079
		x"ff",	--6080
		x"ff",	--6081
		x"ff",	--6082
		x"ff",	--6083
		x"ff",	--6084
		x"ff",	--6085
		x"ff",	--6086
		x"ff",	--6087
		x"ff",	--6088
		x"ff",	--6089
		x"ff",	--6090
		x"ff",	--6091
		x"ff",	--6092
		x"ff",	--6093
		x"ff",	--6094
		x"ff",	--6095
		x"ff",	--6096
		x"ff",	--6097
		x"ff",	--6098
		x"ff",	--6099
		x"ff",	--6100
		x"ff",	--6101
		x"ff",	--6102
		x"ff",	--6103
		x"ff",	--6104
		x"ff",	--6105
		x"ff",	--6106
		x"ff",	--6107
		x"ff",	--6108
		x"ff",	--6109
		x"ff",	--6110
		x"ff",	--6111
		x"ff",	--6112
		x"ff",	--6113
		x"ff",	--6114
		x"ff",	--6115
		x"ff",	--6116
		x"ff",	--6117
		x"ff",	--6118
		x"ff",	--6119
		x"ff",	--6120
		x"ff",	--6121
		x"ff",	--6122
		x"ff",	--6123
		x"ff",	--6124
		x"ff",	--6125
		x"ff",	--6126
		x"ff",	--6127
		x"ff",	--6128
		x"ff",	--6129
		x"ff",	--6130
		x"ff",	--6131
		x"ff",	--6132
		x"ff",	--6133
		x"ff",	--6134
		x"ff",	--6135
		x"ff",	--6136
		x"ff",	--6137
		x"ff",	--6138
		x"ff",	--6139
		x"ff",	--6140
		x"ff",	--6141
		x"ff",	--6142
		x"ff",	--6143
		x"ff",	--6144
		x"ff",	--6145
		x"ff",	--6146
		x"ff",	--6147
		x"ff",	--6148
		x"ff",	--6149
		x"ff",	--6150
		x"ff",	--6151
		x"ff",	--6152
		x"ff",	--6153
		x"ff",	--6154
		x"ff",	--6155
		x"ff",	--6156
		x"ff",	--6157
		x"ff",	--6158
		x"ff",	--6159
		x"ff",	--6160
		x"ff",	--6161
		x"ff",	--6162
		x"ff",	--6163
		x"ff",	--6164
		x"ff",	--6165
		x"ff",	--6166
		x"ff",	--6167
		x"ff",	--6168
		x"ff",	--6169
		x"ff",	--6170
		x"ff",	--6171
		x"ff",	--6172
		x"ff",	--6173
		x"ff",	--6174
		x"ff",	--6175
		x"ff",	--6176
		x"ff",	--6177
		x"ff",	--6178
		x"ff",	--6179
		x"ff",	--6180
		x"ff",	--6181
		x"ff",	--6182
		x"ff",	--6183
		x"ff",	--6184
		x"ff",	--6185
		x"ff",	--6186
		x"ff",	--6187
		x"ff",	--6188
		x"ff",	--6189
		x"ff",	--6190
		x"ff",	--6191
		x"ff",	--6192
		x"ff",	--6193
		x"ff",	--6194
		x"ff",	--6195
		x"ff",	--6196
		x"ff",	--6197
		x"ff",	--6198
		x"ff",	--6199
		x"ff",	--6200
		x"ff",	--6201
		x"ff",	--6202
		x"ff",	--6203
		x"ff",	--6204
		x"ff",	--6205
		x"ff",	--6206
		x"ff",	--6207
		x"ff",	--6208
		x"ff",	--6209
		x"ff",	--6210
		x"ff",	--6211
		x"ff",	--6212
		x"ff",	--6213
		x"ff",	--6214
		x"ff",	--6215
		x"ff",	--6216
		x"ff",	--6217
		x"ff",	--6218
		x"ff",	--6219
		x"ff",	--6220
		x"ff",	--6221
		x"ff",	--6222
		x"ff",	--6223
		x"ff",	--6224
		x"ff",	--6225
		x"ff",	--6226
		x"ff",	--6227
		x"ff",	--6228
		x"ff",	--6229
		x"ff",	--6230
		x"ff",	--6231
		x"ff",	--6232
		x"ff",	--6233
		x"ff",	--6234
		x"ff",	--6235
		x"ff",	--6236
		x"ff",	--6237
		x"ff",	--6238
		x"ff",	--6239
		x"ff",	--6240
		x"ff",	--6241
		x"ff",	--6242
		x"ff",	--6243
		x"ff",	--6244
		x"ff",	--6245
		x"ff",	--6246
		x"ff",	--6247
		x"ff",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"ff",	--6252
		x"ff",	--6253
		x"ff",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"2e",	--8176
		x"2e",	--8177
		x"2e",	--8178
		x"2e",	--8179
		x"2e",	--8180
		x"2e",	--8181
		x"2e",	--8182
		x"54",	--8183
		x"d6",	--8184
		x"2e",	--8185
		x"2e",	--8186
		x"2e",	--8187
		x"2e",	--8188
		x"2e",	--8189
		x"2e",	--8190
		x"00");	--8191
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"e9",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"cd",	--44
		x"12",	--45
		x"c8",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"e6",	--50
		x"12",	--51
		x"cc",	--52
		x"53",	--53
		x"40",	--54
		x"e6",	--55
		x"40",	--56
		x"c5",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"c8",	--61
		x"40",	--62
		x"e6",	--63
		x"40",	--64
		x"c5",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"c8",	--69
		x"40",	--70
		x"e6",	--71
		x"40",	--72
		x"c5",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"c8",	--77
		x"40",	--78
		x"e6",	--79
		x"40",	--80
		x"c3",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"c8",	--85
		x"40",	--86
		x"e6",	--87
		x"40",	--88
		x"c4",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"c8",	--93
		x"40",	--94
		x"e6",	--95
		x"40",	--96
		x"c2",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"c8",	--101
		x"40",	--102
		x"e6",	--103
		x"40",	--104
		x"c2",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"c8",	--109
		x"40",	--110
		x"e6",	--111
		x"40",	--112
		x"c2",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"c8",	--117
		x"43",	--118
		x"43",	--119
		x"12",	--120
		x"c8",	--121
		x"43",	--122
		x"40",	--123
		x"4e",	--124
		x"40",	--125
		x"01",	--126
		x"41",	--127
		x"50",	--128
		x"00",	--129
		x"12",	--130
		x"c7",	--131
		x"41",	--132
		x"50",	--133
		x"00",	--134
		x"12",	--135
		x"c7",	--136
		x"43",	--137
		x"40",	--138
		x"4e",	--139
		x"40",	--140
		x"01",	--141
		x"41",	--142
		x"52",	--143
		x"12",	--144
		x"c7",	--145
		x"41",	--146
		x"52",	--147
		x"12",	--148
		x"c7",	--149
		x"41",	--150
		x"52",	--151
		x"41",	--152
		x"50",	--153
		x"00",	--154
		x"12",	--155
		x"c3",	--156
		x"40",	--157
		x"01",	--158
		x"41",	--159
		x"53",	--160
		x"12",	--161
		x"ca",	--162
		x"40",	--163
		x"01",	--164
		x"41",	--165
		x"12",	--166
		x"ca",	--167
		x"41",	--168
		x"41",	--169
		x"53",	--170
		x"12",	--171
		x"c4",	--172
		x"12",	--173
		x"c9",	--174
		x"40",	--175
		x"00",	--176
		x"40",	--177
		x"c4",	--178
		x"12",	--179
		x"c9",	--180
		x"43",	--181
		x"40",	--182
		x"03",	--183
		x"12",	--184
		x"c9",	--185
		x"43",	--186
		x"43",	--187
		x"43",	--188
		x"41",	--189
		x"50",	--190
		x"00",	--191
		x"12",	--192
		x"c3",	--193
		x"43",	--194
		x"43",	--195
		x"43",	--196
		x"41",	--197
		x"50",	--198
		x"00",	--199
		x"12",	--200
		x"c3",	--201
		x"41",	--202
		x"50",	--203
		x"00",	--204
		x"41",	--205
		x"50",	--206
		x"00",	--207
		x"12",	--208
		x"c2",	--209
		x"40",	--210
		x"ff",	--211
		x"00",	--212
		x"d2",	--213
		x"43",	--214
		x"12",	--215
		x"cd",	--216
		x"93",	--217
		x"27",	--218
		x"12",	--219
		x"cd",	--220
		x"92",	--221
		x"24",	--222
		x"90",	--223
		x"00",	--224
		x"20",	--225
		x"12",	--226
		x"e6",	--227
		x"12",	--228
		x"cc",	--229
		x"53",	--230
		x"40",	--231
		x"00",	--232
		x"51",	--233
		x"5f",	--234
		x"43",	--235
		x"00",	--236
		x"4f",	--237
		x"41",	--238
		x"00",	--239
		x"12",	--240
		x"c8",	--241
		x"43",	--242
		x"3f",	--243
		x"93",	--244
		x"27",	--245
		x"53",	--246
		x"12",	--247
		x"e6",	--248
		x"12",	--249
		x"cc",	--250
		x"53",	--251
		x"3f",	--252
		x"90",	--253
		x"00",	--254
		x"2f",	--255
		x"93",	--256
		x"02",	--257
		x"24",	--258
		x"4f",	--259
		x"11",	--260
		x"12",	--261
		x"12",	--262
		x"e6",	--263
		x"4f",	--264
		x"00",	--265
		x"12",	--266
		x"cc",	--267
		x"52",	--268
		x"41",	--269
		x"00",	--270
		x"40",	--271
		x"00",	--272
		x"51",	--273
		x"5b",	--274
		x"4f",	--275
		x"00",	--276
		x"53",	--277
		x"3f",	--278
		x"40",	--279
		x"e5",	--280
		x"4e",	--281
		x"00",	--282
		x"4d",	--283
		x"00",	--284
		x"4c",	--285
		x"00",	--286
		x"43",	--287
		x"00",	--288
		x"43",	--289
		x"00",	--290
		x"43",	--291
		x"00",	--292
		x"41",	--293
		x"43",	--294
		x"00",	--295
		x"43",	--296
		x"00",	--297
		x"43",	--298
		x"00",	--299
		x"41",	--300
		x"4e",	--301
		x"00",	--302
		x"41",	--303
		x"4e",	--304
		x"00",	--305
		x"41",	--306
		x"4e",	--307
		x"00",	--308
		x"41",	--309
		x"4e",	--310
		x"00",	--311
		x"41",	--312
		x"4f",	--313
		x"00",	--314
		x"8e",	--315
		x"4d",	--316
		x"5f",	--317
		x"00",	--318
		x"4d",	--319
		x"00",	--320
		x"12",	--321
		x"c2",	--322
		x"43",	--323
		x"4e",	--324
		x"01",	--325
		x"4f",	--326
		x"01",	--327
		x"42",	--328
		x"01",	--329
		x"41",	--330
		x"12",	--331
		x"c2",	--332
		x"43",	--333
		x"4d",	--334
		x"01",	--335
		x"4f",	--336
		x"00",	--337
		x"01",	--338
		x"42",	--339
		x"01",	--340
		x"41",	--341
		x"5c",	--342
		x"8f",	--343
		x"00",	--344
		x"12",	--345
		x"c2",	--346
		x"43",	--347
		x"4e",	--348
		x"01",	--349
		x"4f",	--350
		x"00",	--351
		x"01",	--352
		x"42",	--353
		x"01",	--354
		x"41",	--355
		x"5d",	--356
		x"41",	--357
		x"41",	--358
		x"43",	--359
		x"41",	--360
		x"43",	--361
		x"41",	--362
		x"40",	--363
		x"c0",	--364
		x"01",	--365
		x"40",	--366
		x"00",	--367
		x"01",	--368
		x"40",	--369
		x"02",	--370
		x"01",	--371
		x"12",	--372
		x"e5",	--373
		x"12",	--374
		x"cc",	--375
		x"43",	--376
		x"01",	--377
		x"40",	--378
		x"e5",	--379
		x"00",	--380
		x"12",	--381
		x"cc",	--382
		x"53",	--383
		x"43",	--384
		x"41",	--385
		x"12",	--386
		x"c2",	--387
		x"41",	--388
		x"12",	--389
		x"12",	--390
		x"43",	--391
		x"40",	--392
		x"3f",	--393
		x"4a",	--394
		x"4b",	--395
		x"42",	--396
		x"02",	--397
		x"12",	--398
		x"c7",	--399
		x"4a",	--400
		x"4b",	--401
		x"42",	--402
		x"02",	--403
		x"12",	--404
		x"c7",	--405
		x"12",	--406
		x"e5",	--407
		x"12",	--408
		x"cc",	--409
		x"53",	--410
		x"41",	--411
		x"41",	--412
		x"41",	--413
		x"4f",	--414
		x"02",	--415
		x"4e",	--416
		x"02",	--417
		x"41",	--418
		x"12",	--419
		x"12",	--420
		x"83",	--421
		x"4f",	--422
		x"4e",	--423
		x"93",	--424
		x"02",	--425
		x"24",	--426
		x"90",	--427
		x"00",	--428
		x"38",	--429
		x"20",	--430
		x"41",	--431
		x"4b",	--432
		x"00",	--433
		x"12",	--434
		x"c6",	--435
		x"4f",	--436
		x"41",	--437
		x"4b",	--438
		x"00",	--439
		x"12",	--440
		x"c6",	--441
		x"4f",	--442
		x"12",	--443
		x"12",	--444
		x"12",	--445
		x"e6",	--446
		x"12",	--447
		x"cc",	--448
		x"50",	--449
		x"00",	--450
		x"4a",	--451
		x"43",	--452
		x"12",	--453
		x"d5",	--454
		x"43",	--455
		x"40",	--456
		x"42",	--457
		x"12",	--458
		x"d3",	--459
		x"4e",	--460
		x"4f",	--461
		x"42",	--462
		x"02",	--463
		x"12",	--464
		x"c7",	--465
		x"4b",	--466
		x"43",	--467
		x"12",	--468
		x"d5",	--469
		x"43",	--470
		x"40",	--471
		x"42",	--472
		x"12",	--473
		x"d3",	--474
		x"4e",	--475
		x"4f",	--476
		x"42",	--477
		x"02",	--478
		x"12",	--479
		x"c7",	--480
		x"43",	--481
		x"53",	--482
		x"41",	--483
		x"41",	--484
		x"41",	--485
		x"41",	--486
		x"4b",	--487
		x"00",	--488
		x"12",	--489
		x"c6",	--490
		x"43",	--491
		x"4f",	--492
		x"42",	--493
		x"02",	--494
		x"12",	--495
		x"c9",	--496
		x"3f",	--497
		x"43",	--498
		x"40",	--499
		x"c3",	--500
		x"12",	--501
		x"c9",	--502
		x"4f",	--503
		x"02",	--504
		x"3f",	--505
		x"12",	--506
		x"e5",	--507
		x"12",	--508
		x"cc",	--509
		x"40",	--510
		x"e5",	--511
		x"00",	--512
		x"12",	--513
		x"cc",	--514
		x"4b",	--515
		x"00",	--516
		x"12",	--517
		x"e6",	--518
		x"12",	--519
		x"cc",	--520
		x"52",	--521
		x"43",	--522
		x"3f",	--523
		x"12",	--524
		x"12",	--525
		x"42",	--526
		x"02",	--527
		x"12",	--528
		x"ca",	--529
		x"4e",	--530
		x"4f",	--531
		x"42",	--532
		x"02",	--533
		x"12",	--534
		x"ca",	--535
		x"12",	--536
		x"12",	--537
		x"12",	--538
		x"12",	--539
		x"12",	--540
		x"e6",	--541
		x"12",	--542
		x"02",	--543
		x"12",	--544
		x"db",	--545
		x"50",	--546
		x"00",	--547
		x"12",	--548
		x"02",	--549
		x"12",	--550
		x"e6",	--551
		x"12",	--552
		x"cc",	--553
		x"52",	--554
		x"41",	--555
		x"41",	--556
		x"41",	--557
		x"4f",	--558
		x"02",	--559
		x"4e",	--560
		x"02",	--561
		x"41",	--562
		x"12",	--563
		x"12",	--564
		x"12",	--565
		x"83",	--566
		x"4f",	--567
		x"4e",	--568
		x"43",	--569
		x"00",	--570
		x"93",	--571
		x"24",	--572
		x"93",	--573
		x"02",	--574
		x"24",	--575
		x"43",	--576
		x"02",	--577
		x"41",	--578
		x"4b",	--579
		x"00",	--580
		x"12",	--581
		x"c6",	--582
		x"4f",	--583
		x"90",	--584
		x"00",	--585
		x"34",	--586
		x"43",	--587
		x"49",	--588
		x"42",	--589
		x"02",	--590
		x"12",	--591
		x"c9",	--592
		x"43",	--593
		x"53",	--594
		x"41",	--595
		x"41",	--596
		x"41",	--597
		x"41",	--598
		x"93",	--599
		x"02",	--600
		x"24",	--601
		x"43",	--602
		x"02",	--603
		x"42",	--604
		x"02",	--605
		x"12",	--606
		x"c9",	--607
		x"43",	--608
		x"53",	--609
		x"41",	--610
		x"41",	--611
		x"41",	--612
		x"41",	--613
		x"41",	--614
		x"4b",	--615
		x"00",	--616
		x"12",	--617
		x"c6",	--618
		x"4f",	--619
		x"3f",	--620
		x"43",	--621
		x"12",	--622
		x"c4",	--623
		x"43",	--624
		x"53",	--625
		x"41",	--626
		x"41",	--627
		x"41",	--628
		x"41",	--629
		x"43",	--630
		x"40",	--631
		x"c4",	--632
		x"12",	--633
		x"c9",	--634
		x"4f",	--635
		x"02",	--636
		x"3f",	--637
		x"42",	--638
		x"00",	--639
		x"4e",	--640
		x"be",	--641
		x"20",	--642
		x"df",	--643
		x"00",	--644
		x"41",	--645
		x"cf",	--646
		x"00",	--647
		x"41",	--648
		x"43",	--649
		x"93",	--650
		x"02",	--651
		x"24",	--652
		x"43",	--653
		x"4f",	--654
		x"02",	--655
		x"43",	--656
		x"41",	--657
		x"42",	--658
		x"02",	--659
		x"92",	--660
		x"2c",	--661
		x"4e",	--662
		x"5f",	--663
		x"4f",	--664
		x"e6",	--665
		x"43",	--666
		x"00",	--667
		x"90",	--668
		x"00",	--669
		x"38",	--670
		x"43",	--671
		x"02",	--672
		x"41",	--673
		x"53",	--674
		x"4e",	--675
		x"02",	--676
		x"41",	--677
		x"40",	--678
		x"00",	--679
		x"00",	--680
		x"3f",	--681
		x"40",	--682
		x"00",	--683
		x"00",	--684
		x"3f",	--685
		x"42",	--686
		x"00",	--687
		x"3f",	--688
		x"40",	--689
		x"00",	--690
		x"00",	--691
		x"3f",	--692
		x"40",	--693
		x"00",	--694
		x"00",	--695
		x"3f",	--696
		x"40",	--697
		x"00",	--698
		x"00",	--699
		x"3f",	--700
		x"40",	--701
		x"00",	--702
		x"00",	--703
		x"3f",	--704
		x"12",	--705
		x"12",	--706
		x"83",	--707
		x"4f",	--708
		x"4e",	--709
		x"12",	--710
		x"e6",	--711
		x"12",	--712
		x"cc",	--713
		x"53",	--714
		x"90",	--715
		x"00",	--716
		x"38",	--717
		x"41",	--718
		x"4b",	--719
		x"00",	--720
		x"12",	--721
		x"c6",	--722
		x"4f",	--723
		x"41",	--724
		x"4b",	--725
		x"00",	--726
		x"12",	--727
		x"c6",	--728
		x"4f",	--729
		x"12",	--730
		x"12",	--731
		x"12",	--732
		x"e7",	--733
		x"12",	--734
		x"cc",	--735
		x"50",	--736
		x"00",	--737
		x"4b",	--738
		x"00",	--739
		x"43",	--740
		x"53",	--741
		x"41",	--742
		x"41",	--743
		x"41",	--744
		x"12",	--745
		x"e6",	--746
		x"12",	--747
		x"cc",	--748
		x"40",	--749
		x"e6",	--750
		x"00",	--751
		x"12",	--752
		x"cc",	--753
		x"4b",	--754
		x"00",	--755
		x"12",	--756
		x"e6",	--757
		x"12",	--758
		x"cc",	--759
		x"52",	--760
		x"43",	--761
		x"3f",	--762
		x"12",	--763
		x"83",	--764
		x"4e",	--765
		x"93",	--766
		x"24",	--767
		x"38",	--768
		x"12",	--769
		x"e7",	--770
		x"12",	--771
		x"cc",	--772
		x"53",	--773
		x"41",	--774
		x"4b",	--775
		x"00",	--776
		x"12",	--777
		x"c6",	--778
		x"12",	--779
		x"12",	--780
		x"12",	--781
		x"e7",	--782
		x"12",	--783
		x"cc",	--784
		x"50",	--785
		x"00",	--786
		x"43",	--787
		x"53",	--788
		x"41",	--789
		x"41",	--790
		x"12",	--791
		x"e6",	--792
		x"12",	--793
		x"cc",	--794
		x"40",	--795
		x"e6",	--796
		x"00",	--797
		x"12",	--798
		x"cc",	--799
		x"4b",	--800
		x"00",	--801
		x"12",	--802
		x"e7",	--803
		x"12",	--804
		x"cc",	--805
		x"52",	--806
		x"43",	--807
		x"3f",	--808
		x"12",	--809
		x"12",	--810
		x"43",	--811
		x"00",	--812
		x"4f",	--813
		x"93",	--814
		x"24",	--815
		x"53",	--816
		x"43",	--817
		x"43",	--818
		x"3c",	--819
		x"90",	--820
		x"00",	--821
		x"2c",	--822
		x"5c",	--823
		x"5c",	--824
		x"5c",	--825
		x"5c",	--826
		x"11",	--827
		x"5d",	--828
		x"50",	--829
		x"ff",	--830
		x"43",	--831
		x"4f",	--832
		x"93",	--833
		x"24",	--834
		x"90",	--835
		x"00",	--836
		x"24",	--837
		x"4d",	--838
		x"50",	--839
		x"ff",	--840
		x"93",	--841
		x"23",	--842
		x"90",	--843
		x"00",	--844
		x"2c",	--845
		x"5c",	--846
		x"4c",	--847
		x"5b",	--848
		x"5b",	--849
		x"5b",	--850
		x"11",	--851
		x"5d",	--852
		x"50",	--853
		x"ff",	--854
		x"4f",	--855
		x"93",	--856
		x"23",	--857
		x"43",	--858
		x"00",	--859
		x"4c",	--860
		x"41",	--861
		x"41",	--862
		x"41",	--863
		x"43",	--864
		x"3f",	--865
		x"4d",	--866
		x"50",	--867
		x"ff",	--868
		x"90",	--869
		x"00",	--870
		x"2c",	--871
		x"5c",	--872
		x"5c",	--873
		x"5c",	--874
		x"5c",	--875
		x"11",	--876
		x"5d",	--877
		x"50",	--878
		x"ff",	--879
		x"43",	--880
		x"3f",	--881
		x"4d",	--882
		x"50",	--883
		x"ff",	--884
		x"90",	--885
		x"00",	--886
		x"2c",	--887
		x"5c",	--888
		x"5c",	--889
		x"5c",	--890
		x"5c",	--891
		x"11",	--892
		x"5d",	--893
		x"50",	--894
		x"ff",	--895
		x"43",	--896
		x"3f",	--897
		x"11",	--898
		x"12",	--899
		x"12",	--900
		x"e7",	--901
		x"12",	--902
		x"cc",	--903
		x"52",	--904
		x"43",	--905
		x"4c",	--906
		x"41",	--907
		x"41",	--908
		x"41",	--909
		x"43",	--910
		x"3f",	--911
		x"12",	--912
		x"12",	--913
		x"4e",	--914
		x"4c",	--915
		x"4e",	--916
		x"00",	--917
		x"4d",	--918
		x"00",	--919
		x"4c",	--920
		x"00",	--921
		x"4d",	--922
		x"43",	--923
		x"40",	--924
		x"36",	--925
		x"40",	--926
		x"01",	--927
		x"12",	--928
		x"e4",	--929
		x"4e",	--930
		x"00",	--931
		x"12",	--932
		x"c2",	--933
		x"43",	--934
		x"4a",	--935
		x"01",	--936
		x"40",	--937
		x"00",	--938
		x"01",	--939
		x"42",	--940
		x"01",	--941
		x"00",	--942
		x"41",	--943
		x"43",	--944
		x"41",	--945
		x"41",	--946
		x"41",	--947
		x"12",	--948
		x"12",	--949
		x"12",	--950
		x"43",	--951
		x"00",	--952
		x"40",	--953
		x"3f",	--954
		x"00",	--955
		x"4f",	--956
		x"4b",	--957
		x"00",	--958
		x"43",	--959
		x"12",	--960
		x"d5",	--961
		x"43",	--962
		x"40",	--963
		x"3f",	--964
		x"12",	--965
		x"d1",	--966
		x"4e",	--967
		x"4f",	--968
		x"4b",	--969
		x"00",	--970
		x"43",	--971
		x"12",	--972
		x"d5",	--973
		x"4e",	--974
		x"4f",	--975
		x"48",	--976
		x"49",	--977
		x"12",	--978
		x"d1",	--979
		x"12",	--980
		x"ce",	--981
		x"4e",	--982
		x"00",	--983
		x"43",	--984
		x"00",	--985
		x"41",	--986
		x"41",	--987
		x"41",	--988
		x"41",	--989
		x"12",	--990
		x"12",	--991
		x"12",	--992
		x"4d",	--993
		x"4e",	--994
		x"4d",	--995
		x"00",	--996
		x"4e",	--997
		x"00",	--998
		x"4f",	--999
		x"49",	--1000
		x"00",	--1001
		x"43",	--1002
		x"12",	--1003
		x"d5",	--1004
		x"4e",	--1005
		x"4f",	--1006
		x"4a",	--1007
		x"4b",	--1008
		x"12",	--1009
		x"d1",	--1010
		x"4e",	--1011
		x"4f",	--1012
		x"49",	--1013
		x"00",	--1014
		x"43",	--1015
		x"12",	--1016
		x"d5",	--1017
		x"4e",	--1018
		x"4f",	--1019
		x"4a",	--1020
		x"4b",	--1021
		x"12",	--1022
		x"d1",	--1023
		x"12",	--1024
		x"ce",	--1025
		x"4e",	--1026
		x"00",	--1027
		x"41",	--1028
		x"41",	--1029
		x"41",	--1030
		x"41",	--1031
		x"12",	--1032
		x"12",	--1033
		x"93",	--1034
		x"02",	--1035
		x"38",	--1036
		x"40",	--1037
		x"02",	--1038
		x"43",	--1039
		x"12",	--1040
		x"4b",	--1041
		x"ff",	--1042
		x"11",	--1043
		x"12",	--1044
		x"12",	--1045
		x"e7",	--1046
		x"12",	--1047
		x"cc",	--1048
		x"50",	--1049
		x"00",	--1050
		x"53",	--1051
		x"50",	--1052
		x"00",	--1053
		x"92",	--1054
		x"02",	--1055
		x"3b",	--1056
		x"43",	--1057
		x"41",	--1058
		x"41",	--1059
		x"41",	--1060
		x"42",	--1061
		x"02",	--1062
		x"90",	--1063
		x"00",	--1064
		x"34",	--1065
		x"4e",	--1066
		x"5f",	--1067
		x"5e",	--1068
		x"5f",	--1069
		x"50",	--1070
		x"02",	--1071
		x"40",	--1072
		x"00",	--1073
		x"00",	--1074
		x"40",	--1075
		x"c8",	--1076
		x"00",	--1077
		x"40",	--1078
		x"02",	--1079
		x"00",	--1080
		x"53",	--1081
		x"4e",	--1082
		x"02",	--1083
		x"41",	--1084
		x"12",	--1085
		x"42",	--1086
		x"02",	--1087
		x"90",	--1088
		x"00",	--1089
		x"34",	--1090
		x"4b",	--1091
		x"5c",	--1092
		x"5b",	--1093
		x"5c",	--1094
		x"50",	--1095
		x"02",	--1096
		x"4f",	--1097
		x"00",	--1098
		x"4e",	--1099
		x"00",	--1100
		x"4d",	--1101
		x"00",	--1102
		x"53",	--1103
		x"4b",	--1104
		x"02",	--1105
		x"43",	--1106
		x"41",	--1107
		x"41",	--1108
		x"43",	--1109
		x"3f",	--1110
		x"12",	--1111
		x"50",	--1112
		x"ff",	--1113
		x"42",	--1114
		x"02",	--1115
		x"93",	--1116
		x"38",	--1117
		x"92",	--1118
		x"02",	--1119
		x"24",	--1120
		x"40",	--1121
		x"02",	--1122
		x"43",	--1123
		x"3c",	--1124
		x"50",	--1125
		x"00",	--1126
		x"9f",	--1127
		x"ff",	--1128
		x"24",	--1129
		x"53",	--1130
		x"9b",	--1131
		x"23",	--1132
		x"12",	--1133
		x"e7",	--1134
		x"12",	--1135
		x"cc",	--1136
		x"53",	--1137
		x"43",	--1138
		x"50",	--1139
		x"00",	--1140
		x"41",	--1141
		x"41",	--1142
		x"43",	--1143
		x"4e",	--1144
		x"00",	--1145
		x"4e",	--1146
		x"93",	--1147
		x"24",	--1148
		x"53",	--1149
		x"43",	--1150
		x"3c",	--1151
		x"4e",	--1152
		x"93",	--1153
		x"24",	--1154
		x"53",	--1155
		x"92",	--1156
		x"34",	--1157
		x"90",	--1158
		x"00",	--1159
		x"23",	--1160
		x"43",	--1161
		x"ff",	--1162
		x"4f",	--1163
		x"5d",	--1164
		x"51",	--1165
		x"4e",	--1166
		x"00",	--1167
		x"53",	--1168
		x"4e",	--1169
		x"93",	--1170
		x"23",	--1171
		x"4c",	--1172
		x"5e",	--1173
		x"5e",	--1174
		x"5c",	--1175
		x"50",	--1176
		x"02",	--1177
		x"41",	--1178
		x"12",	--1179
		x"00",	--1180
		x"50",	--1181
		x"00",	--1182
		x"41",	--1183
		x"41",	--1184
		x"43",	--1185
		x"3f",	--1186
		x"d0",	--1187
		x"02",	--1188
		x"01",	--1189
		x"40",	--1190
		x"0b",	--1191
		x"01",	--1192
		x"43",	--1193
		x"41",	--1194
		x"12",	--1195
		x"4f",	--1196
		x"42",	--1197
		x"02",	--1198
		x"90",	--1199
		x"00",	--1200
		x"34",	--1201
		x"4f",	--1202
		x"5c",	--1203
		x"4c",	--1204
		x"5d",	--1205
		x"5d",	--1206
		x"5d",	--1207
		x"8c",	--1208
		x"50",	--1209
		x"03",	--1210
		x"43",	--1211
		x"00",	--1212
		x"43",	--1213
		x"00",	--1214
		x"43",	--1215
		x"00",	--1216
		x"4b",	--1217
		x"00",	--1218
		x"4e",	--1219
		x"00",	--1220
		x"4f",	--1221
		x"53",	--1222
		x"4e",	--1223
		x"02",	--1224
		x"41",	--1225
		x"41",	--1226
		x"43",	--1227
		x"3f",	--1228
		x"5f",	--1229
		x"4f",	--1230
		x"5c",	--1231
		x"5c",	--1232
		x"5c",	--1233
		x"8f",	--1234
		x"50",	--1235
		x"03",	--1236
		x"43",	--1237
		x"00",	--1238
		x"4e",	--1239
		x"00",	--1240
		x"43",	--1241
		x"00",	--1242
		x"4d",	--1243
		x"00",	--1244
		x"43",	--1245
		x"00",	--1246
		x"43",	--1247
		x"41",	--1248
		x"5f",	--1249
		x"4f",	--1250
		x"5e",	--1251
		x"5e",	--1252
		x"5e",	--1253
		x"8f",	--1254
		x"43",	--1255
		x"03",	--1256
		x"43",	--1257
		x"41",	--1258
		x"12",	--1259
		x"12",	--1260
		x"12",	--1261
		x"12",	--1262
		x"12",	--1263
		x"12",	--1264
		x"12",	--1265
		x"12",	--1266
		x"12",	--1267
		x"93",	--1268
		x"02",	--1269
		x"38",	--1270
		x"40",	--1271
		x"03",	--1272
		x"4a",	--1273
		x"53",	--1274
		x"4a",	--1275
		x"52",	--1276
		x"4a",	--1277
		x"50",	--1278
		x"00",	--1279
		x"43",	--1280
		x"3c",	--1281
		x"53",	--1282
		x"4f",	--1283
		x"00",	--1284
		x"53",	--1285
		x"50",	--1286
		x"00",	--1287
		x"50",	--1288
		x"00",	--1289
		x"50",	--1290
		x"00",	--1291
		x"50",	--1292
		x"00",	--1293
		x"92",	--1294
		x"02",	--1295
		x"34",	--1296
		x"93",	--1297
		x"00",	--1298
		x"27",	--1299
		x"4b",	--1300
		x"9b",	--1301
		x"00",	--1302
		x"2b",	--1303
		x"43",	--1304
		x"00",	--1305
		x"4b",	--1306
		x"00",	--1307
		x"12",	--1308
		x"00",	--1309
		x"93",	--1310
		x"00",	--1311
		x"27",	--1312
		x"47",	--1313
		x"53",	--1314
		x"4f",	--1315
		x"00",	--1316
		x"98",	--1317
		x"2b",	--1318
		x"43",	--1319
		x"00",	--1320
		x"3f",	--1321
		x"f0",	--1322
		x"ff",	--1323
		x"01",	--1324
		x"41",	--1325
		x"41",	--1326
		x"41",	--1327
		x"41",	--1328
		x"41",	--1329
		x"41",	--1330
		x"41",	--1331
		x"41",	--1332
		x"41",	--1333
		x"13",	--1334
		x"4e",	--1335
		x"00",	--1336
		x"43",	--1337
		x"41",	--1338
		x"4f",	--1339
		x"4f",	--1340
		x"4f",	--1341
		x"00",	--1342
		x"41",	--1343
		x"42",	--1344
		x"00",	--1345
		x"f2",	--1346
		x"23",	--1347
		x"4f",	--1348
		x"00",	--1349
		x"43",	--1350
		x"41",	--1351
		x"f0",	--1352
		x"00",	--1353
		x"4f",	--1354
		x"e8",	--1355
		x"11",	--1356
		x"12",	--1357
		x"ca",	--1358
		x"41",	--1359
		x"12",	--1360
		x"4f",	--1361
		x"4f",	--1362
		x"11",	--1363
		x"11",	--1364
		x"11",	--1365
		x"11",	--1366
		x"4e",	--1367
		x"12",	--1368
		x"ca",	--1369
		x"4b",	--1370
		x"12",	--1371
		x"ca",	--1372
		x"41",	--1373
		x"41",	--1374
		x"12",	--1375
		x"12",	--1376
		x"4f",	--1377
		x"40",	--1378
		x"00",	--1379
		x"4a",	--1380
		x"4b",	--1381
		x"f0",	--1382
		x"00",	--1383
		x"24",	--1384
		x"11",	--1385
		x"53",	--1386
		x"23",	--1387
		x"f3",	--1388
		x"24",	--1389
		x"40",	--1390
		x"00",	--1391
		x"12",	--1392
		x"ca",	--1393
		x"53",	--1394
		x"93",	--1395
		x"23",	--1396
		x"41",	--1397
		x"41",	--1398
		x"41",	--1399
		x"40",	--1400
		x"00",	--1401
		x"3f",	--1402
		x"12",	--1403
		x"4f",	--1404
		x"4f",	--1405
		x"10",	--1406
		x"11",	--1407
		x"4e",	--1408
		x"12",	--1409
		x"ca",	--1410
		x"4b",	--1411
		x"12",	--1412
		x"ca",	--1413
		x"41",	--1414
		x"41",	--1415
		x"12",	--1416
		x"12",	--1417
		x"4e",	--1418
		x"4f",	--1419
		x"4f",	--1420
		x"10",	--1421
		x"11",	--1422
		x"4d",	--1423
		x"12",	--1424
		x"ca",	--1425
		x"4b",	--1426
		x"12",	--1427
		x"ca",	--1428
		x"4b",	--1429
		x"4a",	--1430
		x"10",	--1431
		x"10",	--1432
		x"ec",	--1433
		x"ec",	--1434
		x"4d",	--1435
		x"12",	--1436
		x"ca",	--1437
		x"4a",	--1438
		x"12",	--1439
		x"ca",	--1440
		x"41",	--1441
		x"41",	--1442
		x"41",	--1443
		x"12",	--1444
		x"12",	--1445
		x"12",	--1446
		x"4f",	--1447
		x"93",	--1448
		x"24",	--1449
		x"4e",	--1450
		x"53",	--1451
		x"43",	--1452
		x"4a",	--1453
		x"5b",	--1454
		x"4d",	--1455
		x"11",	--1456
		x"12",	--1457
		x"ca",	--1458
		x"99",	--1459
		x"24",	--1460
		x"53",	--1461
		x"b0",	--1462
		x"00",	--1463
		x"20",	--1464
		x"40",	--1465
		x"00",	--1466
		x"12",	--1467
		x"ca",	--1468
		x"3f",	--1469
		x"40",	--1470
		x"00",	--1471
		x"12",	--1472
		x"ca",	--1473
		x"3f",	--1474
		x"41",	--1475
		x"41",	--1476
		x"41",	--1477
		x"41",	--1478
		x"12",	--1479
		x"12",	--1480
		x"12",	--1481
		x"4f",	--1482
		x"93",	--1483
		x"24",	--1484
		x"4e",	--1485
		x"53",	--1486
		x"43",	--1487
		x"4a",	--1488
		x"11",	--1489
		x"12",	--1490
		x"ca",	--1491
		x"99",	--1492
		x"24",	--1493
		x"53",	--1494
		x"b0",	--1495
		x"00",	--1496
		x"23",	--1497
		x"40",	--1498
		x"00",	--1499
		x"12",	--1500
		x"ca",	--1501
		x"4a",	--1502
		x"11",	--1503
		x"12",	--1504
		x"ca",	--1505
		x"99",	--1506
		x"23",	--1507
		x"41",	--1508
		x"41",	--1509
		x"41",	--1510
		x"41",	--1511
		x"12",	--1512
		x"12",	--1513
		x"12",	--1514
		x"50",	--1515
		x"ff",	--1516
		x"4f",	--1517
		x"93",	--1518
		x"38",	--1519
		x"90",	--1520
		x"00",	--1521
		x"38",	--1522
		x"43",	--1523
		x"41",	--1524
		x"59",	--1525
		x"40",	--1526
		x"00",	--1527
		x"4b",	--1528
		x"12",	--1529
		x"e3",	--1530
		x"50",	--1531
		x"00",	--1532
		x"4f",	--1533
		x"00",	--1534
		x"53",	--1535
		x"40",	--1536
		x"00",	--1537
		x"4b",	--1538
		x"12",	--1539
		x"e3",	--1540
		x"4f",	--1541
		x"90",	--1542
		x"00",	--1543
		x"37",	--1544
		x"49",	--1545
		x"53",	--1546
		x"51",	--1547
		x"40",	--1548
		x"00",	--1549
		x"4b",	--1550
		x"12",	--1551
		x"e3",	--1552
		x"50",	--1553
		x"00",	--1554
		x"4f",	--1555
		x"00",	--1556
		x"53",	--1557
		x"41",	--1558
		x"5a",	--1559
		x"4f",	--1560
		x"11",	--1561
		x"12",	--1562
		x"ca",	--1563
		x"93",	--1564
		x"23",	--1565
		x"50",	--1566
		x"00",	--1567
		x"41",	--1568
		x"41",	--1569
		x"41",	--1570
		x"41",	--1571
		x"40",	--1572
		x"00",	--1573
		x"12",	--1574
		x"ca",	--1575
		x"e3",	--1576
		x"53",	--1577
		x"3f",	--1578
		x"43",	--1579
		x"43",	--1580
		x"3f",	--1581
		x"12",	--1582
		x"12",	--1583
		x"12",	--1584
		x"41",	--1585
		x"52",	--1586
		x"4b",	--1587
		x"49",	--1588
		x"93",	--1589
		x"20",	--1590
		x"3c",	--1591
		x"11",	--1592
		x"12",	--1593
		x"ca",	--1594
		x"49",	--1595
		x"4a",	--1596
		x"53",	--1597
		x"4a",	--1598
		x"00",	--1599
		x"93",	--1600
		x"24",	--1601
		x"90",	--1602
		x"00",	--1603
		x"23",	--1604
		x"49",	--1605
		x"53",	--1606
		x"49",	--1607
		x"00",	--1608
		x"50",	--1609
		x"ff",	--1610
		x"90",	--1611
		x"00",	--1612
		x"2f",	--1613
		x"4f",	--1614
		x"5f",	--1615
		x"4f",	--1616
		x"e7",	--1617
		x"41",	--1618
		x"41",	--1619
		x"41",	--1620
		x"41",	--1621
		x"4b",	--1622
		x"52",	--1623
		x"4b",	--1624
		x"00",	--1625
		x"4b",	--1626
		x"12",	--1627
		x"cb",	--1628
		x"49",	--1629
		x"3f",	--1630
		x"4b",	--1631
		x"53",	--1632
		x"4b",	--1633
		x"12",	--1634
		x"ca",	--1635
		x"49",	--1636
		x"3f",	--1637
		x"4b",	--1638
		x"53",	--1639
		x"4f",	--1640
		x"49",	--1641
		x"93",	--1642
		x"27",	--1643
		x"53",	--1644
		x"11",	--1645
		x"12",	--1646
		x"ca",	--1647
		x"49",	--1648
		x"93",	--1649
		x"23",	--1650
		x"3f",	--1651
		x"4b",	--1652
		x"52",	--1653
		x"4b",	--1654
		x"00",	--1655
		x"4b",	--1656
		x"12",	--1657
		x"cb",	--1658
		x"49",	--1659
		x"3f",	--1660
		x"4b",	--1661
		x"53",	--1662
		x"4b",	--1663
		x"4e",	--1664
		x"10",	--1665
		x"11",	--1666
		x"10",	--1667
		x"11",	--1668
		x"12",	--1669
		x"cb",	--1670
		x"49",	--1671
		x"3f",	--1672
		x"4b",	--1673
		x"53",	--1674
		x"4b",	--1675
		x"12",	--1676
		x"cb",	--1677
		x"49",	--1678
		x"3f",	--1679
		x"4b",	--1680
		x"53",	--1681
		x"4b",	--1682
		x"12",	--1683
		x"ca",	--1684
		x"49",	--1685
		x"3f",	--1686
		x"4b",	--1687
		x"53",	--1688
		x"4b",	--1689
		x"12",	--1690
		x"ca",	--1691
		x"49",	--1692
		x"3f",	--1693
		x"4b",	--1694
		x"53",	--1695
		x"4b",	--1696
		x"12",	--1697
		x"ca",	--1698
		x"49",	--1699
		x"3f",	--1700
		x"40",	--1701
		x"00",	--1702
		x"12",	--1703
		x"ca",	--1704
		x"3f",	--1705
		x"12",	--1706
		x"12",	--1707
		x"42",	--1708
		x"02",	--1709
		x"42",	--1710
		x"00",	--1711
		x"04",	--1712
		x"42",	--1713
		x"02",	--1714
		x"90",	--1715
		x"00",	--1716
		x"34",	--1717
		x"53",	--1718
		x"02",	--1719
		x"42",	--1720
		x"02",	--1721
		x"42",	--1722
		x"02",	--1723
		x"9f",	--1724
		x"20",	--1725
		x"53",	--1726
		x"02",	--1727
		x"40",	--1728
		x"00",	--1729
		x"00",	--1730
		x"41",	--1731
		x"41",	--1732
		x"c0",	--1733
		x"00",	--1734
		x"00",	--1735
		x"13",	--1736
		x"43",	--1737
		x"02",	--1738
		x"3f",	--1739
		x"4e",	--1740
		x"4f",	--1741
		x"40",	--1742
		x"36",	--1743
		x"40",	--1744
		x"01",	--1745
		x"12",	--1746
		x"e3",	--1747
		x"53",	--1748
		x"4e",	--1749
		x"00",	--1750
		x"40",	--1751
		x"00",	--1752
		x"00",	--1753
		x"41",	--1754
		x"42",	--1755
		x"02",	--1756
		x"42",	--1757
		x"02",	--1758
		x"9f",	--1759
		x"38",	--1760
		x"42",	--1761
		x"02",	--1762
		x"82",	--1763
		x"02",	--1764
		x"41",	--1765
		x"42",	--1766
		x"02",	--1767
		x"42",	--1768
		x"02",	--1769
		x"40",	--1770
		x"00",	--1771
		x"8d",	--1772
		x"8e",	--1773
		x"41",	--1774
		x"42",	--1775
		x"02",	--1776
		x"4f",	--1777
		x"04",	--1778
		x"42",	--1779
		x"02",	--1780
		x"42",	--1781
		x"02",	--1782
		x"9e",	--1783
		x"24",	--1784
		x"42",	--1785
		x"02",	--1786
		x"90",	--1787
		x"00",	--1788
		x"38",	--1789
		x"43",	--1790
		x"02",	--1791
		x"41",	--1792
		x"53",	--1793
		x"02",	--1794
		x"41",	--1795
		x"43",	--1796
		x"41",	--1797
		x"12",	--1798
		x"12",	--1799
		x"4e",	--1800
		x"4f",	--1801
		x"43",	--1802
		x"40",	--1803
		x"4f",	--1804
		x"12",	--1805
		x"d4",	--1806
		x"93",	--1807
		x"34",	--1808
		x"4a",	--1809
		x"4b",	--1810
		x"12",	--1811
		x"d5",	--1812
		x"41",	--1813
		x"41",	--1814
		x"41",	--1815
		x"43",	--1816
		x"40",	--1817
		x"4f",	--1818
		x"4a",	--1819
		x"4b",	--1820
		x"12",	--1821
		x"d1",	--1822
		x"12",	--1823
		x"d5",	--1824
		x"53",	--1825
		x"60",	--1826
		x"80",	--1827
		x"41",	--1828
		x"41",	--1829
		x"41",	--1830
		x"12",	--1831
		x"12",	--1832
		x"12",	--1833
		x"12",	--1834
		x"12",	--1835
		x"12",	--1836
		x"12",	--1837
		x"12",	--1838
		x"50",	--1839
		x"ff",	--1840
		x"4d",	--1841
		x"4f",	--1842
		x"93",	--1843
		x"28",	--1844
		x"4e",	--1845
		x"93",	--1846
		x"28",	--1847
		x"92",	--1848
		x"20",	--1849
		x"40",	--1850
		x"d0",	--1851
		x"92",	--1852
		x"24",	--1853
		x"93",	--1854
		x"24",	--1855
		x"93",	--1856
		x"24",	--1857
		x"4f",	--1858
		x"00",	--1859
		x"00",	--1860
		x"4e",	--1861
		x"00",	--1862
		x"4f",	--1863
		x"00",	--1864
		x"4f",	--1865
		x"00",	--1866
		x"4e",	--1867
		x"00",	--1868
		x"4e",	--1869
		x"00",	--1870
		x"41",	--1871
		x"8b",	--1872
		x"4c",	--1873
		x"93",	--1874
		x"38",	--1875
		x"90",	--1876
		x"00",	--1877
		x"34",	--1878
		x"93",	--1879
		x"38",	--1880
		x"46",	--1881
		x"00",	--1882
		x"47",	--1883
		x"00",	--1884
		x"49",	--1885
		x"f0",	--1886
		x"00",	--1887
		x"24",	--1888
		x"46",	--1889
		x"47",	--1890
		x"c3",	--1891
		x"10",	--1892
		x"10",	--1893
		x"53",	--1894
		x"23",	--1895
		x"4a",	--1896
		x"00",	--1897
		x"4b",	--1898
		x"00",	--1899
		x"43",	--1900
		x"43",	--1901
		x"f0",	--1902
		x"00",	--1903
		x"24",	--1904
		x"5c",	--1905
		x"6d",	--1906
		x"53",	--1907
		x"23",	--1908
		x"53",	--1909
		x"63",	--1910
		x"f6",	--1911
		x"f7",	--1912
		x"43",	--1913
		x"43",	--1914
		x"93",	--1915
		x"20",	--1916
		x"93",	--1917
		x"24",	--1918
		x"41",	--1919
		x"00",	--1920
		x"41",	--1921
		x"00",	--1922
		x"da",	--1923
		x"db",	--1924
		x"4f",	--1925
		x"00",	--1926
		x"9e",	--1927
		x"00",	--1928
		x"20",	--1929
		x"4f",	--1930
		x"00",	--1931
		x"41",	--1932
		x"00",	--1933
		x"46",	--1934
		x"47",	--1935
		x"54",	--1936
		x"65",	--1937
		x"4e",	--1938
		x"00",	--1939
		x"4f",	--1940
		x"00",	--1941
		x"40",	--1942
		x"00",	--1943
		x"00",	--1944
		x"93",	--1945
		x"38",	--1946
		x"48",	--1947
		x"50",	--1948
		x"00",	--1949
		x"41",	--1950
		x"41",	--1951
		x"41",	--1952
		x"41",	--1953
		x"41",	--1954
		x"41",	--1955
		x"41",	--1956
		x"41",	--1957
		x"41",	--1958
		x"91",	--1959
		x"38",	--1960
		x"4b",	--1961
		x"00",	--1962
		x"43",	--1963
		x"43",	--1964
		x"4f",	--1965
		x"00",	--1966
		x"9e",	--1967
		x"00",	--1968
		x"27",	--1969
		x"93",	--1970
		x"24",	--1971
		x"46",	--1972
		x"47",	--1973
		x"84",	--1974
		x"75",	--1975
		x"93",	--1976
		x"38",	--1977
		x"43",	--1978
		x"00",	--1979
		x"41",	--1980
		x"00",	--1981
		x"4e",	--1982
		x"00",	--1983
		x"4f",	--1984
		x"00",	--1985
		x"4e",	--1986
		x"4f",	--1987
		x"53",	--1988
		x"63",	--1989
		x"90",	--1990
		x"3f",	--1991
		x"28",	--1992
		x"90",	--1993
		x"40",	--1994
		x"2c",	--1995
		x"93",	--1996
		x"2c",	--1997
		x"48",	--1998
		x"00",	--1999
		x"53",	--2000
		x"5e",	--2001
		x"6f",	--2002
		x"4b",	--2003
		x"53",	--2004
		x"4e",	--2005
		x"4f",	--2006
		x"53",	--2007
		x"63",	--2008
		x"90",	--2009
		x"3f",	--2010
		x"2b",	--2011
		x"24",	--2012
		x"4e",	--2013
		x"00",	--2014
		x"4f",	--2015
		x"00",	--2016
		x"4a",	--2017
		x"00",	--2018
		x"40",	--2019
		x"00",	--2020
		x"00",	--2021
		x"93",	--2022
		x"37",	--2023
		x"4e",	--2024
		x"4f",	--2025
		x"f3",	--2026
		x"f3",	--2027
		x"c3",	--2028
		x"10",	--2029
		x"10",	--2030
		x"4c",	--2031
		x"4d",	--2032
		x"de",	--2033
		x"df",	--2034
		x"4a",	--2035
		x"00",	--2036
		x"4b",	--2037
		x"00",	--2038
		x"53",	--2039
		x"00",	--2040
		x"48",	--2041
		x"3f",	--2042
		x"93",	--2043
		x"23",	--2044
		x"4f",	--2045
		x"00",	--2046
		x"4f",	--2047
		x"00",	--2048
		x"00",	--2049
		x"4f",	--2050
		x"00",	--2051
		x"00",	--2052
		x"4f",	--2053
		x"00",	--2054
		x"00",	--2055
		x"4e",	--2056
		x"00",	--2057
		x"ff",	--2058
		x"00",	--2059
		x"4e",	--2060
		x"00",	--2061
		x"4d",	--2062
		x"3f",	--2063
		x"43",	--2064
		x"43",	--2065
		x"3f",	--2066
		x"e3",	--2067
		x"53",	--2068
		x"90",	--2069
		x"00",	--2070
		x"37",	--2071
		x"3f",	--2072
		x"93",	--2073
		x"2b",	--2074
		x"3f",	--2075
		x"44",	--2076
		x"45",	--2077
		x"86",	--2078
		x"77",	--2079
		x"3f",	--2080
		x"4e",	--2081
		x"3f",	--2082
		x"43",	--2083
		x"00",	--2084
		x"41",	--2085
		x"00",	--2086
		x"e3",	--2087
		x"e3",	--2088
		x"53",	--2089
		x"63",	--2090
		x"4e",	--2091
		x"00",	--2092
		x"4f",	--2093
		x"00",	--2094
		x"3f",	--2095
		x"93",	--2096
		x"27",	--2097
		x"59",	--2098
		x"00",	--2099
		x"44",	--2100
		x"00",	--2101
		x"45",	--2102
		x"00",	--2103
		x"49",	--2104
		x"f0",	--2105
		x"00",	--2106
		x"24",	--2107
		x"4d",	--2108
		x"44",	--2109
		x"45",	--2110
		x"c3",	--2111
		x"10",	--2112
		x"10",	--2113
		x"53",	--2114
		x"23",	--2115
		x"4c",	--2116
		x"00",	--2117
		x"4d",	--2118
		x"00",	--2119
		x"43",	--2120
		x"43",	--2121
		x"f0",	--2122
		x"00",	--2123
		x"24",	--2124
		x"5c",	--2125
		x"6d",	--2126
		x"53",	--2127
		x"23",	--2128
		x"53",	--2129
		x"63",	--2130
		x"f4",	--2131
		x"f5",	--2132
		x"43",	--2133
		x"43",	--2134
		x"93",	--2135
		x"20",	--2136
		x"93",	--2137
		x"20",	--2138
		x"43",	--2139
		x"43",	--2140
		x"41",	--2141
		x"00",	--2142
		x"41",	--2143
		x"00",	--2144
		x"da",	--2145
		x"db",	--2146
		x"3f",	--2147
		x"43",	--2148
		x"43",	--2149
		x"3f",	--2150
		x"92",	--2151
		x"23",	--2152
		x"9e",	--2153
		x"00",	--2154
		x"00",	--2155
		x"27",	--2156
		x"40",	--2157
		x"e8",	--2158
		x"3f",	--2159
		x"50",	--2160
		x"ff",	--2161
		x"4e",	--2162
		x"00",	--2163
		x"4f",	--2164
		x"00",	--2165
		x"4c",	--2166
		x"00",	--2167
		x"4d",	--2168
		x"00",	--2169
		x"41",	--2170
		x"50",	--2171
		x"00",	--2172
		x"41",	--2173
		x"52",	--2174
		x"12",	--2175
		x"d9",	--2176
		x"41",	--2177
		x"50",	--2178
		x"00",	--2179
		x"41",	--2180
		x"12",	--2181
		x"d9",	--2182
		x"41",	--2183
		x"52",	--2184
		x"41",	--2185
		x"50",	--2186
		x"00",	--2187
		x"41",	--2188
		x"50",	--2189
		x"00",	--2190
		x"12",	--2191
		x"ce",	--2192
		x"12",	--2193
		x"d7",	--2194
		x"50",	--2195
		x"00",	--2196
		x"41",	--2197
		x"50",	--2198
		x"ff",	--2199
		x"4e",	--2200
		x"00",	--2201
		x"4f",	--2202
		x"00",	--2203
		x"4c",	--2204
		x"00",	--2205
		x"4d",	--2206
		x"00",	--2207
		x"41",	--2208
		x"50",	--2209
		x"00",	--2210
		x"41",	--2211
		x"52",	--2212
		x"12",	--2213
		x"d9",	--2214
		x"41",	--2215
		x"50",	--2216
		x"00",	--2217
		x"41",	--2218
		x"12",	--2219
		x"d9",	--2220
		x"e3",	--2221
		x"00",	--2222
		x"41",	--2223
		x"52",	--2224
		x"41",	--2225
		x"50",	--2226
		x"00",	--2227
		x"41",	--2228
		x"50",	--2229
		x"00",	--2230
		x"12",	--2231
		x"ce",	--2232
		x"12",	--2233
		x"d7",	--2234
		x"50",	--2235
		x"00",	--2236
		x"41",	--2237
		x"12",	--2238
		x"12",	--2239
		x"12",	--2240
		x"12",	--2241
		x"12",	--2242
		x"12",	--2243
		x"12",	--2244
		x"12",	--2245
		x"50",	--2246
		x"ff",	--2247
		x"4e",	--2248
		x"00",	--2249
		x"4f",	--2250
		x"00",	--2251
		x"4c",	--2252
		x"00",	--2253
		x"4d",	--2254
		x"00",	--2255
		x"41",	--2256
		x"50",	--2257
		x"00",	--2258
		x"41",	--2259
		x"52",	--2260
		x"12",	--2261
		x"d9",	--2262
		x"41",	--2263
		x"50",	--2264
		x"00",	--2265
		x"41",	--2266
		x"12",	--2267
		x"d9",	--2268
		x"41",	--2269
		x"00",	--2270
		x"93",	--2271
		x"28",	--2272
		x"41",	--2273
		x"00",	--2274
		x"93",	--2275
		x"28",	--2276
		x"92",	--2277
		x"24",	--2278
		x"92",	--2279
		x"24",	--2280
		x"93",	--2281
		x"24",	--2282
		x"93",	--2283
		x"24",	--2284
		x"41",	--2285
		x"00",	--2286
		x"41",	--2287
		x"00",	--2288
		x"41",	--2289
		x"00",	--2290
		x"41",	--2291
		x"00",	--2292
		x"40",	--2293
		x"00",	--2294
		x"43",	--2295
		x"43",	--2296
		x"43",	--2297
		x"43",	--2298
		x"43",	--2299
		x"00",	--2300
		x"43",	--2301
		x"00",	--2302
		x"43",	--2303
		x"43",	--2304
		x"4c",	--2305
		x"00",	--2306
		x"3c",	--2307
		x"58",	--2308
		x"69",	--2309
		x"c3",	--2310
		x"10",	--2311
		x"10",	--2312
		x"53",	--2313
		x"00",	--2314
		x"24",	--2315
		x"b3",	--2316
		x"24",	--2317
		x"58",	--2318
		x"69",	--2319
		x"56",	--2320
		x"67",	--2321
		x"43",	--2322
		x"43",	--2323
		x"99",	--2324
		x"28",	--2325
		x"24",	--2326
		x"43",	--2327
		x"43",	--2328
		x"5c",	--2329
		x"6d",	--2330
		x"56",	--2331
		x"67",	--2332
		x"93",	--2333
		x"37",	--2334
		x"d3",	--2335
		x"d3",	--2336
		x"3f",	--2337
		x"98",	--2338
		x"2b",	--2339
		x"3f",	--2340
		x"4a",	--2341
		x"00",	--2342
		x"4b",	--2343
		x"00",	--2344
		x"4f",	--2345
		x"41",	--2346
		x"00",	--2347
		x"51",	--2348
		x"00",	--2349
		x"4a",	--2350
		x"53",	--2351
		x"46",	--2352
		x"00",	--2353
		x"43",	--2354
		x"91",	--2355
		x"00",	--2356
		x"00",	--2357
		x"24",	--2358
		x"4d",	--2359
		x"00",	--2360
		x"93",	--2361
		x"38",	--2362
		x"90",	--2363
		x"40",	--2364
		x"2c",	--2365
		x"41",	--2366
		x"00",	--2367
		x"53",	--2368
		x"41",	--2369
		x"00",	--2370
		x"41",	--2371
		x"00",	--2372
		x"4d",	--2373
		x"5e",	--2374
		x"6f",	--2375
		x"93",	--2376
		x"38",	--2377
		x"5a",	--2378
		x"6b",	--2379
		x"53",	--2380
		x"90",	--2381
		x"40",	--2382
		x"2b",	--2383
		x"4a",	--2384
		x"00",	--2385
		x"4b",	--2386
		x"00",	--2387
		x"4c",	--2388
		x"00",	--2389
		x"4e",	--2390
		x"4f",	--2391
		x"f0",	--2392
		x"00",	--2393
		x"f3",	--2394
		x"90",	--2395
		x"00",	--2396
		x"24",	--2397
		x"4e",	--2398
		x"00",	--2399
		x"4f",	--2400
		x"00",	--2401
		x"40",	--2402
		x"00",	--2403
		x"00",	--2404
		x"41",	--2405
		x"52",	--2406
		x"12",	--2407
		x"d7",	--2408
		x"50",	--2409
		x"00",	--2410
		x"41",	--2411
		x"41",	--2412
		x"41",	--2413
		x"41",	--2414
		x"41",	--2415
		x"41",	--2416
		x"41",	--2417
		x"41",	--2418
		x"41",	--2419
		x"d3",	--2420
		x"d3",	--2421
		x"3f",	--2422
		x"50",	--2423
		x"00",	--2424
		x"4a",	--2425
		x"b3",	--2426
		x"24",	--2427
		x"41",	--2428
		x"00",	--2429
		x"41",	--2430
		x"00",	--2431
		x"c3",	--2432
		x"10",	--2433
		x"10",	--2434
		x"4c",	--2435
		x"4d",	--2436
		x"d3",	--2437
		x"d0",	--2438
		x"80",	--2439
		x"46",	--2440
		x"00",	--2441
		x"47",	--2442
		x"00",	--2443
		x"c3",	--2444
		x"10",	--2445
		x"10",	--2446
		x"53",	--2447
		x"93",	--2448
		x"3b",	--2449
		x"48",	--2450
		x"00",	--2451
		x"3f",	--2452
		x"93",	--2453
		x"24",	--2454
		x"43",	--2455
		x"91",	--2456
		x"00",	--2457
		x"00",	--2458
		x"24",	--2459
		x"4f",	--2460
		x"00",	--2461
		x"41",	--2462
		x"50",	--2463
		x"00",	--2464
		x"3f",	--2465
		x"93",	--2466
		x"23",	--2467
		x"4e",	--2468
		x"4f",	--2469
		x"f0",	--2470
		x"00",	--2471
		x"f3",	--2472
		x"93",	--2473
		x"23",	--2474
		x"93",	--2475
		x"23",	--2476
		x"93",	--2477
		x"00",	--2478
		x"20",	--2479
		x"93",	--2480
		x"00",	--2481
		x"27",	--2482
		x"50",	--2483
		x"00",	--2484
		x"63",	--2485
		x"f0",	--2486
		x"ff",	--2487
		x"f3",	--2488
		x"3f",	--2489
		x"43",	--2490
		x"3f",	--2491
		x"43",	--2492
		x"3f",	--2493
		x"43",	--2494
		x"91",	--2495
		x"00",	--2496
		x"00",	--2497
		x"24",	--2498
		x"4f",	--2499
		x"00",	--2500
		x"41",	--2501
		x"50",	--2502
		x"00",	--2503
		x"3f",	--2504
		x"43",	--2505
		x"3f",	--2506
		x"93",	--2507
		x"23",	--2508
		x"40",	--2509
		x"e8",	--2510
		x"3f",	--2511
		x"12",	--2512
		x"12",	--2513
		x"12",	--2514
		x"12",	--2515
		x"12",	--2516
		x"50",	--2517
		x"ff",	--2518
		x"4e",	--2519
		x"00",	--2520
		x"4f",	--2521
		x"00",	--2522
		x"4c",	--2523
		x"00",	--2524
		x"4d",	--2525
		x"00",	--2526
		x"41",	--2527
		x"50",	--2528
		x"00",	--2529
		x"41",	--2530
		x"52",	--2531
		x"12",	--2532
		x"d9",	--2533
		x"41",	--2534
		x"52",	--2535
		x"41",	--2536
		x"12",	--2537
		x"d9",	--2538
		x"41",	--2539
		x"00",	--2540
		x"93",	--2541
		x"28",	--2542
		x"41",	--2543
		x"00",	--2544
		x"93",	--2545
		x"28",	--2546
		x"e1",	--2547
		x"00",	--2548
		x"00",	--2549
		x"92",	--2550
		x"24",	--2551
		x"93",	--2552
		x"24",	--2553
		x"92",	--2554
		x"24",	--2555
		x"93",	--2556
		x"24",	--2557
		x"41",	--2558
		x"00",	--2559
		x"81",	--2560
		x"00",	--2561
		x"4d",	--2562
		x"00",	--2563
		x"41",	--2564
		x"00",	--2565
		x"41",	--2566
		x"00",	--2567
		x"41",	--2568
		x"00",	--2569
		x"41",	--2570
		x"00",	--2571
		x"99",	--2572
		x"2c",	--2573
		x"5e",	--2574
		x"6f",	--2575
		x"53",	--2576
		x"4d",	--2577
		x"00",	--2578
		x"40",	--2579
		x"00",	--2580
		x"43",	--2581
		x"40",	--2582
		x"40",	--2583
		x"43",	--2584
		x"43",	--2585
		x"3c",	--2586
		x"dc",	--2587
		x"dd",	--2588
		x"88",	--2589
		x"79",	--2590
		x"c3",	--2591
		x"10",	--2592
		x"10",	--2593
		x"5e",	--2594
		x"6f",	--2595
		x"53",	--2596
		x"24",	--2597
		x"99",	--2598
		x"2b",	--2599
		x"23",	--2600
		x"98",	--2601
		x"2b",	--2602
		x"3f",	--2603
		x"9f",	--2604
		x"2b",	--2605
		x"98",	--2606
		x"2f",	--2607
		x"3f",	--2608
		x"4a",	--2609
		x"4b",	--2610
		x"f0",	--2611
		x"00",	--2612
		x"f3",	--2613
		x"90",	--2614
		x"00",	--2615
		x"24",	--2616
		x"4a",	--2617
		x"00",	--2618
		x"4b",	--2619
		x"00",	--2620
		x"41",	--2621
		x"50",	--2622
		x"00",	--2623
		x"12",	--2624
		x"d7",	--2625
		x"50",	--2626
		x"00",	--2627
		x"41",	--2628
		x"41",	--2629
		x"41",	--2630
		x"41",	--2631
		x"41",	--2632
		x"41",	--2633
		x"42",	--2634
		x"00",	--2635
		x"41",	--2636
		x"50",	--2637
		x"00",	--2638
		x"3f",	--2639
		x"9e",	--2640
		x"23",	--2641
		x"40",	--2642
		x"e8",	--2643
		x"3f",	--2644
		x"93",	--2645
		x"23",	--2646
		x"4a",	--2647
		x"4b",	--2648
		x"f0",	--2649
		x"00",	--2650
		x"f3",	--2651
		x"93",	--2652
		x"23",	--2653
		x"93",	--2654
		x"23",	--2655
		x"93",	--2656
		x"20",	--2657
		x"93",	--2658
		x"27",	--2659
		x"50",	--2660
		x"00",	--2661
		x"63",	--2662
		x"f0",	--2663
		x"ff",	--2664
		x"f3",	--2665
		x"3f",	--2666
		x"43",	--2667
		x"00",	--2668
		x"43",	--2669
		x"00",	--2670
		x"43",	--2671
		x"00",	--2672
		x"41",	--2673
		x"50",	--2674
		x"00",	--2675
		x"3f",	--2676
		x"41",	--2677
		x"52",	--2678
		x"3f",	--2679
		x"50",	--2680
		x"ff",	--2681
		x"4e",	--2682
		x"00",	--2683
		x"4f",	--2684
		x"00",	--2685
		x"4c",	--2686
		x"00",	--2687
		x"4d",	--2688
		x"00",	--2689
		x"41",	--2690
		x"50",	--2691
		x"00",	--2692
		x"41",	--2693
		x"52",	--2694
		x"12",	--2695
		x"d9",	--2696
		x"41",	--2697
		x"52",	--2698
		x"41",	--2699
		x"12",	--2700
		x"d9",	--2701
		x"93",	--2702
		x"00",	--2703
		x"28",	--2704
		x"93",	--2705
		x"00",	--2706
		x"28",	--2707
		x"41",	--2708
		x"52",	--2709
		x"41",	--2710
		x"50",	--2711
		x"00",	--2712
		x"12",	--2713
		x"da",	--2714
		x"50",	--2715
		x"00",	--2716
		x"41",	--2717
		x"43",	--2718
		x"3f",	--2719
		x"50",	--2720
		x"ff",	--2721
		x"4e",	--2722
		x"00",	--2723
		x"4f",	--2724
		x"00",	--2725
		x"41",	--2726
		x"52",	--2727
		x"41",	--2728
		x"12",	--2729
		x"d9",	--2730
		x"41",	--2731
		x"00",	--2732
		x"93",	--2733
		x"24",	--2734
		x"28",	--2735
		x"92",	--2736
		x"24",	--2737
		x"41",	--2738
		x"00",	--2739
		x"93",	--2740
		x"38",	--2741
		x"90",	--2742
		x"00",	--2743
		x"38",	--2744
		x"93",	--2745
		x"00",	--2746
		x"20",	--2747
		x"43",	--2748
		x"40",	--2749
		x"7f",	--2750
		x"50",	--2751
		x"00",	--2752
		x"41",	--2753
		x"41",	--2754
		x"00",	--2755
		x"41",	--2756
		x"00",	--2757
		x"40",	--2758
		x"00",	--2759
		x"8d",	--2760
		x"4c",	--2761
		x"f0",	--2762
		x"00",	--2763
		x"20",	--2764
		x"93",	--2765
		x"00",	--2766
		x"27",	--2767
		x"e3",	--2768
		x"e3",	--2769
		x"53",	--2770
		x"63",	--2771
		x"50",	--2772
		x"00",	--2773
		x"41",	--2774
		x"43",	--2775
		x"43",	--2776
		x"50",	--2777
		x"00",	--2778
		x"41",	--2779
		x"c3",	--2780
		x"10",	--2781
		x"10",	--2782
		x"53",	--2783
		x"23",	--2784
		x"3f",	--2785
		x"43",	--2786
		x"40",	--2787
		x"80",	--2788
		x"50",	--2789
		x"00",	--2790
		x"41",	--2791
		x"12",	--2792
		x"12",	--2793
		x"12",	--2794
		x"12",	--2795
		x"82",	--2796
		x"4e",	--2797
		x"4f",	--2798
		x"43",	--2799
		x"00",	--2800
		x"93",	--2801
		x"20",	--2802
		x"93",	--2803
		x"20",	--2804
		x"43",	--2805
		x"00",	--2806
		x"41",	--2807
		x"12",	--2808
		x"d7",	--2809
		x"52",	--2810
		x"41",	--2811
		x"41",	--2812
		x"41",	--2813
		x"41",	--2814
		x"41",	--2815
		x"40",	--2816
		x"00",	--2817
		x"00",	--2818
		x"40",	--2819
		x"00",	--2820
		x"00",	--2821
		x"4a",	--2822
		x"00",	--2823
		x"4b",	--2824
		x"00",	--2825
		x"4a",	--2826
		x"4b",	--2827
		x"12",	--2828
		x"d6",	--2829
		x"53",	--2830
		x"93",	--2831
		x"38",	--2832
		x"27",	--2833
		x"4a",	--2834
		x"00",	--2835
		x"4b",	--2836
		x"00",	--2837
		x"4f",	--2838
		x"f0",	--2839
		x"00",	--2840
		x"20",	--2841
		x"40",	--2842
		x"00",	--2843
		x"8f",	--2844
		x"4e",	--2845
		x"00",	--2846
		x"3f",	--2847
		x"51",	--2848
		x"00",	--2849
		x"00",	--2850
		x"61",	--2851
		x"00",	--2852
		x"00",	--2853
		x"53",	--2854
		x"23",	--2855
		x"3f",	--2856
		x"4f",	--2857
		x"e3",	--2858
		x"53",	--2859
		x"43",	--2860
		x"43",	--2861
		x"4e",	--2862
		x"f0",	--2863
		x"00",	--2864
		x"24",	--2865
		x"5c",	--2866
		x"6d",	--2867
		x"53",	--2868
		x"23",	--2869
		x"53",	--2870
		x"63",	--2871
		x"fa",	--2872
		x"fb",	--2873
		x"43",	--2874
		x"43",	--2875
		x"93",	--2876
		x"20",	--2877
		x"93",	--2878
		x"20",	--2879
		x"43",	--2880
		x"43",	--2881
		x"f0",	--2882
		x"00",	--2883
		x"20",	--2884
		x"48",	--2885
		x"49",	--2886
		x"da",	--2887
		x"db",	--2888
		x"4d",	--2889
		x"00",	--2890
		x"4e",	--2891
		x"00",	--2892
		x"40",	--2893
		x"00",	--2894
		x"8f",	--2895
		x"4e",	--2896
		x"00",	--2897
		x"3f",	--2898
		x"c3",	--2899
		x"10",	--2900
		x"10",	--2901
		x"53",	--2902
		x"23",	--2903
		x"3f",	--2904
		x"12",	--2905
		x"12",	--2906
		x"12",	--2907
		x"93",	--2908
		x"2c",	--2909
		x"90",	--2910
		x"01",	--2911
		x"28",	--2912
		x"40",	--2913
		x"00",	--2914
		x"43",	--2915
		x"42",	--2916
		x"4e",	--2917
		x"4f",	--2918
		x"49",	--2919
		x"93",	--2920
		x"20",	--2921
		x"50",	--2922
		x"e8",	--2923
		x"4c",	--2924
		x"43",	--2925
		x"8e",	--2926
		x"7f",	--2927
		x"4a",	--2928
		x"41",	--2929
		x"41",	--2930
		x"41",	--2931
		x"41",	--2932
		x"90",	--2933
		x"01",	--2934
		x"28",	--2935
		x"42",	--2936
		x"43",	--2937
		x"40",	--2938
		x"00",	--2939
		x"4e",	--2940
		x"4f",	--2941
		x"49",	--2942
		x"93",	--2943
		x"27",	--2944
		x"c3",	--2945
		x"10",	--2946
		x"10",	--2947
		x"53",	--2948
		x"23",	--2949
		x"3f",	--2950
		x"40",	--2951
		x"00",	--2952
		x"43",	--2953
		x"40",	--2954
		x"00",	--2955
		x"3f",	--2956
		x"40",	--2957
		x"00",	--2958
		x"43",	--2959
		x"43",	--2960
		x"3f",	--2961
		x"12",	--2962
		x"12",	--2963
		x"12",	--2964
		x"12",	--2965
		x"12",	--2966
		x"4f",	--2967
		x"4f",	--2968
		x"00",	--2969
		x"4f",	--2970
		x"00",	--2971
		x"4d",	--2972
		x"00",	--2973
		x"4d",	--2974
		x"93",	--2975
		x"28",	--2976
		x"92",	--2977
		x"24",	--2978
		x"93",	--2979
		x"24",	--2980
		x"93",	--2981
		x"24",	--2982
		x"4d",	--2983
		x"00",	--2984
		x"90",	--2985
		x"ff",	--2986
		x"38",	--2987
		x"90",	--2988
		x"00",	--2989
		x"34",	--2990
		x"4e",	--2991
		x"4f",	--2992
		x"f0",	--2993
		x"00",	--2994
		x"f3",	--2995
		x"90",	--2996
		x"00",	--2997
		x"24",	--2998
		x"50",	--2999
		x"00",	--3000
		x"63",	--3001
		x"93",	--3002
		x"38",	--3003
		x"4b",	--3004
		x"50",	--3005
		x"00",	--3006
		x"c3",	--3007
		x"10",	--3008
		x"10",	--3009
		x"c3",	--3010
		x"10",	--3011
		x"10",	--3012
		x"c3",	--3013
		x"10",	--3014
		x"10",	--3015
		x"c3",	--3016
		x"10",	--3017
		x"10",	--3018
		x"c3",	--3019
		x"10",	--3020
		x"10",	--3021
		x"c3",	--3022
		x"10",	--3023
		x"10",	--3024
		x"c3",	--3025
		x"10",	--3026
		x"10",	--3027
		x"f3",	--3028
		x"f0",	--3029
		x"00",	--3030
		x"4d",	--3031
		x"3c",	--3032
		x"93",	--3033
		x"23",	--3034
		x"43",	--3035
		x"43",	--3036
		x"43",	--3037
		x"4d",	--3038
		x"5d",	--3039
		x"5d",	--3040
		x"5d",	--3041
		x"5d",	--3042
		x"5d",	--3043
		x"5d",	--3044
		x"5d",	--3045
		x"4f",	--3046
		x"f0",	--3047
		x"00",	--3048
		x"dd",	--3049
		x"4a",	--3050
		x"11",	--3051
		x"43",	--3052
		x"10",	--3053
		x"4c",	--3054
		x"df",	--3055
		x"4d",	--3056
		x"41",	--3057
		x"41",	--3058
		x"41",	--3059
		x"41",	--3060
		x"41",	--3061
		x"41",	--3062
		x"93",	--3063
		x"23",	--3064
		x"4e",	--3065
		x"4f",	--3066
		x"f0",	--3067
		x"00",	--3068
		x"f3",	--3069
		x"93",	--3070
		x"20",	--3071
		x"93",	--3072
		x"27",	--3073
		x"50",	--3074
		x"00",	--3075
		x"63",	--3076
		x"3f",	--3077
		x"c3",	--3078
		x"10",	--3079
		x"10",	--3080
		x"4b",	--3081
		x"50",	--3082
		x"00",	--3083
		x"3f",	--3084
		x"43",	--3085
		x"43",	--3086
		x"43",	--3087
		x"3f",	--3088
		x"d3",	--3089
		x"d0",	--3090
		x"00",	--3091
		x"f3",	--3092
		x"f0",	--3093
		x"00",	--3094
		x"43",	--3095
		x"3f",	--3096
		x"40",	--3097
		x"ff",	--3098
		x"8b",	--3099
		x"90",	--3100
		x"00",	--3101
		x"34",	--3102
		x"4e",	--3103
		x"4f",	--3104
		x"47",	--3105
		x"f0",	--3106
		x"00",	--3107
		x"24",	--3108
		x"c3",	--3109
		x"10",	--3110
		x"10",	--3111
		x"53",	--3112
		x"23",	--3113
		x"43",	--3114
		x"43",	--3115
		x"f0",	--3116
		x"00",	--3117
		x"24",	--3118
		x"58",	--3119
		x"69",	--3120
		x"53",	--3121
		x"23",	--3122
		x"53",	--3123
		x"63",	--3124
		x"fe",	--3125
		x"ff",	--3126
		x"43",	--3127
		x"43",	--3128
		x"93",	--3129
		x"20",	--3130
		x"93",	--3131
		x"20",	--3132
		x"43",	--3133
		x"43",	--3134
		x"4e",	--3135
		x"4f",	--3136
		x"dc",	--3137
		x"dd",	--3138
		x"48",	--3139
		x"49",	--3140
		x"f0",	--3141
		x"00",	--3142
		x"f3",	--3143
		x"90",	--3144
		x"00",	--3145
		x"24",	--3146
		x"50",	--3147
		x"00",	--3148
		x"63",	--3149
		x"48",	--3150
		x"49",	--3151
		x"c3",	--3152
		x"10",	--3153
		x"10",	--3154
		x"c3",	--3155
		x"10",	--3156
		x"10",	--3157
		x"c3",	--3158
		x"10",	--3159
		x"10",	--3160
		x"c3",	--3161
		x"10",	--3162
		x"10",	--3163
		x"c3",	--3164
		x"10",	--3165
		x"10",	--3166
		x"c3",	--3167
		x"10",	--3168
		x"10",	--3169
		x"c3",	--3170
		x"10",	--3171
		x"10",	--3172
		x"f3",	--3173
		x"f0",	--3174
		x"00",	--3175
		x"43",	--3176
		x"90",	--3177
		x"40",	--3178
		x"2f",	--3179
		x"43",	--3180
		x"3f",	--3181
		x"43",	--3182
		x"43",	--3183
		x"3f",	--3184
		x"93",	--3185
		x"23",	--3186
		x"48",	--3187
		x"49",	--3188
		x"f0",	--3189
		x"00",	--3190
		x"f3",	--3191
		x"93",	--3192
		x"24",	--3193
		x"50",	--3194
		x"00",	--3195
		x"63",	--3196
		x"3f",	--3197
		x"93",	--3198
		x"27",	--3199
		x"3f",	--3200
		x"12",	--3201
		x"12",	--3202
		x"4f",	--3203
		x"4f",	--3204
		x"00",	--3205
		x"f0",	--3206
		x"00",	--3207
		x"4f",	--3208
		x"00",	--3209
		x"c3",	--3210
		x"10",	--3211
		x"c3",	--3212
		x"10",	--3213
		x"c3",	--3214
		x"10",	--3215
		x"c3",	--3216
		x"10",	--3217
		x"c3",	--3218
		x"10",	--3219
		x"c3",	--3220
		x"10",	--3221
		x"c3",	--3222
		x"10",	--3223
		x"4d",	--3224
		x"4f",	--3225
		x"00",	--3226
		x"b0",	--3227
		x"00",	--3228
		x"43",	--3229
		x"6f",	--3230
		x"4f",	--3231
		x"00",	--3232
		x"93",	--3233
		x"20",	--3234
		x"93",	--3235
		x"24",	--3236
		x"40",	--3237
		x"ff",	--3238
		x"00",	--3239
		x"4a",	--3240
		x"4b",	--3241
		x"5c",	--3242
		x"6d",	--3243
		x"5c",	--3244
		x"6d",	--3245
		x"5c",	--3246
		x"6d",	--3247
		x"5c",	--3248
		x"6d",	--3249
		x"5c",	--3250
		x"6d",	--3251
		x"5c",	--3252
		x"6d",	--3253
		x"5c",	--3254
		x"6d",	--3255
		x"40",	--3256
		x"00",	--3257
		x"00",	--3258
		x"90",	--3259
		x"40",	--3260
		x"2c",	--3261
		x"40",	--3262
		x"ff",	--3263
		x"5c",	--3264
		x"6d",	--3265
		x"4f",	--3266
		x"53",	--3267
		x"90",	--3268
		x"40",	--3269
		x"2b",	--3270
		x"4a",	--3271
		x"00",	--3272
		x"4c",	--3273
		x"00",	--3274
		x"4d",	--3275
		x"00",	--3276
		x"41",	--3277
		x"41",	--3278
		x"41",	--3279
		x"90",	--3280
		x"00",	--3281
		x"24",	--3282
		x"50",	--3283
		x"ff",	--3284
		x"4d",	--3285
		x"00",	--3286
		x"40",	--3287
		x"00",	--3288
		x"00",	--3289
		x"4a",	--3290
		x"4b",	--3291
		x"5c",	--3292
		x"6d",	--3293
		x"5c",	--3294
		x"6d",	--3295
		x"5c",	--3296
		x"6d",	--3297
		x"5c",	--3298
		x"6d",	--3299
		x"5c",	--3300
		x"6d",	--3301
		x"5c",	--3302
		x"6d",	--3303
		x"5c",	--3304
		x"6d",	--3305
		x"4c",	--3306
		x"4d",	--3307
		x"d3",	--3308
		x"d0",	--3309
		x"40",	--3310
		x"4a",	--3311
		x"00",	--3312
		x"4b",	--3313
		x"00",	--3314
		x"41",	--3315
		x"41",	--3316
		x"41",	--3317
		x"93",	--3318
		x"23",	--3319
		x"43",	--3320
		x"00",	--3321
		x"41",	--3322
		x"41",	--3323
		x"41",	--3324
		x"93",	--3325
		x"24",	--3326
		x"4a",	--3327
		x"4b",	--3328
		x"f3",	--3329
		x"f0",	--3330
		x"00",	--3331
		x"93",	--3332
		x"20",	--3333
		x"93",	--3334
		x"24",	--3335
		x"43",	--3336
		x"00",	--3337
		x"3f",	--3338
		x"93",	--3339
		x"23",	--3340
		x"42",	--3341
		x"00",	--3342
		x"3f",	--3343
		x"43",	--3344
		x"00",	--3345
		x"3f",	--3346
		x"12",	--3347
		x"4f",	--3348
		x"93",	--3349
		x"28",	--3350
		x"4e",	--3351
		x"93",	--3352
		x"28",	--3353
		x"92",	--3354
		x"24",	--3355
		x"92",	--3356
		x"24",	--3357
		x"93",	--3358
		x"24",	--3359
		x"93",	--3360
		x"24",	--3361
		x"4f",	--3362
		x"00",	--3363
		x"9e",	--3364
		x"00",	--3365
		x"24",	--3366
		x"93",	--3367
		x"20",	--3368
		x"43",	--3369
		x"4e",	--3370
		x"41",	--3371
		x"41",	--3372
		x"93",	--3373
		x"24",	--3374
		x"93",	--3375
		x"00",	--3376
		x"23",	--3377
		x"43",	--3378
		x"4e",	--3379
		x"41",	--3380
		x"41",	--3381
		x"93",	--3382
		x"00",	--3383
		x"27",	--3384
		x"43",	--3385
		x"3f",	--3386
		x"4f",	--3387
		x"00",	--3388
		x"4e",	--3389
		x"00",	--3390
		x"9b",	--3391
		x"3b",	--3392
		x"9c",	--3393
		x"38",	--3394
		x"4f",	--3395
		x"00",	--3396
		x"4f",	--3397
		x"00",	--3398
		x"4e",	--3399
		x"00",	--3400
		x"4e",	--3401
		x"00",	--3402
		x"9f",	--3403
		x"2b",	--3404
		x"9e",	--3405
		x"28",	--3406
		x"9b",	--3407
		x"2b",	--3408
		x"9e",	--3409
		x"28",	--3410
		x"9f",	--3411
		x"28",	--3412
		x"9c",	--3413
		x"28",	--3414
		x"43",	--3415
		x"3f",	--3416
		x"93",	--3417
		x"23",	--3418
		x"43",	--3419
		x"3f",	--3420
		x"92",	--3421
		x"23",	--3422
		x"4e",	--3423
		x"00",	--3424
		x"4f",	--3425
		x"00",	--3426
		x"8f",	--3427
		x"3f",	--3428
		x"42",	--3429
		x"02",	--3430
		x"93",	--3431
		x"38",	--3432
		x"42",	--3433
		x"02",	--3434
		x"4f",	--3435
		x"00",	--3436
		x"53",	--3437
		x"4d",	--3438
		x"02",	--3439
		x"53",	--3440
		x"4e",	--3441
		x"02",	--3442
		x"41",	--3443
		x"43",	--3444
		x"41",	--3445
		x"12",	--3446
		x"12",	--3447
		x"83",	--3448
		x"4e",	--3449
		x"00",	--3450
		x"42",	--3451
		x"02",	--3452
		x"42",	--3453
		x"02",	--3454
		x"4e",	--3455
		x"4f",	--3456
		x"40",	--3457
		x"da",	--3458
		x"12",	--3459
		x"dd",	--3460
		x"9b",	--3461
		x"38",	--3462
		x"4a",	--3463
		x"5b",	--3464
		x"43",	--3465
		x"ff",	--3466
		x"3c",	--3467
		x"42",	--3468
		x"02",	--3469
		x"43",	--3470
		x"00",	--3471
		x"53",	--3472
		x"41",	--3473
		x"41",	--3474
		x"41",	--3475
		x"41",	--3476
		x"00",	--3477
		x"02",	--3478
		x"40",	--3479
		x"7f",	--3480
		x"02",	--3481
		x"41",	--3482
		x"50",	--3483
		x"00",	--3484
		x"41",	--3485
		x"00",	--3486
		x"12",	--3487
		x"da",	--3488
		x"41",	--3489
		x"41",	--3490
		x"00",	--3491
		x"02",	--3492
		x"41",	--3493
		x"00",	--3494
		x"02",	--3495
		x"41",	--3496
		x"52",	--3497
		x"41",	--3498
		x"00",	--3499
		x"12",	--3500
		x"da",	--3501
		x"41",	--3502
		x"4e",	--3503
		x"4f",	--3504
		x"02",	--3505
		x"40",	--3506
		x"7f",	--3507
		x"02",	--3508
		x"4d",	--3509
		x"4c",	--3510
		x"12",	--3511
		x"da",	--3512
		x"41",	--3513
		x"4f",	--3514
		x"02",	--3515
		x"4e",	--3516
		x"02",	--3517
		x"4c",	--3518
		x"4d",	--3519
		x"12",	--3520
		x"da",	--3521
		x"41",	--3522
		x"12",	--3523
		x"12",	--3524
		x"12",	--3525
		x"12",	--3526
		x"12",	--3527
		x"12",	--3528
		x"12",	--3529
		x"12",	--3530
		x"82",	--3531
		x"4f",	--3532
		x"4e",	--3533
		x"00",	--3534
		x"4d",	--3535
		x"41",	--3536
		x"00",	--3537
		x"41",	--3538
		x"00",	--3539
		x"4d",	--3540
		x"4d",	--3541
		x"10",	--3542
		x"44",	--3543
		x"4f",	--3544
		x"b0",	--3545
		x"00",	--3546
		x"24",	--3547
		x"40",	--3548
		x"00",	--3549
		x"00",	--3550
		x"4f",	--3551
		x"10",	--3552
		x"f3",	--3553
		x"24",	--3554
		x"40",	--3555
		x"00",	--3556
		x"3c",	--3557
		x"40",	--3558
		x"00",	--3559
		x"4e",	--3560
		x"00",	--3561
		x"41",	--3562
		x"53",	--3563
		x"3c",	--3564
		x"f0",	--3565
		x"00",	--3566
		x"24",	--3567
		x"40",	--3568
		x"00",	--3569
		x"00",	--3570
		x"3c",	--3571
		x"93",	--3572
		x"24",	--3573
		x"4d",	--3574
		x"00",	--3575
		x"41",	--3576
		x"53",	--3577
		x"3c",	--3578
		x"41",	--3579
		x"4c",	--3580
		x"10",	--3581
		x"11",	--3582
		x"10",	--3583
		x"11",	--3584
		x"4c",	--3585
		x"41",	--3586
		x"41",	--3587
		x"10",	--3588
		x"11",	--3589
		x"10",	--3590
		x"11",	--3591
		x"4c",	--3592
		x"86",	--3593
		x"77",	--3594
		x"4f",	--3595
		x"10",	--3596
		x"4e",	--3597
		x"00",	--3598
		x"f2",	--3599
		x"24",	--3600
		x"45",	--3601
		x"3c",	--3602
		x"43",	--3603
		x"4f",	--3604
		x"b0",	--3605
		x"00",	--3606
		x"20",	--3607
		x"41",	--3608
		x"00",	--3609
		x"53",	--3610
		x"53",	--3611
		x"93",	--3612
		x"00",	--3613
		x"23",	--3614
		x"81",	--3615
		x"00",	--3616
		x"9a",	--3617
		x"28",	--3618
		x"8a",	--3619
		x"3c",	--3620
		x"43",	--3621
		x"b3",	--3622
		x"00",	--3623
		x"24",	--3624
		x"95",	--3625
		x"28",	--3626
		x"85",	--3627
		x"3c",	--3628
		x"43",	--3629
		x"4d",	--3630
		x"9d",	--3631
		x"2c",	--3632
		x"47",	--3633
		x"93",	--3634
		x"38",	--3635
		x"40",	--3636
		x"00",	--3637
		x"00",	--3638
		x"43",	--3639
		x"43",	--3640
		x"3c",	--3641
		x"41",	--3642
		x"56",	--3643
		x"4f",	--3644
		x"11",	--3645
		x"53",	--3646
		x"12",	--3647
		x"3c",	--3648
		x"43",	--3649
		x"9a",	--3650
		x"3b",	--3651
		x"4a",	--3652
		x"40",	--3653
		x"00",	--3654
		x"00",	--3655
		x"8b",	--3656
		x"3c",	--3657
		x"41",	--3658
		x"00",	--3659
		x"11",	--3660
		x"12",	--3661
		x"53",	--3662
		x"45",	--3663
		x"5b",	--3664
		x"99",	--3665
		x"2b",	--3666
		x"3c",	--3667
		x"43",	--3668
		x"43",	--3669
		x"3c",	--3670
		x"53",	--3671
		x"41",	--3672
		x"56",	--3673
		x"4f",	--3674
		x"11",	--3675
		x"53",	--3676
		x"12",	--3677
		x"9a",	--3678
		x"3b",	--3679
		x"b3",	--3680
		x"00",	--3681
		x"24",	--3682
		x"44",	--3683
		x"3c",	--3684
		x"41",	--3685
		x"00",	--3686
		x"8b",	--3687
		x"3c",	--3688
		x"40",	--3689
		x"00",	--3690
		x"12",	--3691
		x"53",	--3692
		x"93",	--3693
		x"23",	--3694
		x"44",	--3695
		x"54",	--3696
		x"3f",	--3697
		x"53",	--3698
		x"11",	--3699
		x"12",	--3700
		x"53",	--3701
		x"4a",	--3702
		x"5b",	--3703
		x"4f",	--3704
		x"93",	--3705
		x"24",	--3706
		x"93",	--3707
		x"23",	--3708
		x"3c",	--3709
		x"40",	--3710
		x"00",	--3711
		x"12",	--3712
		x"53",	--3713
		x"99",	--3714
		x"2b",	--3715
		x"4b",	--3716
		x"52",	--3717
		x"41",	--3718
		x"41",	--3719
		x"41",	--3720
		x"41",	--3721
		x"41",	--3722
		x"41",	--3723
		x"41",	--3724
		x"41",	--3725
		x"41",	--3726
		x"12",	--3727
		x"12",	--3728
		x"12",	--3729
		x"12",	--3730
		x"12",	--3731
		x"12",	--3732
		x"12",	--3733
		x"12",	--3734
		x"50",	--3735
		x"ff",	--3736
		x"4f",	--3737
		x"00",	--3738
		x"4e",	--3739
		x"4d",	--3740
		x"4e",	--3741
		x"00",	--3742
		x"43",	--3743
		x"00",	--3744
		x"43",	--3745
		x"00",	--3746
		x"43",	--3747
		x"00",	--3748
		x"43",	--3749
		x"00",	--3750
		x"43",	--3751
		x"00",	--3752
		x"43",	--3753
		x"00",	--3754
		x"43",	--3755
		x"43",	--3756
		x"00",	--3757
		x"41",	--3758
		x"50",	--3759
		x"00",	--3760
		x"4e",	--3761
		x"00",	--3762
		x"40",	--3763
		x"e3",	--3764
		x"46",	--3765
		x"53",	--3766
		x"4f",	--3767
		x"00",	--3768
		x"93",	--3769
		x"20",	--3770
		x"90",	--3771
		x"00",	--3772
		x"20",	--3773
		x"43",	--3774
		x"00",	--3775
		x"43",	--3776
		x"00",	--3777
		x"46",	--3778
		x"00",	--3779
		x"43",	--3780
		x"00",	--3781
		x"43",	--3782
		x"00",	--3783
		x"43",	--3784
		x"00",	--3785
		x"43",	--3786
		x"00",	--3787
		x"43",	--3788
		x"00",	--3789
		x"40",	--3790
		x"e3",	--3791
		x"47",	--3792
		x"11",	--3793
		x"4e",	--3794
		x"12",	--3795
		x"00",	--3796
		x"53",	--3797
		x"00",	--3798
		x"40",	--3799
		x"e3",	--3800
		x"90",	--3801
		x"00",	--3802
		x"24",	--3803
		x"90",	--3804
		x"00",	--3805
		x"34",	--3806
		x"90",	--3807
		x"00",	--3808
		x"24",	--3809
		x"90",	--3810
		x"00",	--3811
		x"34",	--3812
		x"90",	--3813
		x"00",	--3814
		x"24",	--3815
		x"90",	--3816
		x"00",	--3817
		x"34",	--3818
		x"90",	--3819
		x"00",	--3820
		x"24",	--3821
		x"90",	--3822
		x"00",	--3823
		x"27",	--3824
		x"90",	--3825
		x"00",	--3826
		x"20",	--3827
		x"3c",	--3828
		x"90",	--3829
		x"00",	--3830
		x"24",	--3831
		x"90",	--3832
		x"00",	--3833
		x"24",	--3834
		x"90",	--3835
		x"00",	--3836
		x"20",	--3837
		x"3c",	--3838
		x"90",	--3839
		x"00",	--3840
		x"38",	--3841
		x"90",	--3842
		x"00",	--3843
		x"20",	--3844
		x"3c",	--3845
		x"90",	--3846
		x"00",	--3847
		x"24",	--3848
		x"90",	--3849
		x"00",	--3850
		x"34",	--3851
		x"90",	--3852
		x"00",	--3853
		x"24",	--3854
		x"90",	--3855
		x"00",	--3856
		x"24",	--3857
		x"90",	--3858
		x"00",	--3859
		x"20",	--3860
		x"3c",	--3861
		x"90",	--3862
		x"00",	--3863
		x"24",	--3864
		x"90",	--3865
		x"00",	--3866
		x"34",	--3867
		x"90",	--3868
		x"00",	--3869
		x"20",	--3870
		x"3c",	--3871
		x"90",	--3872
		x"00",	--3873
		x"24",	--3874
		x"90",	--3875
		x"00",	--3876
		x"24",	--3877
		x"41",	--3878
		x"00",	--3879
		x"41",	--3880
		x"00",	--3881
		x"89",	--3882
		x"40",	--3883
		x"e3",	--3884
		x"42",	--3885
		x"00",	--3886
		x"3c",	--3887
		x"d2",	--3888
		x"00",	--3889
		x"40",	--3890
		x"e3",	--3891
		x"41",	--3892
		x"f3",	--3893
		x"41",	--3894
		x"24",	--3895
		x"f0",	--3896
		x"ff",	--3897
		x"d3",	--3898
		x"3c",	--3899
		x"d3",	--3900
		x"4e",	--3901
		x"00",	--3902
		x"40",	--3903
		x"e3",	--3904
		x"d0",	--3905
		x"00",	--3906
		x"00",	--3907
		x"40",	--3908
		x"e3",	--3909
		x"40",	--3910
		x"00",	--3911
		x"00",	--3912
		x"40",	--3913
		x"e3",	--3914
		x"90",	--3915
		x"00",	--3916
		x"00",	--3917
		x"20",	--3918
		x"40",	--3919
		x"e3",	--3920
		x"40",	--3921
		x"00",	--3922
		x"00",	--3923
		x"40",	--3924
		x"e3",	--3925
		x"93",	--3926
		x"00",	--3927
		x"24",	--3928
		x"40",	--3929
		x"e3",	--3930
		x"43",	--3931
		x"00",	--3932
		x"40",	--3933
		x"e3",	--3934
		x"45",	--3935
		x"53",	--3936
		x"45",	--3937
		x"93",	--3938
		x"38",	--3939
		x"4a",	--3940
		x"00",	--3941
		x"3c",	--3942
		x"93",	--3943
		x"00",	--3944
		x"24",	--3945
		x"40",	--3946
		x"e3",	--3947
		x"d0",	--3948
		x"00",	--3949
		x"00",	--3950
		x"e3",	--3951
		x"4a",	--3952
		x"00",	--3953
		x"53",	--3954
		x"00",	--3955
		x"4e",	--3956
		x"3c",	--3957
		x"93",	--3958
		x"00",	--3959
		x"20",	--3960
		x"93",	--3961
		x"00",	--3962
		x"20",	--3963
		x"41",	--3964
		x"f0",	--3965
		x"00",	--3966
		x"43",	--3967
		x"24",	--3968
		x"43",	--3969
		x"4e",	--3970
		x"11",	--3971
		x"43",	--3972
		x"10",	--3973
		x"41",	--3974
		x"f0",	--3975
		x"00",	--3976
		x"de",	--3977
		x"4a",	--3978
		x"00",	--3979
		x"40",	--3980
		x"e3",	--3981
		x"41",	--3982
		x"00",	--3983
		x"5a",	--3984
		x"4a",	--3985
		x"5c",	--3986
		x"5c",	--3987
		x"5c",	--3988
		x"4a",	--3989
		x"00",	--3990
		x"50",	--3991
		x"ff",	--3992
		x"00",	--3993
		x"11",	--3994
		x"5e",	--3995
		x"00",	--3996
		x"43",	--3997
		x"00",	--3998
		x"40",	--3999
		x"e3",	--4000
		x"45",	--4001
		x"53",	--4002
		x"45",	--4003
		x"93",	--4004
		x"00",	--4005
		x"20",	--4006
		x"93",	--4007
		x"00",	--4008
		x"27",	--4009
		x"4e",	--4010
		x"00",	--4011
		x"43",	--4012
		x"00",	--4013
		x"41",	--4014
		x"52",	--4015
		x"3c",	--4016
		x"45",	--4017
		x"53",	--4018
		x"45",	--4019
		x"93",	--4020
		x"00",	--4021
		x"24",	--4022
		x"d2",	--4023
		x"00",	--4024
		x"41",	--4025
		x"00",	--4026
		x"4f",	--4027
		x"00",	--4028
		x"3c",	--4029
		x"93",	--4030
		x"00",	--4031
		x"24",	--4032
		x"41",	--4033
		x"00",	--4034
		x"00",	--4035
		x"93",	--4036
		x"20",	--4037
		x"40",	--4038
		x"e9",	--4039
		x"12",	--4040
		x"00",	--4041
		x"12",	--4042
		x"00",	--4043
		x"41",	--4044
		x"00",	--4045
		x"41",	--4046
		x"00",	--4047
		x"12",	--4048
		x"db",	--4049
		x"52",	--4050
		x"5f",	--4051
		x"00",	--4052
		x"47",	--4053
		x"40",	--4054
		x"e3",	--4055
		x"45",	--4056
		x"53",	--4057
		x"45",	--4058
		x"49",	--4059
		x"00",	--4060
		x"43",	--4061
		x"93",	--4062
		x"20",	--4063
		x"43",	--4064
		x"5e",	--4065
		x"5e",	--4066
		x"5e",	--4067
		x"41",	--4068
		x"f0",	--4069
		x"ff",	--4070
		x"de",	--4071
		x"4a",	--4072
		x"00",	--4073
		x"47",	--4074
		x"40",	--4075
		x"00",	--4076
		x"00",	--4077
		x"3c",	--4078
		x"d3",	--4079
		x"00",	--4080
		x"3c",	--4081
		x"d2",	--4082
		x"00",	--4083
		x"40",	--4084
		x"00",	--4085
		x"00",	--4086
		x"3c",	--4087
		x"40",	--4088
		x"00",	--4089
		x"00",	--4090
		x"41",	--4091
		x"b3",	--4092
		x"24",	--4093
		x"45",	--4094
		x"52",	--4095
		x"45",	--4096
		x"45",	--4097
		x"00",	--4098
		x"45",	--4099
		x"00",	--4100
		x"45",	--4101
		x"00",	--4102
		x"48",	--4103
		x"00",	--4104
		x"47",	--4105
		x"00",	--4106
		x"46",	--4107
		x"00",	--4108
		x"4b",	--4109
		x"00",	--4110
		x"43",	--4111
		x"00",	--4112
		x"93",	--4113
		x"20",	--4114
		x"93",	--4115
		x"20",	--4116
		x"93",	--4117
		x"20",	--4118
		x"93",	--4119
		x"24",	--4120
		x"43",	--4121
		x"00",	--4122
		x"5b",	--4123
		x"43",	--4124
		x"6b",	--4125
		x"4b",	--4126
		x"00",	--4127
		x"4c",	--4128
		x"3c",	--4129
		x"f3",	--4130
		x"45",	--4131
		x"24",	--4132
		x"52",	--4133
		x"45",	--4134
		x"45",	--4135
		x"00",	--4136
		x"48",	--4137
		x"00",	--4138
		x"4b",	--4139
		x"00",	--4140
		x"43",	--4141
		x"00",	--4142
		x"93",	--4143
		x"20",	--4144
		x"3c",	--4145
		x"53",	--4146
		x"45",	--4147
		x"4b",	--4148
		x"00",	--4149
		x"43",	--4150
		x"00",	--4151
		x"93",	--4152
		x"24",	--4153
		x"43",	--4154
		x"00",	--4155
		x"5b",	--4156
		x"43",	--4157
		x"6b",	--4158
		x"4b",	--4159
		x"00",	--4160
		x"47",	--4161
		x"b2",	--4162
		x"00",	--4163
		x"24",	--4164
		x"93",	--4165
		x"00",	--4166
		x"20",	--4167
		x"41",	--4168
		x"90",	--4169
		x"00",	--4170
		x"00",	--4171
		x"20",	--4172
		x"d0",	--4173
		x"00",	--4174
		x"3c",	--4175
		x"92",	--4176
		x"00",	--4177
		x"20",	--4178
		x"d0",	--4179
		x"00",	--4180
		x"48",	--4181
		x"00",	--4182
		x"41",	--4183
		x"b2",	--4184
		x"24",	--4185
		x"93",	--4186
		x"00",	--4187
		x"24",	--4188
		x"40",	--4189
		x"00",	--4190
		x"00",	--4191
		x"b3",	--4192
		x"24",	--4193
		x"e3",	--4194
		x"00",	--4195
		x"e3",	--4196
		x"00",	--4197
		x"e3",	--4198
		x"00",	--4199
		x"e3",	--4200
		x"00",	--4201
		x"53",	--4202
		x"00",	--4203
		x"63",	--4204
		x"00",	--4205
		x"63",	--4206
		x"00",	--4207
		x"63",	--4208
		x"00",	--4209
		x"3c",	--4210
		x"b3",	--4211
		x"24",	--4212
		x"41",	--4213
		x"00",	--4214
		x"41",	--4215
		x"00",	--4216
		x"e3",	--4217
		x"e3",	--4218
		x"4a",	--4219
		x"4b",	--4220
		x"53",	--4221
		x"63",	--4222
		x"4e",	--4223
		x"00",	--4224
		x"4f",	--4225
		x"00",	--4226
		x"3c",	--4227
		x"41",	--4228
		x"00",	--4229
		x"e3",	--4230
		x"53",	--4231
		x"4a",	--4232
		x"00",	--4233
		x"43",	--4234
		x"00",	--4235
		x"b3",	--4236
		x"24",	--4237
		x"41",	--4238
		x"00",	--4239
		x"41",	--4240
		x"00",	--4241
		x"00",	--4242
		x"41",	--4243
		x"00",	--4244
		x"41",	--4245
		x"00",	--4246
		x"41",	--4247
		x"50",	--4248
		x"00",	--4249
		x"46",	--4250
		x"41",	--4251
		x"00",	--4252
		x"00",	--4253
		x"41",	--4254
		x"00",	--4255
		x"10",	--4256
		x"11",	--4257
		x"10",	--4258
		x"11",	--4259
		x"4b",	--4260
		x"00",	--4261
		x"4b",	--4262
		x"00",	--4263
		x"4b",	--4264
		x"00",	--4265
		x"12",	--4266
		x"00",	--4267
		x"12",	--4268
		x"00",	--4269
		x"12",	--4270
		x"00",	--4271
		x"12",	--4272
		x"00",	--4273
		x"49",	--4274
		x"41",	--4275
		x"00",	--4276
		x"48",	--4277
		x"44",	--4278
		x"12",	--4279
		x"e5",	--4280
		x"52",	--4281
		x"4c",	--4282
		x"90",	--4283
		x"00",	--4284
		x"34",	--4285
		x"50",	--4286
		x"00",	--4287
		x"4b",	--4288
		x"00",	--4289
		x"3c",	--4290
		x"4c",	--4291
		x"b3",	--4292
		x"00",	--4293
		x"24",	--4294
		x"40",	--4295
		x"00",	--4296
		x"3c",	--4297
		x"40",	--4298
		x"00",	--4299
		x"5b",	--4300
		x"4a",	--4301
		x"00",	--4302
		x"47",	--4303
		x"53",	--4304
		x"12",	--4305
		x"00",	--4306
		x"12",	--4307
		x"00",	--4308
		x"12",	--4309
		x"00",	--4310
		x"12",	--4311
		x"00",	--4312
		x"49",	--4313
		x"41",	--4314
		x"00",	--4315
		x"48",	--4316
		x"44",	--4317
		x"12",	--4318
		x"e5",	--4319
		x"52",	--4320
		x"4c",	--4321
		x"4d",	--4322
		x"00",	--4323
		x"4e",	--4324
		x"4f",	--4325
		x"53",	--4326
		x"93",	--4327
		x"23",	--4328
		x"93",	--4329
		x"23",	--4330
		x"93",	--4331
		x"23",	--4332
		x"93",	--4333
		x"23",	--4334
		x"43",	--4335
		x"00",	--4336
		x"43",	--4337
		x"00",	--4338
		x"43",	--4339
		x"00",	--4340
		x"43",	--4341
		x"00",	--4342
		x"3c",	--4343
		x"b3",	--4344
		x"24",	--4345
		x"41",	--4346
		x"00",	--4347
		x"41",	--4348
		x"00",	--4349
		x"41",	--4350
		x"50",	--4351
		x"00",	--4352
		x"41",	--4353
		x"00",	--4354
		x"10",	--4355
		x"11",	--4356
		x"10",	--4357
		x"11",	--4358
		x"41",	--4359
		x"00",	--4360
		x"49",	--4361
		x"44",	--4362
		x"47",	--4363
		x"12",	--4364
		x"e4",	--4365
		x"4e",	--4366
		x"90",	--4367
		x"00",	--4368
		x"34",	--4369
		x"50",	--4370
		x"00",	--4371
		x"4b",	--4372
		x"00",	--4373
		x"3c",	--4374
		x"4e",	--4375
		x"b3",	--4376
		x"00",	--4377
		x"24",	--4378
		x"40",	--4379
		x"00",	--4380
		x"3c",	--4381
		x"40",	--4382
		x"00",	--4383
		x"5b",	--4384
		x"4a",	--4385
		x"00",	--4386
		x"48",	--4387
		x"53",	--4388
		x"41",	--4389
		x"00",	--4390
		x"49",	--4391
		x"44",	--4392
		x"47",	--4393
		x"12",	--4394
		x"e3",	--4395
		x"4e",	--4396
		x"4f",	--4397
		x"53",	--4398
		x"93",	--4399
		x"23",	--4400
		x"93",	--4401
		x"23",	--4402
		x"43",	--4403
		x"00",	--4404
		x"43",	--4405
		x"00",	--4406
		x"3c",	--4407
		x"41",	--4408
		x"00",	--4409
		x"41",	--4410
		x"50",	--4411
		x"00",	--4412
		x"41",	--4413
		x"00",	--4414
		x"47",	--4415
		x"12",	--4416
		x"e4",	--4417
		x"4f",	--4418
		x"90",	--4419
		x"00",	--4420
		x"34",	--4421
		x"50",	--4422
		x"00",	--4423
		x"4d",	--4424
		x"00",	--4425
		x"3c",	--4426
		x"4f",	--4427
		x"b3",	--4428
		x"00",	--4429
		x"24",	--4430
		x"40",	--4431
		x"00",	--4432
		x"3c",	--4433
		x"40",	--4434
		x"00",	--4435
		x"5d",	--4436
		x"4c",	--4437
		x"00",	--4438
		x"48",	--4439
		x"53",	--4440
		x"41",	--4441
		x"00",	--4442
		x"47",	--4443
		x"12",	--4444
		x"e4",	--4445
		x"4f",	--4446
		x"53",	--4447
		x"93",	--4448
		x"23",	--4449
		x"43",	--4450
		x"00",	--4451
		x"90",	--4452
		x"00",	--4453
		x"00",	--4454
		x"24",	--4455
		x"43",	--4456
		x"00",	--4457
		x"93",	--4458
		x"00",	--4459
		x"24",	--4460
		x"41",	--4461
		x"50",	--4462
		x"00",	--4463
		x"4f",	--4464
		x"00",	--4465
		x"41",	--4466
		x"00",	--4467
		x"10",	--4468
		x"11",	--4469
		x"10",	--4470
		x"11",	--4471
		x"4a",	--4472
		x"00",	--4473
		x"46",	--4474
		x"00",	--4475
		x"46",	--4476
		x"10",	--4477
		x"11",	--4478
		x"10",	--4479
		x"11",	--4480
		x"4a",	--4481
		x"00",	--4482
		x"41",	--4483
		x"00",	--4484
		x"41",	--4485
		x"00",	--4486
		x"81",	--4487
		x"00",	--4488
		x"71",	--4489
		x"00",	--4490
		x"83",	--4491
		x"91",	--4492
		x"00",	--4493
		x"2c",	--4494
		x"d3",	--4495
		x"00",	--4496
		x"41",	--4497
		x"00",	--4498
		x"8c",	--4499
		x"4e",	--4500
		x"00",	--4501
		x"3c",	--4502
		x"93",	--4503
		x"00",	--4504
		x"24",	--4505
		x"41",	--4506
		x"00",	--4507
		x"00",	--4508
		x"12",	--4509
		x"00",	--4510
		x"12",	--4511
		x"00",	--4512
		x"41",	--4513
		x"00",	--4514
		x"46",	--4515
		x"53",	--4516
		x"41",	--4517
		x"00",	--4518
		x"12",	--4519
		x"db",	--4520
		x"52",	--4521
		x"5f",	--4522
		x"00",	--4523
		x"3c",	--4524
		x"49",	--4525
		x"11",	--4526
		x"12",	--4527
		x"00",	--4528
		x"49",	--4529
		x"58",	--4530
		x"91",	--4531
		x"00",	--4532
		x"2b",	--4533
		x"49",	--4534
		x"00",	--4535
		x"4e",	--4536
		x"00",	--4537
		x"43",	--4538
		x"3c",	--4539
		x"41",	--4540
		x"00",	--4541
		x"00",	--4542
		x"43",	--4543
		x"00",	--4544
		x"43",	--4545
		x"00",	--4546
		x"3c",	--4547
		x"4e",	--4548
		x"43",	--4549
		x"00",	--4550
		x"43",	--4551
		x"00",	--4552
		x"43",	--4553
		x"41",	--4554
		x"00",	--4555
		x"46",	--4556
		x"93",	--4557
		x"24",	--4558
		x"40",	--4559
		x"dd",	--4560
		x"41",	--4561
		x"00",	--4562
		x"50",	--4563
		x"00",	--4564
		x"41",	--4565
		x"41",	--4566
		x"41",	--4567
		x"41",	--4568
		x"41",	--4569
		x"41",	--4570
		x"41",	--4571
		x"41",	--4572
		x"41",	--4573
		x"43",	--4574
		x"93",	--4575
		x"34",	--4576
		x"40",	--4577
		x"00",	--4578
		x"e3",	--4579
		x"53",	--4580
		x"93",	--4581
		x"34",	--4582
		x"e3",	--4583
		x"e3",	--4584
		x"53",	--4585
		x"12",	--4586
		x"12",	--4587
		x"e4",	--4588
		x"41",	--4589
		x"b3",	--4590
		x"24",	--4591
		x"e3",	--4592
		x"53",	--4593
		x"b3",	--4594
		x"24",	--4595
		x"e3",	--4596
		x"53",	--4597
		x"41",	--4598
		x"12",	--4599
		x"e3",	--4600
		x"4e",	--4601
		x"41",	--4602
		x"12",	--4603
		x"12",	--4604
		x"12",	--4605
		x"40",	--4606
		x"00",	--4607
		x"4c",	--4608
		x"4d",	--4609
		x"43",	--4610
		x"43",	--4611
		x"5e",	--4612
		x"6f",	--4613
		x"6c",	--4614
		x"6d",	--4615
		x"9b",	--4616
		x"28",	--4617
		x"20",	--4618
		x"9a",	--4619
		x"28",	--4620
		x"8a",	--4621
		x"7b",	--4622
		x"d3",	--4623
		x"83",	--4624
		x"23",	--4625
		x"41",	--4626
		x"41",	--4627
		x"41",	--4628
		x"41",	--4629
		x"12",	--4630
		x"e3",	--4631
		x"4c",	--4632
		x"4d",	--4633
		x"41",	--4634
		x"12",	--4635
		x"43",	--4636
		x"93",	--4637
		x"34",	--4638
		x"40",	--4639
		x"00",	--4640
		x"e3",	--4641
		x"e3",	--4642
		x"53",	--4643
		x"63",	--4644
		x"93",	--4645
		x"34",	--4646
		x"e3",	--4647
		x"e3",	--4648
		x"e3",	--4649
		x"53",	--4650
		x"63",	--4651
		x"12",	--4652
		x"e3",	--4653
		x"b3",	--4654
		x"24",	--4655
		x"e3",	--4656
		x"e3",	--4657
		x"53",	--4658
		x"63",	--4659
		x"b3",	--4660
		x"24",	--4661
		x"e3",	--4662
		x"e3",	--4663
		x"53",	--4664
		x"63",	--4665
		x"41",	--4666
		x"41",	--4667
		x"12",	--4668
		x"e4",	--4669
		x"4c",	--4670
		x"4d",	--4671
		x"41",	--4672
		x"40",	--4673
		x"00",	--4674
		x"4e",	--4675
		x"43",	--4676
		x"5f",	--4677
		x"6e",	--4678
		x"9d",	--4679
		x"28",	--4680
		x"8d",	--4681
		x"d3",	--4682
		x"83",	--4683
		x"23",	--4684
		x"41",	--4685
		x"12",	--4686
		x"e4",	--4687
		x"4e",	--4688
		x"41",	--4689
		x"12",	--4690
		x"12",	--4691
		x"12",	--4692
		x"12",	--4693
		x"12",	--4694
		x"00",	--4695
		x"48",	--4696
		x"49",	--4697
		x"4a",	--4698
		x"4b",	--4699
		x"43",	--4700
		x"43",	--4701
		x"43",	--4702
		x"43",	--4703
		x"5c",	--4704
		x"6d",	--4705
		x"6e",	--4706
		x"6f",	--4707
		x"68",	--4708
		x"69",	--4709
		x"6a",	--4710
		x"6b",	--4711
		x"97",	--4712
		x"28",	--4713
		x"20",	--4714
		x"96",	--4715
		x"28",	--4716
		x"20",	--4717
		x"95",	--4718
		x"28",	--4719
		x"20",	--4720
		x"94",	--4721
		x"28",	--4722
		x"84",	--4723
		x"75",	--4724
		x"76",	--4725
		x"77",	--4726
		x"d3",	--4727
		x"83",	--4728
		x"00",	--4729
		x"23",	--4730
		x"53",	--4731
		x"41",	--4732
		x"41",	--4733
		x"41",	--4734
		x"41",	--4735
		x"41",	--4736
		x"12",	--4737
		x"12",	--4738
		x"12",	--4739
		x"12",	--4740
		x"41",	--4741
		x"00",	--4742
		x"41",	--4743
		x"00",	--4744
		x"41",	--4745
		x"00",	--4746
		x"41",	--4747
		x"00",	--4748
		x"12",	--4749
		x"e4",	--4750
		x"41",	--4751
		x"41",	--4752
		x"41",	--4753
		x"41",	--4754
		x"41",	--4755
		x"12",	--4756
		x"12",	--4757
		x"12",	--4758
		x"12",	--4759
		x"41",	--4760
		x"00",	--4761
		x"41",	--4762
		x"00",	--4763
		x"41",	--4764
		x"00",	--4765
		x"41",	--4766
		x"00",	--4767
		x"12",	--4768
		x"e4",	--4769
		x"48",	--4770
		x"49",	--4771
		x"4a",	--4772
		x"4b",	--4773
		x"41",	--4774
		x"41",	--4775
		x"41",	--4776
		x"41",	--4777
		x"41",	--4778
		x"12",	--4779
		x"12",	--4780
		x"12",	--4781
		x"12",	--4782
		x"12",	--4783
		x"41",	--4784
		x"00",	--4785
		x"41",	--4786
		x"00",	--4787
		x"41",	--4788
		x"00",	--4789
		x"41",	--4790
		x"00",	--4791
		x"12",	--4792
		x"e4",	--4793
		x"41",	--4794
		x"00",	--4795
		x"48",	--4796
		x"00",	--4797
		x"49",	--4798
		x"00",	--4799
		x"4a",	--4800
		x"00",	--4801
		x"4b",	--4802
		x"00",	--4803
		x"41",	--4804
		x"41",	--4805
		x"41",	--4806
		x"41",	--4807
		x"41",	--4808
		x"41",	--4809
		x"13",	--4810
		x"d0",	--4811
		x"00",	--4812
		x"3f",	--4813
		x"61",	--4814
		x"74",	--4815
		x"6e",	--4816
		x"20",	--4817
		x"6f",	--4818
		x"20",	--4819
		x"20",	--4820
		x"65",	--4821
		x"20",	--4822
		x"62",	--4823
		x"6e",	--4824
		x"66",	--4825
		x"6c",	--4826
		x"0d",	--4827
		x"00",	--4828
		x"65",	--4829
		x"73",	--4830
		x"6f",	--4831
		x"6c",	--4832
		x"20",	--4833
		x"6f",	--4834
		x"20",	--4835
		x"65",	--4836
		x"20",	--4837
		x"68",	--4838
		x"74",	--4839
		x"0a",	--4840
		x"53",	--4841
		x"6f",	--4842
		x"0d",	--4843
		x"00",	--4844
		x"72",	--4845
		x"6f",	--4846
		x"3a",	--4847
		x"6d",	--4848
		x"73",	--4849
		x"69",	--4850
		x"67",	--4851
		x"61",	--4852
		x"67",	--4853
		x"6d",	--4854
		x"6e",	--4855
		x"0d",	--4856
		x"00",	--4857
		x"6f",	--4858
		x"72",	--4859
		x"63",	--4860
		x"20",	--4861
		x"73",	--4862
		x"67",	--4863
		x"3a",	--4864
		x"0a",	--4865
		x"09",	--4866
		x"73",	--4867
		x"4c",	--4868
		x"46",	--4869
		x"20",	--4870
		x"49",	--4871
		x"48",	--4872
		x"20",	--4873
		x"54",	--4874
		x"4d",	--4875
		x"4f",	--4876
		x"54",	--4877
		x"0d",	--4878
		x"00",	--4879
		x"64",	--4880
		x"25",	--4881
		x"0d",	--4882
		x"00",	--4883
		x"6c",	--4884
		x"20",	--4885
		x"6c",	--4886
		x"00",	--4887
		x"73",	--4888
		x"0a",	--4889
		x"00",	--4890
		x"c5",	--4891
		x"c5",	--4892
		x"c5",	--4893
		x"c5",	--4894
		x"c5",	--4895
		x"c5",	--4896
		x"c5",	--4897
		x"c5",	--4898
		x"0a",	--4899
		x"3d",	--4900
		x"3d",	--4901
		x"3d",	--4902
		x"4d",	--4903
		x"72",	--4904
		x"65",	--4905
		x"20",	--4906
		x"43",	--4907
		x"20",	--4908
		x"3d",	--4909
		x"3d",	--4910
		x"3d",	--4911
		x"0a",	--4912
		x"69",	--4913
		x"74",	--4914
		x"72",	--4915
		x"63",	--4916
		x"69",	--4917
		x"65",	--4918
		x"6d",	--4919
		x"64",	--4920
		x"00",	--4921
		x"72",	--4922
		x"74",	--4923
		x"00",	--4924
		x"65",	--4925
		x"64",	--4926
		x"70",	--4927
		x"6d",	--4928
		x"65",	--4929
		x"63",	--4930
		x"64",	--4931
		x"72",	--4932
		x"73",	--4933
		x"65",	--4934
		x"64",	--4935
		x"63",	--4936
		x"6e",	--4937
		x"72",	--4938
		x"6c",	--4939
		x"65",	--4940
		x"00",	--4941
		x"70",	--4942
		x"65",	--4943
		x"20",	--4944
		x"6f",	--4945
		x"66",	--4946
		x"67",	--4947
		x"72",	--4948
		x"74",	--4949
		x"6f",	--4950
		x"00",	--4951
		x"6f",	--4952
		x"74",	--4953
		x"6f",	--4954
		x"64",	--4955
		x"72",	--4956
		x"0d",	--4957
		x"00",	--4958
		x"20",	--4959
		x"00",	--4960
		x"63",	--4961
		x"00",	--4962
		x"72",	--4963
		x"74",	--4964
		x"0a",	--4965
		x"00",	--4966
		x"72",	--4967
		x"6f",	--4968
		x"3a",	--4969
		x"6d",	--4970
		x"73",	--4971
		x"69",	--4972
		x"67",	--4973
		x"61",	--4974
		x"67",	--4975
		x"6d",	--4976
		x"6e",	--4977
		x"0d",	--4978
		x"00",	--4979
		x"6f",	--4980
		x"72",	--4981
		x"63",	--4982
		x"20",	--4983
		x"73",	--4984
		x"67",	--4985
		x"3a",	--4986
		x"0a",	--4987
		x"09",	--4988
		x"73",	--4989
		x"52",	--4990
		x"47",	--4991
		x"53",	--4992
		x"45",	--4993
		x"20",	--4994
		x"41",	--4995
		x"55",	--4996
		x"0d",	--4997
		x"00",	--4998
		x"3d",	--4999
		x"64",	--5000
		x"76",	--5001
		x"25",	--5002
		x"0d",	--5003
		x"00",	--5004
		x"25",	--5005
		x"20",	--5006
		x"45",	--5007
		x"49",	--5008
		x"54",	--5009
		x"52",	--5010
		x"0a",	--5011
		x"72",	--5012
		x"61",	--5013
		x"0a",	--5014
		x"00",	--5015
		x"63",	--5016
		x"69",	--5017
		x"20",	--5018
		x"6f",	--5019
		x"20",	--5020
		x"20",	--5021
		x"75",	--5022
		x"62",	--5023
		x"72",	--5024
		x"0a",	--5025
		x"25",	--5026
		x"20",	--5027
		x"73",	--5028
		x"0a",	--5029
		x"25",	--5030
		x"3a",	--5031
		x"6e",	--5032
		x"20",	--5033
		x"75",	--5034
		x"68",	--5035
		x"63",	--5036
		x"6d",	--5037
		x"61",	--5038
		x"64",	--5039
		x"0a",	--5040
		x"00",	--5041
		x"cd",	--5042
		x"cc",	--5043
		x"cc",	--5044
		x"cc",	--5045
		x"cc",	--5046
		x"cc",	--5047
		x"cc",	--5048
		x"cc",	--5049
		x"cc",	--5050
		x"cc",	--5051
		x"cc",	--5052
		x"cc",	--5053
		x"cc",	--5054
		x"cc",	--5055
		x"cc",	--5056
		x"cc",	--5057
		x"cc",	--5058
		x"cc",	--5059
		x"cc",	--5060
		x"cc",	--5061
		x"cc",	--5062
		x"cc",	--5063
		x"cc",	--5064
		x"cc",	--5065
		x"cc",	--5066
		x"cc",	--5067
		x"cc",	--5068
		x"cc",	--5069
		x"cc",	--5070
		x"cd",	--5071
		x"cc",	--5072
		x"cc",	--5073
		x"cc",	--5074
		x"cc",	--5075
		x"cc",	--5076
		x"cc",	--5077
		x"cc",	--5078
		x"cc",	--5079
		x"cc",	--5080
		x"cc",	--5081
		x"cc",	--5082
		x"cc",	--5083
		x"cc",	--5084
		x"cc",	--5085
		x"cc",	--5086
		x"cc",	--5087
		x"cc",	--5088
		x"cc",	--5089
		x"cc",	--5090
		x"cc",	--5091
		x"cc",	--5092
		x"cc",	--5093
		x"cc",	--5094
		x"cc",	--5095
		x"cc",	--5096
		x"cc",	--5097
		x"cc",	--5098
		x"cc",	--5099
		x"cc",	--5100
		x"cc",	--5101
		x"cc",	--5102
		x"cd",	--5103
		x"cd",	--5104
		x"cd",	--5105
		x"cc",	--5106
		x"cc",	--5107
		x"cc",	--5108
		x"cc",	--5109
		x"cc",	--5110
		x"cc",	--5111
		x"cc",	--5112
		x"cc",	--5113
		x"cc",	--5114
		x"cc",	--5115
		x"cc",	--5116
		x"cc",	--5117
		x"cc",	--5118
		x"cc",	--5119
		x"cc",	--5120
		x"cc",	--5121
		x"cc",	--5122
		x"cc",	--5123
		x"cc",	--5124
		x"cc",	--5125
		x"31",	--5126
		x"33",	--5127
		x"35",	--5128
		x"37",	--5129
		x"39",	--5130
		x"62",	--5131
		x"64",	--5132
		x"66",	--5133
		x"00",	--5134
		x"00",	--5135
		x"00",	--5136
		x"00",	--5137
		x"00",	--5138
		x"01",	--5139
		x"02",	--5140
		x"03",	--5141
		x"03",	--5142
		x"04",	--5143
		x"04",	--5144
		x"04",	--5145
		x"04",	--5146
		x"05",	--5147
		x"05",	--5148
		x"05",	--5149
		x"05",	--5150
		x"05",	--5151
		x"05",	--5152
		x"05",	--5153
		x"05",	--5154
		x"06",	--5155
		x"06",	--5156
		x"06",	--5157
		x"06",	--5158
		x"06",	--5159
		x"06",	--5160
		x"06",	--5161
		x"06",	--5162
		x"06",	--5163
		x"06",	--5164
		x"06",	--5165
		x"06",	--5166
		x"06",	--5167
		x"06",	--5168
		x"06",	--5169
		x"06",	--5170
		x"07",	--5171
		x"07",	--5172
		x"07",	--5173
		x"07",	--5174
		x"07",	--5175
		x"07",	--5176
		x"07",	--5177
		x"07",	--5178
		x"07",	--5179
		x"07",	--5180
		x"07",	--5181
		x"07",	--5182
		x"07",	--5183
		x"07",	--5184
		x"07",	--5185
		x"07",	--5186
		x"07",	--5187
		x"07",	--5188
		x"07",	--5189
		x"07",	--5190
		x"07",	--5191
		x"07",	--5192
		x"07",	--5193
		x"07",	--5194
		x"07",	--5195
		x"07",	--5196
		x"07",	--5197
		x"07",	--5198
		x"07",	--5199
		x"07",	--5200
		x"07",	--5201
		x"07",	--5202
		x"08",	--5203
		x"08",	--5204
		x"08",	--5205
		x"08",	--5206
		x"08",	--5207
		x"08",	--5208
		x"08",	--5209
		x"08",	--5210
		x"08",	--5211
		x"08",	--5212
		x"08",	--5213
		x"08",	--5214
		x"08",	--5215
		x"08",	--5216
		x"08",	--5217
		x"08",	--5218
		x"08",	--5219
		x"08",	--5220
		x"08",	--5221
		x"08",	--5222
		x"08",	--5223
		x"08",	--5224
		x"08",	--5225
		x"08",	--5226
		x"08",	--5227
		x"08",	--5228
		x"08",	--5229
		x"08",	--5230
		x"08",	--5231
		x"08",	--5232
		x"08",	--5233
		x"08",	--5234
		x"08",	--5235
		x"08",	--5236
		x"08",	--5237
		x"08",	--5238
		x"08",	--5239
		x"08",	--5240
		x"08",	--5241
		x"08",	--5242
		x"08",	--5243
		x"08",	--5244
		x"08",	--5245
		x"08",	--5246
		x"08",	--5247
		x"08",	--5248
		x"08",	--5249
		x"08",	--5250
		x"08",	--5251
		x"08",	--5252
		x"08",	--5253
		x"08",	--5254
		x"08",	--5255
		x"08",	--5256
		x"08",	--5257
		x"08",	--5258
		x"08",	--5259
		x"08",	--5260
		x"08",	--5261
		x"08",	--5262
		x"08",	--5263
		x"08",	--5264
		x"08",	--5265
		x"08",	--5266
		x"6e",	--5267
		x"6c",	--5268
		x"29",	--5269
		x"00",	--5270
		x"ff",	--5271
		x"ff",	--5272
		x"65",	--5273
		x"70",	--5274
		x"00",	--5275
		x"ff",	--5276
		x"ff",	--5277
		x"ff",	--5278
		x"ff",	--5279
		x"ff",	--5280
		x"ff",	--5281
		x"ff",	--5282
		x"ff",	--5283
		x"ff",	--5284
		x"ff",	--5285
		x"ff",	--5286
		x"ff",	--5287
		x"ff",	--5288
		x"ff",	--5289
		x"ff",	--5290
		x"ff",	--5291
		x"ff",	--5292
		x"ff",	--5293
		x"ff",	--5294
		x"ff",	--5295
		x"ff",	--5296
		x"ff",	--5297
		x"ff",	--5298
		x"ff",	--5299
		x"ff",	--5300
		x"ff",	--5301
		x"ff",	--5302
		x"ff",	--5303
		x"ff",	--5304
		x"ff",	--5305
		x"ff",	--5306
		x"ff",	--5307
		x"ff",	--5308
		x"ff",	--5309
		x"ff",	--5310
		x"ff",	--5311
		x"ff",	--5312
		x"ff",	--5313
		x"ff",	--5314
		x"ff",	--5315
		x"ff",	--5316
		x"ff",	--5317
		x"ff",	--5318
		x"ff",	--5319
		x"ff",	--5320
		x"ff",	--5321
		x"ff",	--5322
		x"ff",	--5323
		x"ff",	--5324
		x"ff",	--5325
		x"ff",	--5326
		x"ff",	--5327
		x"ff",	--5328
		x"ff",	--5329
		x"ff",	--5330
		x"ff",	--5331
		x"ff",	--5332
		x"ff",	--5333
		x"ff",	--5334
		x"ff",	--5335
		x"ff",	--5336
		x"ff",	--5337
		x"ff",	--5338
		x"ff",	--5339
		x"ff",	--5340
		x"ff",	--5341
		x"ff",	--5342
		x"ff",	--5343
		x"ff",	--5344
		x"ff",	--5345
		x"ff",	--5346
		x"ff",	--5347
		x"ff",	--5348
		x"ff",	--5349
		x"ff",	--5350
		x"ff",	--5351
		x"ff",	--5352
		x"ff",	--5353
		x"ff",	--5354
		x"ff",	--5355
		x"ff",	--5356
		x"ff",	--5357
		x"ff",	--5358
		x"ff",	--5359
		x"ff",	--5360
		x"ff",	--5361
		x"ff",	--5362
		x"ff",	--5363
		x"ff",	--5364
		x"ff",	--5365
		x"ff",	--5366
		x"ff",	--5367
		x"ff",	--5368
		x"ff",	--5369
		x"ff",	--5370
		x"ff",	--5371
		x"ff",	--5372
		x"ff",	--5373
		x"ff",	--5374
		x"ff",	--5375
		x"ff",	--5376
		x"ff",	--5377
		x"ff",	--5378
		x"ff",	--5379
		x"ff",	--5380
		x"ff",	--5381
		x"ff",	--5382
		x"ff",	--5383
		x"ff",	--5384
		x"ff",	--5385
		x"ff",	--5386
		x"ff",	--5387
		x"ff",	--5388
		x"ff",	--5389
		x"ff",	--5390
		x"ff",	--5391
		x"ff",	--5392
		x"ff",	--5393
		x"ff",	--5394
		x"ff",	--5395
		x"ff",	--5396
		x"ff",	--5397
		x"ff",	--5398
		x"ff",	--5399
		x"ff",	--5400
		x"ff",	--5401
		x"ff",	--5402
		x"ff",	--5403
		x"ff",	--5404
		x"ff",	--5405
		x"ff",	--5406
		x"ff",	--5407
		x"ff",	--5408
		x"ff",	--5409
		x"ff",	--5410
		x"ff",	--5411
		x"ff",	--5412
		x"ff",	--5413
		x"ff",	--5414
		x"ff",	--5415
		x"ff",	--5416
		x"ff",	--5417
		x"ff",	--5418
		x"ff",	--5419
		x"ff",	--5420
		x"ff",	--5421
		x"ff",	--5422
		x"ff",	--5423
		x"ff",	--5424
		x"ff",	--5425
		x"ff",	--5426
		x"ff",	--5427
		x"ff",	--5428
		x"ff",	--5429
		x"ff",	--5430
		x"ff",	--5431
		x"ff",	--5432
		x"ff",	--5433
		x"ff",	--5434
		x"ff",	--5435
		x"ff",	--5436
		x"ff",	--5437
		x"ff",	--5438
		x"ff",	--5439
		x"ff",	--5440
		x"ff",	--5441
		x"ff",	--5442
		x"ff",	--5443
		x"ff",	--5444
		x"ff",	--5445
		x"ff",	--5446
		x"ff",	--5447
		x"ff",	--5448
		x"ff",	--5449
		x"ff",	--5450
		x"ff",	--5451
		x"ff",	--5452
		x"ff",	--5453
		x"ff",	--5454
		x"ff",	--5455
		x"ff",	--5456
		x"ff",	--5457
		x"ff",	--5458
		x"ff",	--5459
		x"ff",	--5460
		x"ff",	--5461
		x"ff",	--5462
		x"ff",	--5463
		x"ff",	--5464
		x"ff",	--5465
		x"ff",	--5466
		x"ff",	--5467
		x"ff",	--5468
		x"ff",	--5469
		x"ff",	--5470
		x"ff",	--5471
		x"ff",	--5472
		x"ff",	--5473
		x"ff",	--5474
		x"ff",	--5475
		x"ff",	--5476
		x"ff",	--5477
		x"ff",	--5478
		x"ff",	--5479
		x"ff",	--5480
		x"ff",	--5481
		x"ff",	--5482
		x"ff",	--5483
		x"ff",	--5484
		x"ff",	--5485
		x"ff",	--5486
		x"ff",	--5487
		x"ff",	--5488
		x"ff",	--5489
		x"ff",	--5490
		x"ff",	--5491
		x"ff",	--5492
		x"ff",	--5493
		x"ff",	--5494
		x"ff",	--5495
		x"ff",	--5496
		x"ff",	--5497
		x"ff",	--5498
		x"ff",	--5499
		x"ff",	--5500
		x"ff",	--5501
		x"ff",	--5502
		x"ff",	--5503
		x"ff",	--5504
		x"ff",	--5505
		x"ff",	--5506
		x"ff",	--5507
		x"ff",	--5508
		x"ff",	--5509
		x"ff",	--5510
		x"ff",	--5511
		x"ff",	--5512
		x"ff",	--5513
		x"ff",	--5514
		x"ff",	--5515
		x"ff",	--5516
		x"ff",	--5517
		x"ff",	--5518
		x"ff",	--5519
		x"ff",	--5520
		x"ff",	--5521
		x"ff",	--5522
		x"ff",	--5523
		x"ff",	--5524
		x"ff",	--5525
		x"ff",	--5526
		x"ff",	--5527
		x"ff",	--5528
		x"ff",	--5529
		x"ff",	--5530
		x"ff",	--5531
		x"ff",	--5532
		x"ff",	--5533
		x"ff",	--5534
		x"ff",	--5535
		x"ff",	--5536
		x"ff",	--5537
		x"ff",	--5538
		x"ff",	--5539
		x"ff",	--5540
		x"ff",	--5541
		x"ff",	--5542
		x"ff",	--5543
		x"ff",	--5544
		x"ff",	--5545
		x"ff",	--5546
		x"ff",	--5547
		x"ff",	--5548
		x"ff",	--5549
		x"ff",	--5550
		x"ff",	--5551
		x"ff",	--5552
		x"ff",	--5553
		x"ff",	--5554
		x"ff",	--5555
		x"ff",	--5556
		x"ff",	--5557
		x"ff",	--5558
		x"ff",	--5559
		x"ff",	--5560
		x"ff",	--5561
		x"ff",	--5562
		x"ff",	--5563
		x"ff",	--5564
		x"ff",	--5565
		x"ff",	--5566
		x"ff",	--5567
		x"ff",	--5568
		x"ff",	--5569
		x"ff",	--5570
		x"ff",	--5571
		x"ff",	--5572
		x"ff",	--5573
		x"ff",	--5574
		x"ff",	--5575
		x"ff",	--5576
		x"ff",	--5577
		x"ff",	--5578
		x"ff",	--5579
		x"ff",	--5580
		x"ff",	--5581
		x"ff",	--5582
		x"ff",	--5583
		x"ff",	--5584
		x"ff",	--5585
		x"ff",	--5586
		x"ff",	--5587
		x"ff",	--5588
		x"ff",	--5589
		x"ff",	--5590
		x"ff",	--5591
		x"ff",	--5592
		x"ff",	--5593
		x"ff",	--5594
		x"ff",	--5595
		x"ff",	--5596
		x"ff",	--5597
		x"ff",	--5598
		x"ff",	--5599
		x"ff",	--5600
		x"ff",	--5601
		x"ff",	--5602
		x"ff",	--5603
		x"ff",	--5604
		x"ff",	--5605
		x"ff",	--5606
		x"ff",	--5607
		x"ff",	--5608
		x"ff",	--5609
		x"ff",	--5610
		x"ff",	--5611
		x"ff",	--5612
		x"ff",	--5613
		x"ff",	--5614
		x"ff",	--5615
		x"ff",	--5616
		x"ff",	--5617
		x"ff",	--5618
		x"ff",	--5619
		x"ff",	--5620
		x"ff",	--5621
		x"ff",	--5622
		x"ff",	--5623
		x"ff",	--5624
		x"ff",	--5625
		x"ff",	--5626
		x"ff",	--5627
		x"ff",	--5628
		x"ff",	--5629
		x"ff",	--5630
		x"ff",	--5631
		x"ff",	--5632
		x"ff",	--5633
		x"ff",	--5634
		x"ff",	--5635
		x"ff",	--5636
		x"ff",	--5637
		x"ff",	--5638
		x"ff",	--5639
		x"ff",	--5640
		x"ff",	--5641
		x"ff",	--5642
		x"ff",	--5643
		x"ff",	--5644
		x"ff",	--5645
		x"ff",	--5646
		x"ff",	--5647
		x"ff",	--5648
		x"ff",	--5649
		x"ff",	--5650
		x"ff",	--5651
		x"ff",	--5652
		x"ff",	--5653
		x"ff",	--5654
		x"ff",	--5655
		x"ff",	--5656
		x"ff",	--5657
		x"ff",	--5658
		x"ff",	--5659
		x"ff",	--5660
		x"ff",	--5661
		x"ff",	--5662
		x"ff",	--5663
		x"ff",	--5664
		x"ff",	--5665
		x"ff",	--5666
		x"ff",	--5667
		x"ff",	--5668
		x"ff",	--5669
		x"ff",	--5670
		x"ff",	--5671
		x"ff",	--5672
		x"ff",	--5673
		x"ff",	--5674
		x"ff",	--5675
		x"ff",	--5676
		x"ff",	--5677
		x"ff",	--5678
		x"ff",	--5679
		x"ff",	--5680
		x"ff",	--5681
		x"ff",	--5682
		x"ff",	--5683
		x"ff",	--5684
		x"ff",	--5685
		x"ff",	--5686
		x"ff",	--5687
		x"ff",	--5688
		x"ff",	--5689
		x"ff",	--5690
		x"ff",	--5691
		x"ff",	--5692
		x"ff",	--5693
		x"ff",	--5694
		x"ff",	--5695
		x"ff",	--5696
		x"ff",	--5697
		x"ff",	--5698
		x"ff",	--5699
		x"ff",	--5700
		x"ff",	--5701
		x"ff",	--5702
		x"ff",	--5703
		x"ff",	--5704
		x"ff",	--5705
		x"ff",	--5706
		x"ff",	--5707
		x"ff",	--5708
		x"ff",	--5709
		x"ff",	--5710
		x"ff",	--5711
		x"ff",	--5712
		x"ff",	--5713
		x"ff",	--5714
		x"ff",	--5715
		x"ff",	--5716
		x"ff",	--5717
		x"ff",	--5718
		x"ff",	--5719
		x"ff",	--5720
		x"ff",	--5721
		x"ff",	--5722
		x"ff",	--5723
		x"ff",	--5724
		x"ff",	--5725
		x"ff",	--5726
		x"ff",	--5727
		x"ff",	--5728
		x"ff",	--5729
		x"ff",	--5730
		x"ff",	--5731
		x"ff",	--5732
		x"ff",	--5733
		x"ff",	--5734
		x"ff",	--5735
		x"ff",	--5736
		x"ff",	--5737
		x"ff",	--5738
		x"ff",	--5739
		x"ff",	--5740
		x"ff",	--5741
		x"ff",	--5742
		x"ff",	--5743
		x"ff",	--5744
		x"ff",	--5745
		x"ff",	--5746
		x"ff",	--5747
		x"ff",	--5748
		x"ff",	--5749
		x"ff",	--5750
		x"ff",	--5751
		x"ff",	--5752
		x"ff",	--5753
		x"ff",	--5754
		x"ff",	--5755
		x"ff",	--5756
		x"ff",	--5757
		x"ff",	--5758
		x"ff",	--5759
		x"ff",	--5760
		x"ff",	--5761
		x"ff",	--5762
		x"ff",	--5763
		x"ff",	--5764
		x"ff",	--5765
		x"ff",	--5766
		x"ff",	--5767
		x"ff",	--5768
		x"ff",	--5769
		x"ff",	--5770
		x"ff",	--5771
		x"ff",	--5772
		x"ff",	--5773
		x"ff",	--5774
		x"ff",	--5775
		x"ff",	--5776
		x"ff",	--5777
		x"ff",	--5778
		x"ff",	--5779
		x"ff",	--5780
		x"ff",	--5781
		x"ff",	--5782
		x"ff",	--5783
		x"ff",	--5784
		x"ff",	--5785
		x"ff",	--5786
		x"ff",	--5787
		x"ff",	--5788
		x"ff",	--5789
		x"ff",	--5790
		x"ff",	--5791
		x"ff",	--5792
		x"ff",	--5793
		x"ff",	--5794
		x"ff",	--5795
		x"ff",	--5796
		x"ff",	--5797
		x"ff",	--5798
		x"ff",	--5799
		x"ff",	--5800
		x"ff",	--5801
		x"ff",	--5802
		x"ff",	--5803
		x"ff",	--5804
		x"ff",	--5805
		x"ff",	--5806
		x"ff",	--5807
		x"ff",	--5808
		x"ff",	--5809
		x"ff",	--5810
		x"ff",	--5811
		x"ff",	--5812
		x"ff",	--5813
		x"ff",	--5814
		x"ff",	--5815
		x"ff",	--5816
		x"ff",	--5817
		x"ff",	--5818
		x"ff",	--5819
		x"ff",	--5820
		x"ff",	--5821
		x"ff",	--5822
		x"ff",	--5823
		x"ff",	--5824
		x"ff",	--5825
		x"ff",	--5826
		x"ff",	--5827
		x"ff",	--5828
		x"ff",	--5829
		x"ff",	--5830
		x"ff",	--5831
		x"ff",	--5832
		x"ff",	--5833
		x"ff",	--5834
		x"ff",	--5835
		x"ff",	--5836
		x"ff",	--5837
		x"ff",	--5838
		x"ff",	--5839
		x"ff",	--5840
		x"ff",	--5841
		x"ff",	--5842
		x"ff",	--5843
		x"ff",	--5844
		x"ff",	--5845
		x"ff",	--5846
		x"ff",	--5847
		x"ff",	--5848
		x"ff",	--5849
		x"ff",	--5850
		x"ff",	--5851
		x"ff",	--5852
		x"ff",	--5853
		x"ff",	--5854
		x"ff",	--5855
		x"ff",	--5856
		x"ff",	--5857
		x"ff",	--5858
		x"ff",	--5859
		x"ff",	--5860
		x"ff",	--5861
		x"ff",	--5862
		x"ff",	--5863
		x"ff",	--5864
		x"ff",	--5865
		x"ff",	--5866
		x"ff",	--5867
		x"ff",	--5868
		x"ff",	--5869
		x"ff",	--5870
		x"ff",	--5871
		x"ff",	--5872
		x"ff",	--5873
		x"ff",	--5874
		x"ff",	--5875
		x"ff",	--5876
		x"ff",	--5877
		x"ff",	--5878
		x"ff",	--5879
		x"ff",	--5880
		x"ff",	--5881
		x"ff",	--5882
		x"ff",	--5883
		x"ff",	--5884
		x"ff",	--5885
		x"ff",	--5886
		x"ff",	--5887
		x"ff",	--5888
		x"ff",	--5889
		x"ff",	--5890
		x"ff",	--5891
		x"ff",	--5892
		x"ff",	--5893
		x"ff",	--5894
		x"ff",	--5895
		x"ff",	--5896
		x"ff",	--5897
		x"ff",	--5898
		x"ff",	--5899
		x"ff",	--5900
		x"ff",	--5901
		x"ff",	--5902
		x"ff",	--5903
		x"ff",	--5904
		x"ff",	--5905
		x"ff",	--5906
		x"ff",	--5907
		x"ff",	--5908
		x"ff",	--5909
		x"ff",	--5910
		x"ff",	--5911
		x"ff",	--5912
		x"ff",	--5913
		x"ff",	--5914
		x"ff",	--5915
		x"ff",	--5916
		x"ff",	--5917
		x"ff",	--5918
		x"ff",	--5919
		x"ff",	--5920
		x"ff",	--5921
		x"ff",	--5922
		x"ff",	--5923
		x"ff",	--5924
		x"ff",	--5925
		x"ff",	--5926
		x"ff",	--5927
		x"ff",	--5928
		x"ff",	--5929
		x"ff",	--5930
		x"ff",	--5931
		x"ff",	--5932
		x"ff",	--5933
		x"ff",	--5934
		x"ff",	--5935
		x"ff",	--5936
		x"ff",	--5937
		x"ff",	--5938
		x"ff",	--5939
		x"ff",	--5940
		x"ff",	--5941
		x"ff",	--5942
		x"ff",	--5943
		x"ff",	--5944
		x"ff",	--5945
		x"ff",	--5946
		x"ff",	--5947
		x"ff",	--5948
		x"ff",	--5949
		x"ff",	--5950
		x"ff",	--5951
		x"ff",	--5952
		x"ff",	--5953
		x"ff",	--5954
		x"ff",	--5955
		x"ff",	--5956
		x"ff",	--5957
		x"ff",	--5958
		x"ff",	--5959
		x"ff",	--5960
		x"ff",	--5961
		x"ff",	--5962
		x"ff",	--5963
		x"ff",	--5964
		x"ff",	--5965
		x"ff",	--5966
		x"ff",	--5967
		x"ff",	--5968
		x"ff",	--5969
		x"ff",	--5970
		x"ff",	--5971
		x"ff",	--5972
		x"ff",	--5973
		x"ff",	--5974
		x"ff",	--5975
		x"ff",	--5976
		x"ff",	--5977
		x"ff",	--5978
		x"ff",	--5979
		x"ff",	--5980
		x"ff",	--5981
		x"ff",	--5982
		x"ff",	--5983
		x"ff",	--5984
		x"ff",	--5985
		x"ff",	--5986
		x"ff",	--5987
		x"ff",	--5988
		x"ff",	--5989
		x"ff",	--5990
		x"ff",	--5991
		x"ff",	--5992
		x"ff",	--5993
		x"ff",	--5994
		x"ff",	--5995
		x"ff",	--5996
		x"ff",	--5997
		x"ff",	--5998
		x"ff",	--5999
		x"ff",	--6000
		x"ff",	--6001
		x"ff",	--6002
		x"ff",	--6003
		x"ff",	--6004
		x"ff",	--6005
		x"ff",	--6006
		x"ff",	--6007
		x"ff",	--6008
		x"ff",	--6009
		x"ff",	--6010
		x"ff",	--6011
		x"ff",	--6012
		x"ff",	--6013
		x"ff",	--6014
		x"ff",	--6015
		x"ff",	--6016
		x"ff",	--6017
		x"ff",	--6018
		x"ff",	--6019
		x"ff",	--6020
		x"ff",	--6021
		x"ff",	--6022
		x"ff",	--6023
		x"ff",	--6024
		x"ff",	--6025
		x"ff",	--6026
		x"ff",	--6027
		x"ff",	--6028
		x"ff",	--6029
		x"ff",	--6030
		x"ff",	--6031
		x"ff",	--6032
		x"ff",	--6033
		x"ff",	--6034
		x"ff",	--6035
		x"ff",	--6036
		x"ff",	--6037
		x"ff",	--6038
		x"ff",	--6039
		x"ff",	--6040
		x"ff",	--6041
		x"ff",	--6042
		x"ff",	--6043
		x"ff",	--6044
		x"ff",	--6045
		x"ff",	--6046
		x"ff",	--6047
		x"ff",	--6048
		x"ff",	--6049
		x"ff",	--6050
		x"ff",	--6051
		x"ff",	--6052
		x"ff",	--6053
		x"ff",	--6054
		x"ff",	--6055
		x"ff",	--6056
		x"ff",	--6057
		x"ff",	--6058
		x"ff",	--6059
		x"ff",	--6060
		x"ff",	--6061
		x"ff",	--6062
		x"ff",	--6063
		x"ff",	--6064
		x"ff",	--6065
		x"ff",	--6066
		x"ff",	--6067
		x"ff",	--6068
		x"ff",	--6069
		x"ff",	--6070
		x"ff",	--6071
		x"ff",	--6072
		x"ff",	--6073
		x"ff",	--6074
		x"ff",	--6075
		x"ff",	--6076
		x"ff",	--6077
		x"ff",	--6078
		x"ff",	--6079
		x"ff",	--6080
		x"ff",	--6081
		x"ff",	--6082
		x"ff",	--6083
		x"ff",	--6084
		x"ff",	--6085
		x"ff",	--6086
		x"ff",	--6087
		x"ff",	--6088
		x"ff",	--6089
		x"ff",	--6090
		x"ff",	--6091
		x"ff",	--6092
		x"ff",	--6093
		x"ff",	--6094
		x"ff",	--6095
		x"ff",	--6096
		x"ff",	--6097
		x"ff",	--6098
		x"ff",	--6099
		x"ff",	--6100
		x"ff",	--6101
		x"ff",	--6102
		x"ff",	--6103
		x"ff",	--6104
		x"ff",	--6105
		x"ff",	--6106
		x"ff",	--6107
		x"ff",	--6108
		x"ff",	--6109
		x"ff",	--6110
		x"ff",	--6111
		x"ff",	--6112
		x"ff",	--6113
		x"ff",	--6114
		x"ff",	--6115
		x"ff",	--6116
		x"ff",	--6117
		x"ff",	--6118
		x"ff",	--6119
		x"ff",	--6120
		x"ff",	--6121
		x"ff",	--6122
		x"ff",	--6123
		x"ff",	--6124
		x"ff",	--6125
		x"ff",	--6126
		x"ff",	--6127
		x"ff",	--6128
		x"ff",	--6129
		x"ff",	--6130
		x"ff",	--6131
		x"ff",	--6132
		x"ff",	--6133
		x"ff",	--6134
		x"ff",	--6135
		x"ff",	--6136
		x"ff",	--6137
		x"ff",	--6138
		x"ff",	--6139
		x"ff",	--6140
		x"ff",	--6141
		x"ff",	--6142
		x"ff",	--6143
		x"ff",	--6144
		x"ff",	--6145
		x"ff",	--6146
		x"ff",	--6147
		x"ff",	--6148
		x"ff",	--6149
		x"ff",	--6150
		x"ff",	--6151
		x"ff",	--6152
		x"ff",	--6153
		x"ff",	--6154
		x"ff",	--6155
		x"ff",	--6156
		x"ff",	--6157
		x"ff",	--6158
		x"ff",	--6159
		x"ff",	--6160
		x"ff",	--6161
		x"ff",	--6162
		x"ff",	--6163
		x"ff",	--6164
		x"ff",	--6165
		x"ff",	--6166
		x"ff",	--6167
		x"ff",	--6168
		x"ff",	--6169
		x"ff",	--6170
		x"ff",	--6171
		x"ff",	--6172
		x"ff",	--6173
		x"ff",	--6174
		x"ff",	--6175
		x"ff",	--6176
		x"ff",	--6177
		x"ff",	--6178
		x"ff",	--6179
		x"ff",	--6180
		x"ff",	--6181
		x"ff",	--6182
		x"ff",	--6183
		x"ff",	--6184
		x"ff",	--6185
		x"ff",	--6186
		x"ff",	--6187
		x"ff",	--6188
		x"ff",	--6189
		x"ff",	--6190
		x"ff",	--6191
		x"ff",	--6192
		x"ff",	--6193
		x"ff",	--6194
		x"ff",	--6195
		x"ff",	--6196
		x"ff",	--6197
		x"ff",	--6198
		x"ff",	--6199
		x"ff",	--6200
		x"ff",	--6201
		x"ff",	--6202
		x"ff",	--6203
		x"ff",	--6204
		x"ff",	--6205
		x"ff",	--6206
		x"ff",	--6207
		x"ff",	--6208
		x"ff",	--6209
		x"ff",	--6210
		x"ff",	--6211
		x"ff",	--6212
		x"ff",	--6213
		x"ff",	--6214
		x"ff",	--6215
		x"ff",	--6216
		x"ff",	--6217
		x"ff",	--6218
		x"ff",	--6219
		x"ff",	--6220
		x"ff",	--6221
		x"ff",	--6222
		x"ff",	--6223
		x"ff",	--6224
		x"ff",	--6225
		x"ff",	--6226
		x"ff",	--6227
		x"ff",	--6228
		x"ff",	--6229
		x"ff",	--6230
		x"ff",	--6231
		x"ff",	--6232
		x"ff",	--6233
		x"ff",	--6234
		x"ff",	--6235
		x"ff",	--6236
		x"ff",	--6237
		x"ff",	--6238
		x"ff",	--6239
		x"ff",	--6240
		x"ff",	--6241
		x"ff",	--6242
		x"ff",	--6243
		x"ff",	--6244
		x"ff",	--6245
		x"ff",	--6246
		x"ff",	--6247
		x"ff",	--6248
		x"ff",	--6249
		x"ff",	--6250
		x"ff",	--6251
		x"ff",	--6252
		x"ff",	--6253
		x"ff",	--6254
		x"ff",	--6255
		x"ff",	--6256
		x"ff",	--6257
		x"ff",	--6258
		x"ff",	--6259
		x"ff",	--6260
		x"ff",	--6261
		x"ff",	--6262
		x"ff",	--6263
		x"ff",	--6264
		x"ff",	--6265
		x"ff",	--6266
		x"ff",	--6267
		x"ff",	--6268
		x"ff",	--6269
		x"ff",	--6270
		x"ff",	--6271
		x"ff",	--6272
		x"ff",	--6273
		x"ff",	--6274
		x"ff",	--6275
		x"ff",	--6276
		x"ff",	--6277
		x"ff",	--6278
		x"ff",	--6279
		x"ff",	--6280
		x"ff",	--6281
		x"ff",	--6282
		x"ff",	--6283
		x"ff",	--6284
		x"ff",	--6285
		x"ff",	--6286
		x"ff",	--6287
		x"ff",	--6288
		x"ff",	--6289
		x"ff",	--6290
		x"ff",	--6291
		x"ff",	--6292
		x"ff",	--6293
		x"ff",	--6294
		x"ff",	--6295
		x"ff",	--6296
		x"ff",	--6297
		x"ff",	--6298
		x"ff",	--6299
		x"ff",	--6300
		x"ff",	--6301
		x"ff",	--6302
		x"ff",	--6303
		x"ff",	--6304
		x"ff",	--6305
		x"ff",	--6306
		x"ff",	--6307
		x"ff",	--6308
		x"ff",	--6309
		x"ff",	--6310
		x"ff",	--6311
		x"ff",	--6312
		x"ff",	--6313
		x"ff",	--6314
		x"ff",	--6315
		x"ff",	--6316
		x"ff",	--6317
		x"ff",	--6318
		x"ff",	--6319
		x"ff",	--6320
		x"ff",	--6321
		x"ff",	--6322
		x"ff",	--6323
		x"ff",	--6324
		x"ff",	--6325
		x"ff",	--6326
		x"ff",	--6327
		x"ff",	--6328
		x"ff",	--6329
		x"ff",	--6330
		x"ff",	--6331
		x"ff",	--6332
		x"ff",	--6333
		x"ff",	--6334
		x"ff",	--6335
		x"ff",	--6336
		x"ff",	--6337
		x"ff",	--6338
		x"ff",	--6339
		x"ff",	--6340
		x"ff",	--6341
		x"ff",	--6342
		x"ff",	--6343
		x"ff",	--6344
		x"ff",	--6345
		x"ff",	--6346
		x"ff",	--6347
		x"ff",	--6348
		x"ff",	--6349
		x"ff",	--6350
		x"ff",	--6351
		x"ff",	--6352
		x"ff",	--6353
		x"ff",	--6354
		x"ff",	--6355
		x"ff",	--6356
		x"ff",	--6357
		x"ff",	--6358
		x"ff",	--6359
		x"ff",	--6360
		x"ff",	--6361
		x"ff",	--6362
		x"ff",	--6363
		x"ff",	--6364
		x"ff",	--6365
		x"ff",	--6366
		x"ff",	--6367
		x"ff",	--6368
		x"ff",	--6369
		x"ff",	--6370
		x"ff",	--6371
		x"ff",	--6372
		x"ff",	--6373
		x"ff",	--6374
		x"ff",	--6375
		x"ff",	--6376
		x"ff",	--6377
		x"ff",	--6378
		x"ff",	--6379
		x"ff",	--6380
		x"ff",	--6381
		x"ff",	--6382
		x"ff",	--6383
		x"ff",	--6384
		x"ff",	--6385
		x"ff",	--6386
		x"ff",	--6387
		x"ff",	--6388
		x"ff",	--6389
		x"ff",	--6390
		x"ff",	--6391
		x"ff",	--6392
		x"ff",	--6393
		x"ff",	--6394
		x"ff",	--6395
		x"ff",	--6396
		x"ff",	--6397
		x"ff",	--6398
		x"ff",	--6399
		x"ff",	--6400
		x"ff",	--6401
		x"ff",	--6402
		x"ff",	--6403
		x"ff",	--6404
		x"ff",	--6405
		x"ff",	--6406
		x"ff",	--6407
		x"ff",	--6408
		x"ff",	--6409
		x"ff",	--6410
		x"ff",	--6411
		x"ff",	--6412
		x"ff",	--6413
		x"ff",	--6414
		x"ff",	--6415
		x"ff",	--6416
		x"ff",	--6417
		x"ff",	--6418
		x"ff",	--6419
		x"ff",	--6420
		x"ff",	--6421
		x"ff",	--6422
		x"ff",	--6423
		x"ff",	--6424
		x"ff",	--6425
		x"ff",	--6426
		x"ff",	--6427
		x"ff",	--6428
		x"ff",	--6429
		x"ff",	--6430
		x"ff",	--6431
		x"ff",	--6432
		x"ff",	--6433
		x"ff",	--6434
		x"ff",	--6435
		x"ff",	--6436
		x"ff",	--6437
		x"ff",	--6438
		x"ff",	--6439
		x"ff",	--6440
		x"ff",	--6441
		x"ff",	--6442
		x"ff",	--6443
		x"ff",	--6444
		x"ff",	--6445
		x"ff",	--6446
		x"ff",	--6447
		x"ff",	--6448
		x"ff",	--6449
		x"ff",	--6450
		x"ff",	--6451
		x"ff",	--6452
		x"ff",	--6453
		x"ff",	--6454
		x"ff",	--6455
		x"ff",	--6456
		x"ff",	--6457
		x"ff",	--6458
		x"ff",	--6459
		x"ff",	--6460
		x"ff",	--6461
		x"ff",	--6462
		x"ff",	--6463
		x"ff",	--6464
		x"ff",	--6465
		x"ff",	--6466
		x"ff",	--6467
		x"ff",	--6468
		x"ff",	--6469
		x"ff",	--6470
		x"ff",	--6471
		x"ff",	--6472
		x"ff",	--6473
		x"ff",	--6474
		x"ff",	--6475
		x"ff",	--6476
		x"ff",	--6477
		x"ff",	--6478
		x"ff",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"ff",	--6484
		x"ff",	--6485
		x"ff",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"c2",	--8176
		x"c2",	--8177
		x"c2",	--8178
		x"c2",	--8179
		x"c2",	--8180
		x"c2",	--8181
		x"c2",	--8182
		x"cd",	--8183
		x"c9",	--8184
		x"c2",	--8185
		x"c2",	--8186
		x"c2",	--8187
		x"c2",	--8188
		x"c2",	--8189
		x"c2",	--8190
		x"c0");	--8191

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
