library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"4a",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"1a",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"4a",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"b6",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"30",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"4a",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"1a",	--29
		x"f9",	--30
		x"31",	--31
		x"3e",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"d0",	--44
		x"b0",	--45
		x"0c",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"e4",	--50
		x"b0",	--51
		x"94",	--52
		x"21",	--53
		x"3d",	--54
		x"01",	--55
		x"3e",	--56
		x"76",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"3c",	--61
		x"3d",	--62
		x"12",	--63
		x"3e",	--64
		x"4e",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"3c",	--69
		x"3d",	--70
		x"18",	--71
		x"3e",	--72
		x"c2",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"3c",	--77
		x"3d",	--78
		x"1d",	--79
		x"3e",	--80
		x"22",	--81
		x"7f",	--82
		x"61",	--83
		x"b0",	--84
		x"3c",	--85
		x"3d",	--86
		x"24",	--87
		x"3e",	--88
		x"84",	--89
		x"7f",	--90
		x"70",	--91
		x"b0",	--92
		x"3c",	--93
		x"3d",	--94
		x"28",	--95
		x"3e",	--96
		x"c4",	--97
		x"7f",	--98
		x"65",	--99
		x"b0",	--100
		x"3c",	--101
		x"3d",	--102
		x"30",	--103
		x"3e",	--104
		x"54",	--105
		x"7f",	--106
		x"73",	--107
		x"b0",	--108
		x"3c",	--109
		x"3d",	--110
		x"41",	--111
		x"3e",	--112
		x"06",	--113
		x"7f",	--114
		x"7a",	--115
		x"b0",	--116
		x"3c",	--117
		x"3d",	--118
		x"4a",	--119
		x"3e",	--120
		x"7c",	--121
		x"7f",	--122
		x"63",	--123
		x"b0",	--124
		x"3c",	--125
		x"3d",	--126
		x"5e",	--127
		x"3e",	--128
		x"ae",	--129
		x"7f",	--130
		x"6f",	--131
		x"b0",	--132
		x"3c",	--133
		x"3d",	--134
		x"71",	--135
		x"3e",	--136
		x"54",	--137
		x"7f",	--138
		x"74",	--139
		x"b0",	--140
		x"3c",	--141
		x"3d",	--142
		x"76",	--143
		x"3e",	--144
		x"8a",	--145
		x"7f",	--146
		x"62",	--147
		x"b0",	--148
		x"3c",	--149
		x"0e",	--150
		x"0f",	--151
		x"b0",	--152
		x"d2",	--153
		x"2c",	--154
		x"3d",	--155
		x"20",	--156
		x"3e",	--157
		x"80",	--158
		x"0f",	--159
		x"3f",	--160
		x"12",	--161
		x"b0",	--162
		x"da",	--163
		x"0f",	--164
		x"3f",	--165
		x"12",	--166
		x"b0",	--167
		x"22",	--168
		x"2c",	--169
		x"3d",	--170
		x"20",	--171
		x"3e",	--172
		x"88",	--173
		x"0f",	--174
		x"3f",	--175
		x"b0",	--176
		x"da",	--177
		x"0f",	--178
		x"3f",	--179
		x"b0",	--180
		x"22",	--181
		x"0e",	--182
		x"3e",	--183
		x"0f",	--184
		x"3f",	--185
		x"12",	--186
		x"b0",	--187
		x"7a",	--188
		x"3e",	--189
		x"98",	--190
		x"0f",	--191
		x"3f",	--192
		x"06",	--193
		x"b0",	--194
		x"76",	--195
		x"3e",	--196
		x"9c",	--197
		x"0f",	--198
		x"2f",	--199
		x"b0",	--200
		x"76",	--201
		x"0e",	--202
		x"2e",	--203
		x"0f",	--204
		x"3f",	--205
		x"06",	--206
		x"b0",	--207
		x"b0",	--208
		x"0e",	--209
		x"3e",	--210
		x"0f",	--211
		x"3f",	--212
		x"12",	--213
		x"b0",	--214
		x"ba",	--215
		x"b0",	--216
		x"4e",	--217
		x"3e",	--218
		x"a0",	--219
		x"0f",	--220
		x"2f",	--221
		x"b0",	--222
		x"8e",	--223
		x"0f",	--224
		x"2f",	--225
		x"b0",	--226
		x"1c",	--227
		x"3d",	--228
		x"64",	--229
		x"3e",	--230
		x"2a",	--231
		x"0f",	--232
		x"2f",	--233
		x"b0",	--234
		x"a2",	--235
		x"3e",	--236
		x"b0",	--237
		x"0f",	--238
		x"b0",	--239
		x"08",	--240
		x"0f",	--241
		x"b0",	--242
		x"a8",	--243
		x"30",	--244
		x"20",	--245
		x"03",	--246
		x"03",	--247
		x"03",	--248
		x"30",	--249
		x"d1",	--250
		x"30",	--251
		x"17",	--252
		x"30",	--253
		x"1d",	--254
		x"30",	--255
		x"52",	--256
		x"3c",	--257
		x"32",	--258
		x"0d",	--259
		x"3d",	--260
		x"16",	--261
		x"0e",	--262
		x"3e",	--263
		x"22",	--264
		x"0f",	--265
		x"3f",	--266
		x"a4",	--267
		x"b0",	--268
		x"92",	--269
		x"31",	--270
		x"10",	--271
		x"30",	--272
		x"20",	--273
		x"03",	--274
		x"03",	--275
		x"03",	--276
		x"30",	--277
		x"d1",	--278
		x"30",	--279
		x"17",	--280
		x"30",	--281
		x"1d",	--282
		x"30",	--283
		x"52",	--284
		x"3c",	--285
		x"32",	--286
		x"0d",	--287
		x"3d",	--288
		x"14",	--289
		x"0e",	--290
		x"3e",	--291
		x"18",	--292
		x"0f",	--293
		x"3f",	--294
		x"78",	--295
		x"b0",	--296
		x"92",	--297
		x"31",	--298
		x"10",	--299
		x"0e",	--300
		x"3e",	--301
		x"68",	--302
		x"0f",	--303
		x"3f",	--304
		x"94",	--305
		x"b0",	--306
		x"44",	--307
		x"0f",	--308
		x"b0",	--309
		x"4e",	--310
		x"b0",	--311
		x"1c",	--312
		x"30",	--313
		x"b0",	--314
		x"30",	--315
		x"19",	--316
		x"30",	--317
		x"9a",	--318
		x"3d",	--319
		x"8f",	--320
		x"3e",	--321
		x"75",	--322
		x"0f",	--323
		x"3f",	--324
		x"22",	--325
		x"b0",	--326
		x"a8",	--327
		x"31",	--328
		x"06",	--329
		x"0d",	--330
		x"3d",	--331
		x"06",	--332
		x"0e",	--333
		x"2e",	--334
		x"0f",	--335
		x"3f",	--336
		x"1c",	--337
		x"b0",	--338
		x"00",	--339
		x"3e",	--340
		x"64",	--341
		x"0f",	--342
		x"3f",	--343
		x"1c",	--344
		x"b0",	--345
		x"c4",	--346
		x"0f",	--347
		x"3f",	--348
		x"1c",	--349
		x"b0",	--350
		x"00",	--351
		x"0e",	--352
		x"3e",	--353
		x"68",	--354
		x"0f",	--355
		x"3f",	--356
		x"94",	--357
		x"b0",	--358
		x"26",	--359
		x"0f",	--360
		x"b0",	--361
		x"30",	--362
		x"3f",	--363
		x"64",	--364
		x"b0",	--365
		x"36",	--366
		x"f2",	--367
		x"80",	--368
		x"19",	--369
		x"32",	--370
		x"0b",	--371
		x"0a",	--372
		x"05",	--373
		x"1b",	--374
		x"03",	--375
		x"2b",	--376
		x"01",	--377
		x"0b",	--378
		x"b0",	--379
		x"ee",	--380
		x"0f",	--381
		x"fc",	--382
		x"b0",	--383
		x"16",	--384
		x"0b",	--385
		x"3e",	--386
		x"7f",	--387
		x"0d",	--388
		x"06",	--389
		x"7f",	--390
		x"1b",	--391
		x"ed",	--392
		x"7f",	--393
		x"1c",	--394
		x"12",	--395
		x"30",	--396
		x"81",	--397
		x"b0",	--398
		x"94",	--399
		x"21",	--400
		x"3f",	--401
		x"40",	--402
		x"0f",	--403
		x"0a",	--404
		x"ca",	--405
		x"00",	--406
		x"0e",	--407
		x"5f",	--408
		x"40",	--409
		x"b0",	--410
		x"70",	--411
		x"0a",	--412
		x"dd",	--413
		x"0a",	--414
		x"db",	--415
		x"3a",	--416
		x"30",	--417
		x"84",	--418
		x"b0",	--419
		x"94",	--420
		x"21",	--421
		x"d4",	--422
		x"3a",	--423
		x"28",	--424
		x"d1",	--425
		x"82",	--426
		x"1c",	--427
		x"0c",	--428
		x"4e",	--429
		x"8e",	--430
		x"0e",	--431
		x"30",	--432
		x"88",	--433
		x"81",	--434
		x"c4",	--435
		x"b0",	--436
		x"94",	--437
		x"21",	--438
		x"1f",	--439
		x"c0",	--440
		x"3e",	--441
		x"40",	--442
		x"0e",	--443
		x"0e",	--444
		x"ce",	--445
		x"00",	--446
		x"1a",	--447
		x"ba",	--448
		x"1b",	--449
		x"04",	--450
		x"7f",	--451
		x"5b",	--452
		x"b5",	--453
		x"b1",	--454
		x"2b",	--455
		x"b2",	--456
		x"7f",	--457
		x"42",	--458
		x"17",	--459
		x"7f",	--460
		x"43",	--461
		x"04",	--462
		x"7f",	--463
		x"41",	--464
		x"a8",	--465
		x"07",	--466
		x"7f",	--467
		x"43",	--468
		x"16",	--469
		x"7f",	--470
		x"44",	--471
		x"a1",	--472
		x"1b",	--473
		x"30",	--474
		x"8b",	--475
		x"b0",	--476
		x"94",	--477
		x"21",	--478
		x"b0",	--479
		x"dc",	--480
		x"0b",	--481
		x"98",	--482
		x"30",	--483
		x"90",	--484
		x"b0",	--485
		x"94",	--486
		x"21",	--487
		x"b0",	--488
		x"04",	--489
		x"0b",	--490
		x"8f",	--491
		x"30",	--492
		x"97",	--493
		x"b0",	--494
		x"94",	--495
		x"21",	--496
		x"b0",	--497
		x"2c",	--498
		x"0b",	--499
		x"86",	--500
		x"30",	--501
		x"9f",	--502
		x"b0",	--503
		x"94",	--504
		x"21",	--505
		x"b0",	--506
		x"54",	--507
		x"0b",	--508
		x"7d",	--509
		x"30",	--510
		x"b0",	--511
		x"82",	--512
		x"36",	--513
		x"30",	--514
		x"0b",	--515
		x"1b",	--516
		x"36",	--517
		x"0c",	--518
		x"3d",	--519
		x"7a",	--520
		x"1e",	--521
		x"12",	--522
		x"1f",	--523
		x"14",	--524
		x"b0",	--525
		x"b2",	--526
		x"b0",	--527
		x"5c",	--528
		x"0e",	--529
		x"0c",	--530
		x"3d",	--531
		x"7a",	--532
		x"1e",	--533
		x"0e",	--534
		x"1f",	--535
		x"10",	--536
		x"b0",	--537
		x"b2",	--538
		x"b0",	--539
		x"5c",	--540
		x"0e",	--541
		x"0c",	--542
		x"3d",	--543
		x"7a",	--544
		x"1e",	--545
		x"0a",	--546
		x"1f",	--547
		x"0c",	--548
		x"b0",	--549
		x"b2",	--550
		x"b0",	--551
		x"5c",	--552
		x"0e",	--553
		x"30",	--554
		x"b8",	--555
		x"30",	--556
		x"38",	--557
		x"b0",	--558
		x"44",	--559
		x"31",	--560
		x"0a",	--561
		x"30",	--562
		x"38",	--563
		x"30",	--564
		x"c7",	--565
		x"b0",	--566
		x"94",	--567
		x"21",	--568
		x"0f",	--569
		x"3b",	--570
		x"30",	--571
		x"0b",	--572
		x"0b",	--573
		x"0e",	--574
		x"1f",	--575
		x"36",	--576
		x"b0",	--577
		x"18",	--578
		x"0f",	--579
		x"30",	--580
		x"cc",	--581
		x"b0",	--582
		x"94",	--583
		x"21",	--584
		x"1b",	--585
		x"3b",	--586
		x"05",	--587
		x"f1",	--588
		x"30",	--589
		x"d0",	--590
		x"b0",	--591
		x"94",	--592
		x"21",	--593
		x"3b",	--594
		x"30",	--595
		x"82",	--596
		x"36",	--597
		x"30",	--598
		x"0b",	--599
		x"21",	--600
		x"0b",	--601
		x"81",	--602
		x"00",	--603
		x"1f",	--604
		x"14",	--605
		x"b2",	--606
		x"00",	--607
		x"25",	--608
		x"92",	--609
		x"1a",	--610
		x"0e",	--611
		x"1f",	--612
		x"02",	--613
		x"b0",	--614
		x"b8",	--615
		x"0d",	--616
		x"0e",	--617
		x"1f",	--618
		x"00",	--619
		x"b0",	--620
		x"a2",	--621
		x"0f",	--622
		x"21",	--623
		x"3b",	--624
		x"30",	--625
		x"82",	--626
		x"1a",	--627
		x"0a",	--628
		x"82",	--629
		x"1a",	--630
		x"1f",	--631
		x"00",	--632
		x"b0",	--633
		x"ca",	--634
		x"0f",	--635
		x"21",	--636
		x"3b",	--637
		x"30",	--638
		x"0f",	--639
		x"b0",	--640
		x"78",	--641
		x"0f",	--642
		x"21",	--643
		x"3b",	--644
		x"30",	--645
		x"0e",	--646
		x"3f",	--647
		x"78",	--648
		x"b0",	--649
		x"5e",	--650
		x"82",	--651
		x"00",	--652
		x"d3",	--653
		x"82",	--654
		x"78",	--655
		x"30",	--656
		x"0b",	--657
		x"0a",	--658
		x"21",	--659
		x"0a",	--660
		x"0b",	--661
		x"2f",	--662
		x"1b",	--663
		x"0e",	--664
		x"1f",	--665
		x"02",	--666
		x"b0",	--667
		x"b8",	--668
		x"0d",	--669
		x"2a",	--670
		x"18",	--671
		x"0e",	--672
		x"1f",	--673
		x"04",	--674
		x"81",	--675
		x"02",	--676
		x"b0",	--677
		x"b8",	--678
		x"0e",	--679
		x"1d",	--680
		x"02",	--681
		x"1f",	--682
		x"78",	--683
		x"b0",	--684
		x"a2",	--685
		x"0f",	--686
		x"21",	--687
		x"3a",	--688
		x"3b",	--689
		x"30",	--690
		x"3d",	--691
		x"64",	--692
		x"3e",	--693
		x"2a",	--694
		x"f2",	--695
		x"3e",	--696
		x"2a",	--697
		x"ef",	--698
		x"1f",	--699
		x"82",	--700
		x"1c",	--701
		x"01",	--702
		x"0f",	--703
		x"82",	--704
		x"1c",	--705
		x"0f",	--706
		x"30",	--707
		x"5e",	--708
		x"19",	--709
		x"4e",	--710
		x"0f",	--711
		x"03",	--712
		x"c2",	--713
		x"19",	--714
		x"30",	--715
		x"c2",	--716
		x"19",	--717
		x"30",	--718
		x"1e",	--719
		x"1e",	--720
		x"3e",	--721
		x"06",	--722
		x"0f",	--723
		x"0f",	--724
		x"10",	--725
		x"d4",	--726
		x"c2",	--727
		x"19",	--728
		x"3e",	--729
		x"07",	--730
		x"03",	--731
		x"82",	--732
		x"1e",	--733
		x"30",	--734
		x"1e",	--735
		x"82",	--736
		x"1e",	--737
		x"30",	--738
		x"f2",	--739
		x"0e",	--740
		x"19",	--741
		x"f2",	--742
		x"f2",	--743
		x"0a",	--744
		x"19",	--745
		x"ee",	--746
		x"e2",	--747
		x"19",	--748
		x"eb",	--749
		x"f2",	--750
		x"0d",	--751
		x"19",	--752
		x"e7",	--753
		x"f2",	--754
		x"09",	--755
		x"19",	--756
		x"e3",	--757
		x"f2",	--758
		x"03",	--759
		x"19",	--760
		x"df",	--761
		x"f2",	--762
		x"07",	--763
		x"19",	--764
		x"db",	--765
		x"0e",	--766
		x"1f",	--767
		x"7c",	--768
		x"b0",	--769
		x"26",	--770
		x"0e",	--771
		x"1f",	--772
		x"7a",	--773
		x"b0",	--774
		x"26",	--775
		x"30",	--776
		x"a6",	--777
		x"b0",	--778
		x"94",	--779
		x"21",	--780
		x"30",	--781
		x"b2",	--782
		x"02",	--783
		x"09",	--784
		x"1f",	--785
		x"7c",	--786
		x"b0",	--787
		x"e2",	--788
		x"1f",	--789
		x"7a",	--790
		x"b0",	--791
		x"e2",	--792
		x"30",	--793
		x"0e",	--794
		x"3f",	--795
		x"fc",	--796
		x"b0",	--797
		x"5e",	--798
		x"82",	--799
		x"02",	--800
		x"ef",	--801
		x"82",	--802
		x"7c",	--803
		x"82",	--804
		x"7a",	--805
		x"30",	--806
		x"82",	--807
		x"7e",	--808
		x"30",	--809
		x"0b",	--810
		x"0a",	--811
		x"21",	--812
		x"0b",	--813
		x"3f",	--814
		x"03",	--815
		x"30",	--816
		x"23",	--817
		x"0e",	--818
		x"1f",	--819
		x"02",	--820
		x"b0",	--821
		x"86",	--822
		x"0a",	--823
		x"0e",	--824
		x"1f",	--825
		x"04",	--826
		x"b0",	--827
		x"86",	--828
		x"0b",	--829
		x"0f",	--830
		x"0a",	--831
		x"30",	--832
		x"dd",	--833
		x"b0",	--834
		x"94",	--835
		x"31",	--836
		x"06",	--837
		x"0e",	--838
		x"1f",	--839
		x"7c",	--840
		x"b0",	--841
		x"26",	--842
		x"0e",	--843
		x"1f",	--844
		x"7a",	--845
		x"b0",	--846
		x"26",	--847
		x"0f",	--848
		x"21",	--849
		x"3a",	--850
		x"3b",	--851
		x"30",	--852
		x"0e",	--853
		x"1f",	--854
		x"06",	--855
		x"b0",	--856
		x"b8",	--857
		x"1d",	--858
		x"0e",	--859
		x"1f",	--860
		x"02",	--861
		x"b0",	--862
		x"a2",	--863
		x"d1",	--864
		x"30",	--865
		x"ad",	--866
		x"b0",	--867
		x"94",	--868
		x"a1",	--869
		x"00",	--870
		x"30",	--871
		x"be",	--872
		x"b0",	--873
		x"94",	--874
		x"21",	--875
		x"3f",	--876
		x"e3",	--877
		x"3e",	--878
		x"64",	--879
		x"1f",	--880
		x"7c",	--881
		x"b0",	--882
		x"26",	--883
		x"3e",	--884
		x"9c",	--885
		x"1f",	--886
		x"7a",	--887
		x"b0",	--888
		x"26",	--889
		x"1d",	--890
		x"3e",	--891
		x"c8",	--892
		x"1f",	--893
		x"02",	--894
		x"b0",	--895
		x"a2",	--896
		x"30",	--897
		x"3e",	--898
		x"9c",	--899
		x"1f",	--900
		x"7c",	--901
		x"b0",	--902
		x"26",	--903
		x"3e",	--904
		x"64",	--905
		x"1f",	--906
		x"7a",	--907
		x"b0",	--908
		x"26",	--909
		x"1d",	--910
		x"3e",	--911
		x"c8",	--912
		x"1f",	--913
		x"02",	--914
		x"b0",	--915
		x"a2",	--916
		x"30",	--917
		x"3e",	--918
		x"c4",	--919
		x"1f",	--920
		x"7c",	--921
		x"b0",	--922
		x"26",	--923
		x"3e",	--924
		x"c4",	--925
		x"1f",	--926
		x"7a",	--927
		x"b0",	--928
		x"26",	--929
		x"1d",	--930
		x"3e",	--931
		x"c8",	--932
		x"1f",	--933
		x"02",	--934
		x"b0",	--935
		x"a2",	--936
		x"30",	--937
		x"3e",	--938
		x"3c",	--939
		x"1f",	--940
		x"7c",	--941
		x"b0",	--942
		x"26",	--943
		x"3e",	--944
		x"3c",	--945
		x"1f",	--946
		x"7a",	--947
		x"b0",	--948
		x"26",	--949
		x"1d",	--950
		x"3e",	--951
		x"c8",	--952
		x"1f",	--953
		x"02",	--954
		x"b0",	--955
		x"a2",	--956
		x"30",	--957
		x"30",	--958
		x"e5",	--959
		x"b0",	--960
		x"94",	--961
		x"21",	--962
		x"0f",	--963
		x"30",	--964
		x"b2",	--965
		x"00",	--966
		x"92",	--967
		x"b2",	--968
		x"30",	--969
		x"94",	--970
		x"b2",	--971
		x"41",	--972
		x"96",	--973
		x"30",	--974
		x"fb",	--975
		x"b0",	--976
		x"94",	--977
		x"92",	--978
		x"90",	--979
		x"b1",	--980
		x"19",	--981
		x"00",	--982
		x"b0",	--983
		x"94",	--984
		x"21",	--985
		x"0f",	--986
		x"30",	--987
		x"0b",	--988
		x"0a",	--989
		x"8e",	--990
		x"00",	--991
		x"6d",	--992
		x"4d",	--993
		x"5e",	--994
		x"1f",	--995
		x"0a",	--996
		x"0c",	--997
		x"0f",	--998
		x"7b",	--999
		x"0a",	--1000
		x"2b",	--1001
		x"0c",	--1002
		x"0c",	--1003
		x"0c",	--1004
		x"0c",	--1005
		x"8d",	--1006
		x"0c",	--1007
		x"3c",	--1008
		x"d0",	--1009
		x"1a",	--1010
		x"7d",	--1011
		x"4d",	--1012
		x"17",	--1013
		x"7d",	--1014
		x"78",	--1015
		x"1a",	--1016
		x"4b",	--1017
		x"7b",	--1018
		x"d0",	--1019
		x"0a",	--1020
		x"e9",	--1021
		x"7b",	--1022
		x"0a",	--1023
		x"34",	--1024
		x"0c",	--1025
		x"0b",	--1026
		x"0b",	--1027
		x"0b",	--1028
		x"0c",	--1029
		x"8d",	--1030
		x"0c",	--1031
		x"3c",	--1032
		x"d0",	--1033
		x"7d",	--1034
		x"4d",	--1035
		x"e9",	--1036
		x"9e",	--1037
		x"00",	--1038
		x"0f",	--1039
		x"3a",	--1040
		x"3b",	--1041
		x"30",	--1042
		x"1a",	--1043
		x"de",	--1044
		x"4b",	--1045
		x"7b",	--1046
		x"9f",	--1047
		x"7b",	--1048
		x"06",	--1049
		x"0a",	--1050
		x"0c",	--1051
		x"0c",	--1052
		x"0c",	--1053
		x"0c",	--1054
		x"8d",	--1055
		x"0c",	--1056
		x"3c",	--1057
		x"a9",	--1058
		x"1a",	--1059
		x"ce",	--1060
		x"4b",	--1061
		x"7b",	--1062
		x"bf",	--1063
		x"7b",	--1064
		x"06",	--1065
		x"0a",	--1066
		x"0c",	--1067
		x"0c",	--1068
		x"0c",	--1069
		x"0c",	--1070
		x"8d",	--1071
		x"0c",	--1072
		x"3c",	--1073
		x"c9",	--1074
		x"1a",	--1075
		x"be",	--1076
		x"8d",	--1077
		x"0d",	--1078
		x"30",	--1079
		x"32",	--1080
		x"b0",	--1081
		x"94",	--1082
		x"21",	--1083
		x"0c",	--1084
		x"0f",	--1085
		x"3a",	--1086
		x"3b",	--1087
		x"30",	--1088
		x"0c",	--1089
		x"ca",	--1090
		x"0b",	--1091
		x"0a",	--1092
		x"8e",	--1093
		x"00",	--1094
		x"6b",	--1095
		x"4b",	--1096
		x"37",	--1097
		x"1f",	--1098
		x"1a",	--1099
		x"0c",	--1100
		x"12",	--1101
		x"4d",	--1102
		x"7d",	--1103
		x"d0",	--1104
		x"7d",	--1105
		x"0a",	--1106
		x"22",	--1107
		x"0c",	--1108
		x"0d",	--1109
		x"0d",	--1110
		x"0d",	--1111
		x"0c",	--1112
		x"8b",	--1113
		x"0c",	--1114
		x"3c",	--1115
		x"d0",	--1116
		x"7b",	--1117
		x"4b",	--1118
		x"07",	--1119
		x"7b",	--1120
		x"2d",	--1121
		x"eb",	--1122
		x"3a",	--1123
		x"7b",	--1124
		x"4b",	--1125
		x"f9",	--1126
		x"02",	--1127
		x"32",	--1128
		x"03",	--1129
		x"82",	--1130
		x"32",	--1131
		x"82",	--1132
		x"38",	--1133
		x"1f",	--1134
		x"3a",	--1135
		x"32",	--1136
		x"9e",	--1137
		x"00",	--1138
		x"3a",	--1139
		x"3b",	--1140
		x"30",	--1141
		x"8b",	--1142
		x"0b",	--1143
		x"30",	--1144
		x"32",	--1145
		x"b0",	--1146
		x"94",	--1147
		x"21",	--1148
		x"0f",	--1149
		x"3a",	--1150
		x"3b",	--1151
		x"30",	--1152
		x"0f",	--1153
		x"ee",	--1154
		x"0b",	--1155
		x"0a",	--1156
		x"09",	--1157
		x"09",	--1158
		x"1f",	--1159
		x"22",	--1160
		x"b0",	--1161
		x"7e",	--1162
		x"0a",	--1163
		x"0b",	--1164
		x"1e",	--1165
		x"24",	--1166
		x"1f",	--1167
		x"26",	--1168
		x"b0",	--1169
		x"b6",	--1170
		x"89",	--1171
		x"24",	--1172
		x"89",	--1173
		x"26",	--1174
		x"0d",	--1175
		x"0e",	--1176
		x"0f",	--1177
		x"b0",	--1178
		x"30",	--1179
		x"0c",	--1180
		x"3d",	--1181
		x"00",	--1182
		x"b0",	--1183
		x"16",	--1184
		x"0a",	--1185
		x"0b",	--1186
		x"3c",	--1187
		x"66",	--1188
		x"3d",	--1189
		x"66",	--1190
		x"b0",	--1191
		x"76",	--1192
		x"0f",	--1193
		x"01",	--1194
		x"18",	--1195
		x"3c",	--1196
		x"cd",	--1197
		x"3d",	--1198
		x"cc",	--1199
		x"0e",	--1200
		x"0f",	--1201
		x"b0",	--1202
		x"16",	--1203
		x"0f",	--1204
		x"04",	--1205
		x"3a",	--1206
		x"cd",	--1207
		x"3b",	--1208
		x"cc",	--1209
		x"0d",	--1210
		x"0e",	--1211
		x"1f",	--1212
		x"20",	--1213
		x"b0",	--1214
		x"76",	--1215
		x"39",	--1216
		x"3a",	--1217
		x"3b",	--1218
		x"30",	--1219
		x"3a",	--1220
		x"66",	--1221
		x"3b",	--1222
		x"66",	--1223
		x"f1",	--1224
		x"0b",	--1225
		x"0a",	--1226
		x"0b",	--1227
		x"0a",	--1228
		x"8f",	--1229
		x"20",	--1230
		x"8f",	--1231
		x"22",	--1232
		x"11",	--1233
		x"16",	--1234
		x"11",	--1235
		x"16",	--1236
		x"11",	--1237
		x"16",	--1238
		x"11",	--1239
		x"16",	--1240
		x"11",	--1241
		x"16",	--1242
		x"11",	--1243
		x"16",	--1244
		x"1d",	--1245
		x"12",	--1246
		x"1e",	--1247
		x"14",	--1248
		x"b0",	--1249
		x"96",	--1250
		x"31",	--1251
		x"0c",	--1252
		x"8b",	--1253
		x"28",	--1254
		x"0e",	--1255
		x"3f",	--1256
		x"06",	--1257
		x"b0",	--1258
		x"5e",	--1259
		x"8b",	--1260
		x"2a",	--1261
		x"3a",	--1262
		x"3b",	--1263
		x"30",	--1264
		x"0b",	--1265
		x"0b",	--1266
		x"1f",	--1267
		x"22",	--1268
		x"b0",	--1269
		x"7e",	--1270
		x"8b",	--1271
		x"24",	--1272
		x"8b",	--1273
		x"26",	--1274
		x"0d",	--1275
		x"1e",	--1276
		x"28",	--1277
		x"1f",	--1278
		x"2a",	--1279
		x"b0",	--1280
		x"a2",	--1281
		x"3b",	--1282
		x"30",	--1283
		x"0b",	--1284
		x"0b",	--1285
		x"0d",	--1286
		x"3e",	--1287
		x"00",	--1288
		x"1f",	--1289
		x"20",	--1290
		x"b0",	--1291
		x"76",	--1292
		x"1f",	--1293
		x"2a",	--1294
		x"b0",	--1295
		x"ca",	--1296
		x"3b",	--1297
		x"30",	--1298
		x"0b",	--1299
		x"0b",	--1300
		x"0d",	--1301
		x"8d",	--1302
		x"8d",	--1303
		x"8d",	--1304
		x"8d",	--1305
		x"0f",	--1306
		x"b0",	--1307
		x"b6",	--1308
		x"0d",	--1309
		x"0e",	--1310
		x"0f",	--1311
		x"b0",	--1312
		x"1c",	--1313
		x"3b",	--1314
		x"30",	--1315
		x"0b",	--1316
		x"0a",	--1317
		x"0a",	--1318
		x"3b",	--1319
		x"00",	--1320
		x"0d",	--1321
		x"0e",	--1322
		x"1f",	--1323
		x"82",	--1324
		x"b0",	--1325
		x"76",	--1326
		x"0d",	--1327
		x"0e",	--1328
		x"1f",	--1329
		x"80",	--1330
		x"b0",	--1331
		x"76",	--1332
		x"30",	--1333
		x"47",	--1334
		x"b0",	--1335
		x"94",	--1336
		x"21",	--1337
		x"3a",	--1338
		x"3b",	--1339
		x"30",	--1340
		x"82",	--1341
		x"82",	--1342
		x"82",	--1343
		x"80",	--1344
		x"30",	--1345
		x"0b",	--1346
		x"0a",	--1347
		x"21",	--1348
		x"0a",	--1349
		x"0b",	--1350
		x"b2",	--1351
		x"04",	--1352
		x"4e",	--1353
		x"3a",	--1354
		x"03",	--1355
		x"53",	--1356
		x"3e",	--1357
		x"0e",	--1358
		x"1f",	--1359
		x"02",	--1360
		x"b0",	--1361
		x"b8",	--1362
		x"0a",	--1363
		x"0e",	--1364
		x"1f",	--1365
		x"04",	--1366
		x"b0",	--1367
		x"b8",	--1368
		x"0b",	--1369
		x"0f",	--1370
		x"0a",	--1371
		x"30",	--1372
		x"94",	--1373
		x"b0",	--1374
		x"94",	--1375
		x"31",	--1376
		x"06",	--1377
		x"0e",	--1378
		x"0f",	--1379
		x"b0",	--1380
		x"ec",	--1381
		x"0c",	--1382
		x"3d",	--1383
		x"c8",	--1384
		x"b0",	--1385
		x"d6",	--1386
		x"0c",	--1387
		x"0d",	--1388
		x"0e",	--1389
		x"3f",	--1390
		x"80",	--1391
		x"b0",	--1392
		x"62",	--1393
		x"0d",	--1394
		x"0e",	--1395
		x"1f",	--1396
		x"82",	--1397
		x"b0",	--1398
		x"76",	--1399
		x"0e",	--1400
		x"0f",	--1401
		x"b0",	--1402
		x"ec",	--1403
		x"0c",	--1404
		x"3d",	--1405
		x"c8",	--1406
		x"b0",	--1407
		x"d6",	--1408
		x"0d",	--1409
		x"0e",	--1410
		x"1f",	--1411
		x"80",	--1412
		x"b0",	--1413
		x"76",	--1414
		x"0f",	--1415
		x"21",	--1416
		x"3a",	--1417
		x"3b",	--1418
		x"30",	--1419
		x"0e",	--1420
		x"1f",	--1421
		x"06",	--1422
		x"b0",	--1423
		x"b8",	--1424
		x"1d",	--1425
		x"0e",	--1426
		x"1f",	--1427
		x"04",	--1428
		x"b0",	--1429
		x"a2",	--1430
		x"b6",	--1431
		x"0e",	--1432
		x"3f",	--1433
		x"48",	--1434
		x"b0",	--1435
		x"5e",	--1436
		x"82",	--1437
		x"04",	--1438
		x"aa",	--1439
		x"30",	--1440
		x"4e",	--1441
		x"b0",	--1442
		x"94",	--1443
		x"b1",	--1444
		x"68",	--1445
		x"00",	--1446
		x"b0",	--1447
		x"94",	--1448
		x"a1",	--1449
		x"00",	--1450
		x"30",	--1451
		x"79",	--1452
		x"b0",	--1453
		x"94",	--1454
		x"21",	--1455
		x"3f",	--1456
		x"d6",	--1457
		x"0b",	--1458
		x"0a",	--1459
		x"1f",	--1460
		x"86",	--1461
		x"b0",	--1462
		x"7e",	--1463
		x"0a",	--1464
		x"0b",	--1465
		x"1f",	--1466
		x"84",	--1467
		x"b0",	--1468
		x"7e",	--1469
		x"0b",	--1470
		x"0a",	--1471
		x"3e",	--1472
		x"3f",	--1473
		x"1e",	--1474
		x"0f",	--1475
		x"0f",	--1476
		x"0e",	--1477
		x"30",	--1478
		x"9c",	--1479
		x"30",	--1480
		x"38",	--1481
		x"b0",	--1482
		x"44",	--1483
		x"31",	--1484
		x"0c",	--1485
		x"30",	--1486
		x"38",	--1487
		x"30",	--1488
		x"a4",	--1489
		x"b0",	--1490
		x"94",	--1491
		x"21",	--1492
		x"3a",	--1493
		x"3b",	--1494
		x"30",	--1495
		x"82",	--1496
		x"84",	--1497
		x"82",	--1498
		x"86",	--1499
		x"30",	--1500
		x"82",	--1501
		x"82",	--1502
		x"82",	--1503
		x"80",	--1504
		x"30",	--1505
		x"0b",	--1506
		x"0a",	--1507
		x"09",	--1508
		x"08",	--1509
		x"21",	--1510
		x"0a",	--1511
		x"0b",	--1512
		x"81",	--1513
		x"00",	--1514
		x"1f",	--1515
		x"1c",	--1516
		x"b2",	--1517
		x"06",	--1518
		x"6f",	--1519
		x"92",	--1520
		x"20",	--1521
		x"0e",	--1522
		x"1f",	--1523
		x"02",	--1524
		x"b0",	--1525
		x"b8",	--1526
		x"08",	--1527
		x"3a",	--1528
		x"03",	--1529
		x"1e",	--1530
		x"09",	--1531
		x"0d",	--1532
		x"0e",	--1533
		x"1f",	--1534
		x"06",	--1535
		x"b0",	--1536
		x"a2",	--1537
		x"0f",	--1538
		x"21",	--1539
		x"38",	--1540
		x"39",	--1541
		x"3a",	--1542
		x"3b",	--1543
		x"30",	--1544
		x"82",	--1545
		x"20",	--1546
		x"49",	--1547
		x"82",	--1548
		x"20",	--1549
		x"1f",	--1550
		x"06",	--1551
		x"b0",	--1552
		x"ca",	--1553
		x"0f",	--1554
		x"21",	--1555
		x"38",	--1556
		x"39",	--1557
		x"3a",	--1558
		x"3b",	--1559
		x"30",	--1560
		x"0e",	--1561
		x"1f",	--1562
		x"04",	--1563
		x"b0",	--1564
		x"b8",	--1565
		x"09",	--1566
		x"3a",	--1567
		x"05",	--1568
		x"da",	--1569
		x"0e",	--1570
		x"1f",	--1571
		x"06",	--1572
		x"b0",	--1573
		x"b8",	--1574
		x"0a",	--1575
		x"0e",	--1576
		x"1f",	--1577
		x"08",	--1578
		x"b0",	--1579
		x"b8",	--1580
		x"0b",	--1581
		x"0f",	--1582
		x"0a",	--1583
		x"30",	--1584
		x"a9",	--1585
		x"b0",	--1586
		x"94",	--1587
		x"31",	--1588
		x"06",	--1589
		x"0e",	--1590
		x"0f",	--1591
		x"b0",	--1592
		x"ec",	--1593
		x"0c",	--1594
		x"3d",	--1595
		x"c8",	--1596
		x"b0",	--1597
		x"d6",	--1598
		x"0d",	--1599
		x"0e",	--1600
		x"1f",	--1601
		x"82",	--1602
		x"b0",	--1603
		x"76",	--1604
		x"0e",	--1605
		x"0f",	--1606
		x"b0",	--1607
		x"ec",	--1608
		x"0c",	--1609
		x"3d",	--1610
		x"c8",	--1611
		x"b0",	--1612
		x"d6",	--1613
		x"0d",	--1614
		x"0e",	--1615
		x"1f",	--1616
		x"80",	--1617
		x"b0",	--1618
		x"76",	--1619
		x"a7",	--1620
		x"0f",	--1621
		x"b0",	--1622
		x"64",	--1623
		x"0f",	--1624
		x"21",	--1625
		x"38",	--1626
		x"39",	--1627
		x"3a",	--1628
		x"3b",	--1629
		x"30",	--1630
		x"0e",	--1631
		x"3f",	--1632
		x"64",	--1633
		x"b0",	--1634
		x"5e",	--1635
		x"82",	--1636
		x"06",	--1637
		x"89",	--1638
		x"0b",	--1639
		x"0a",	--1640
		x"09",	--1641
		x"08",	--1642
		x"08",	--1643
		x"3a",	--1644
		x"08",	--1645
		x"09",	--1646
		x"0b",	--1647
		x"0e",	--1648
		x"0f",	--1649
		x"b0",	--1650
		x"18",	--1651
		x"2f",	--1652
		x"09",	--1653
		x"1e",	--1654
		x"4d",	--1655
		x"7d",	--1656
		x"0f",	--1657
		x"03",	--1658
		x"0e",	--1659
		x"7d",	--1660
		x"fd",	--1661
		x"09",	--1662
		x"1b",	--1663
		x"2a",	--1664
		x"3b",	--1665
		x"05",	--1666
		x"ec",	--1667
		x"0f",	--1668
		x"38",	--1669
		x"39",	--1670
		x"3a",	--1671
		x"3b",	--1672
		x"30",	--1673
		x"0b",	--1674
		x"0a",	--1675
		x"82",	--1676
		x"26",	--1677
		x"03",	--1678
		x"3a",	--1679
		x"3b",	--1680
		x"30",	--1681
		x"1f",	--1682
		x"7e",	--1683
		x"b0",	--1684
		x"ce",	--1685
		x"0a",	--1686
		x"0b",	--1687
		x"0e",	--1688
		x"1f",	--1689
		x"7e",	--1690
		x"b0",	--1691
		x"18",	--1692
		x"0f",	--1693
		x"30",	--1694
		x"b1",	--1695
		x"b0",	--1696
		x"94",	--1697
		x"21",	--1698
		x"1b",	--1699
		x"3b",	--1700
		x"05",	--1701
		x"f1",	--1702
		x"30",	--1703
		x"b5",	--1704
		x"b0",	--1705
		x"94",	--1706
		x"21",	--1707
		x"1f",	--1708
		x"28",	--1709
		x"0f",	--1710
		x"23",	--1711
		x"0a",	--1712
		x"75",	--1713
		x"3a",	--1714
		x"18",	--1715
		x"7f",	--1716
		x"2a",	--1717
		x"83",	--1718
		x"1a",	--1719
		x"99",	--1720
		x"2a",	--1721
		x"47",	--1722
		x"a2",	--1723
		x"28",	--1724
		x"0e",	--1725
		x"1f",	--1726
		x"7c",	--1727
		x"b0",	--1728
		x"26",	--1729
		x"0e",	--1730
		x"1f",	--1731
		x"7a",	--1732
		x"b0",	--1733
		x"26",	--1734
		x"b2",	--1735
		x"14",	--1736
		x"24",	--1737
		x"b2",	--1738
		x"0f",	--1739
		x"22",	--1740
		x"30",	--1741
		x"00",	--1742
		x"b0",	--1743
		x"94",	--1744
		x"21",	--1745
		x"bc",	--1746
		x"82",	--1747
		x"24",	--1748
		x"12",	--1749
		x"1e",	--1750
		x"22",	--1751
		x"0e",	--1752
		x"0b",	--1753
		x"1f",	--1754
		x"8f",	--1755
		x"2f",	--1756
		x"a1",	--1757
		x"3f",	--1758
		x"03",	--1759
		x"32",	--1760
		x"3e",	--1761
		x"82",	--1762
		x"22",	--1763
		x"aa",	--1764
		x"82",	--1765
		x"28",	--1766
		x"a7",	--1767
		x"0e",	--1768
		x"1f",	--1769
		x"7c",	--1770
		x"b0",	--1771
		x"26",	--1772
		x"0e",	--1773
		x"1f",	--1774
		x"7a",	--1775
		x"b0",	--1776
		x"26",	--1777
		x"30",	--1778
		x"16",	--1779
		x"b0",	--1780
		x"94",	--1781
		x"21",	--1782
		x"b2",	--1783
		x"24",	--1784
		x"0a",	--1785
		x"94",	--1786
		x"82",	--1787
		x"24",	--1788
		x"82",	--1789
		x"22",	--1790
		x"82",	--1791
		x"28",	--1792
		x"8d",	--1793
		x"0e",	--1794
		x"1f",	--1795
		x"7c",	--1796
		x"b0",	--1797
		x"26",	--1798
		x"0e",	--1799
		x"1f",	--1800
		x"7a",	--1801
		x"b0",	--1802
		x"26",	--1803
		x"0a",	--1804
		x"30",	--1805
		x"11",	--1806
		x"b0",	--1807
		x"94",	--1808
		x"21",	--1809
		x"7c",	--1810
		x"3e",	--1811
		x"1e",	--1812
		x"1f",	--1813
		x"7c",	--1814
		x"b0",	--1815
		x"26",	--1816
		x"3e",	--1817
		x"1e",	--1818
		x"1f",	--1819
		x"7a",	--1820
		x"b0",	--1821
		x"26",	--1822
		x"30",	--1823
		x"3e",	--1824
		x"b0",	--1825
		x"94",	--1826
		x"21",	--1827
		x"1e",	--1828
		x"22",	--1829
		x"ba",	--1830
		x"3e",	--1831
		x"3c",	--1832
		x"1f",	--1833
		x"7c",	--1834
		x"b0",	--1835
		x"26",	--1836
		x"3e",	--1837
		x"c4",	--1838
		x"1f",	--1839
		x"7a",	--1840
		x"b0",	--1841
		x"26",	--1842
		x"5b",	--1843
		x"30",	--1844
		x"b8",	--1845
		x"b0",	--1846
		x"94",	--1847
		x"21",	--1848
		x"55",	--1849
		x"92",	--1850
		x"28",	--1851
		x"0e",	--1852
		x"1f",	--1853
		x"7c",	--1854
		x"b0",	--1855
		x"26",	--1856
		x"0e",	--1857
		x"1f",	--1858
		x"7a",	--1859
		x"b0",	--1860
		x"26",	--1861
		x"b2",	--1862
		x"14",	--1863
		x"24",	--1864
		x"b2",	--1865
		x"14",	--1866
		x"22",	--1867
		x"30",	--1868
		x"e0",	--1869
		x"b0",	--1870
		x"94",	--1871
		x"21",	--1872
		x"3d",	--1873
		x"b2",	--1874
		x"03",	--1875
		x"28",	--1876
		x"0e",	--1877
		x"1f",	--1878
		x"7c",	--1879
		x"b0",	--1880
		x"26",	--1881
		x"0e",	--1882
		x"1f",	--1883
		x"7a",	--1884
		x"b0",	--1885
		x"26",	--1886
		x"b2",	--1887
		x"14",	--1888
		x"24",	--1889
		x"b2",	--1890
		x"0f",	--1891
		x"22",	--1892
		x"30",	--1893
		x"ee",	--1894
		x"b0",	--1895
		x"94",	--1896
		x"21",	--1897
		x"24",	--1898
		x"3e",	--1899
		x"1e",	--1900
		x"1f",	--1901
		x"7c",	--1902
		x"b0",	--1903
		x"26",	--1904
		x"3e",	--1905
		x"1e",	--1906
		x"1f",	--1907
		x"7a",	--1908
		x"b0",	--1909
		x"26",	--1910
		x"30",	--1911
		x"1d",	--1912
		x"b0",	--1913
		x"94",	--1914
		x"21",	--1915
		x"1e",	--1916
		x"22",	--1917
		x"62",	--1918
		x"3e",	--1919
		x"e2",	--1920
		x"1f",	--1921
		x"7c",	--1922
		x"b0",	--1923
		x"26",	--1924
		x"3e",	--1925
		x"e2",	--1926
		x"1f",	--1927
		x"7a",	--1928
		x"b0",	--1929
		x"26",	--1930
		x"30",	--1931
		x"2e",	--1932
		x"b0",	--1933
		x"94",	--1934
		x"21",	--1935
		x"1e",	--1936
		x"22",	--1937
		x"4e",	--1938
		x"82",	--1939
		x"7c",	--1940
		x"82",	--1941
		x"7a",	--1942
		x"30",	--1943
		x"82",	--1944
		x"7e",	--1945
		x"30",	--1946
		x"0b",	--1947
		x"0b",	--1948
		x"0e",	--1949
		x"3f",	--1950
		x"14",	--1951
		x"b0",	--1952
		x"5e",	--1953
		x"82",	--1954
		x"88",	--1955
		x"0d",	--1956
		x"0e",	--1957
		x"b0",	--1958
		x"a2",	--1959
		x"3b",	--1960
		x"30",	--1961
		x"1f",	--1962
		x"82",	--1963
		x"26",	--1964
		x"01",	--1965
		x"0f",	--1966
		x"82",	--1967
		x"26",	--1968
		x"0f",	--1969
		x"11",	--1970
		x"0e",	--1971
		x"1f",	--1972
		x"7c",	--1973
		x"b0",	--1974
		x"26",	--1975
		x"0e",	--1976
		x"1f",	--1977
		x"7a",	--1978
		x"b0",	--1979
		x"26",	--1980
		x"30",	--1981
		x"63",	--1982
		x"b0",	--1983
		x"94",	--1984
		x"21",	--1985
		x"0f",	--1986
		x"30",	--1987
		x"30",	--1988
		x"4f",	--1989
		x"b0",	--1990
		x"94",	--1991
		x"21",	--1992
		x"0f",	--1993
		x"30",	--1994
		x"8f",	--1995
		x"00",	--1996
		x"8f",	--1997
		x"02",	--1998
		x"9f",	--1999
		x"02",	--2000
		x"04",	--2001
		x"9f",	--2002
		x"04",	--2003
		x"06",	--2004
		x"9f",	--2005
		x"06",	--2006
		x"08",	--2007
		x"9f",	--2008
		x"08",	--2009
		x"0a",	--2010
		x"9f",	--2011
		x"0a",	--2012
		x"10",	--2013
		x"9f",	--2014
		x"0c",	--2015
		x"12",	--2016
		x"8f",	--2017
		x"14",	--2018
		x"8f",	--2019
		x"16",	--2020
		x"8f",	--2021
		x"0c",	--2022
		x"8f",	--2023
		x"0e",	--2024
		x"8f",	--2025
		x"18",	--2026
		x"8f",	--2027
		x"1a",	--2028
		x"8f",	--2029
		x"1c",	--2030
		x"8f",	--2031
		x"1e",	--2032
		x"30",	--2033
		x"8f",	--2034
		x"0c",	--2035
		x"8f",	--2036
		x"0e",	--2037
		x"8f",	--2038
		x"18",	--2039
		x"8f",	--2040
		x"1a",	--2041
		x"8f",	--2042
		x"1c",	--2043
		x"8f",	--2044
		x"1e",	--2045
		x"30",	--2046
		x"8f",	--2047
		x"00",	--2048
		x"8f",	--2049
		x"02",	--2050
		x"30",	--2051
		x"8f",	--2052
		x"04",	--2053
		x"8f",	--2054
		x"06",	--2055
		x"30",	--2056
		x"8f",	--2057
		x"08",	--2058
		x"8f",	--2059
		x"0a",	--2060
		x"30",	--2061
		x"8f",	--2062
		x"0c",	--2063
		x"8f",	--2064
		x"0e",	--2065
		x"30",	--2066
		x"8f",	--2067
		x"10",	--2068
		x"8f",	--2069
		x"12",	--2070
		x"30",	--2071
		x"0b",	--2072
		x"0a",	--2073
		x"09",	--2074
		x"07",	--2075
		x"06",	--2076
		x"05",	--2077
		x"04",	--2078
		x"09",	--2079
		x"04",	--2080
		x"05",	--2081
		x"16",	--2082
		x"14",	--2083
		x"17",	--2084
		x"16",	--2085
		x"1a",	--2086
		x"0c",	--2087
		x"1b",	--2088
		x"0e",	--2089
		x"0c",	--2090
		x"0d",	--2091
		x"0e",	--2092
		x"0f",	--2093
		x"b0",	--2094
		x"16",	--2095
		x"1c",	--2096
		x"10",	--2097
		x"1d",	--2098
		x"12",	--2099
		x"0f",	--2100
		x"5b",	--2101
		x"0e",	--2102
		x"0f",	--2103
		x"b0",	--2104
		x"16",	--2105
		x"06",	--2106
		x"07",	--2107
		x"89",	--2108
		x"14",	--2109
		x"89",	--2110
		x"16",	--2111
		x"0c",	--2112
		x"0d",	--2113
		x"0e",	--2114
		x"0f",	--2115
		x"b0",	--2116
		x"16",	--2117
		x"0f",	--2118
		x"5c",	--2119
		x"89",	--2120
		x"14",	--2121
		x"89",	--2122
		x"16",	--2123
		x"0c",	--2124
		x"0d",	--2125
		x"0e",	--2126
		x"0f",	--2127
		x"b0",	--2128
		x"62",	--2129
		x"0a",	--2130
		x"0b",	--2131
		x"1c",	--2132
		x"18",	--2133
		x"1d",	--2134
		x"1a",	--2135
		x"b0",	--2136
		x"16",	--2137
		x"06",	--2138
		x"07",	--2139
		x"89",	--2140
		x"18",	--2141
		x"89",	--2142
		x"1a",	--2143
		x"2c",	--2144
		x"1d",	--2145
		x"02",	--2146
		x"0e",	--2147
		x"0f",	--2148
		x"b0",	--2149
		x"b2",	--2150
		x"04",	--2151
		x"05",	--2152
		x"1c",	--2153
		x"04",	--2154
		x"1d",	--2155
		x"06",	--2156
		x"0e",	--2157
		x"0f",	--2158
		x"b0",	--2159
		x"b2",	--2160
		x"0c",	--2161
		x"0d",	--2162
		x"b0",	--2163
		x"16",	--2164
		x"06",	--2165
		x"07",	--2166
		x"1c",	--2167
		x"1c",	--2168
		x"1d",	--2169
		x"1e",	--2170
		x"0e",	--2171
		x"0f",	--2172
		x"b0",	--2173
		x"62",	--2174
		x"1c",	--2175
		x"08",	--2176
		x"1d",	--2177
		x"0a",	--2178
		x"b0",	--2179
		x"b2",	--2180
		x"0c",	--2181
		x"0d",	--2182
		x"b0",	--2183
		x"16",	--2184
		x"34",	--2185
		x"35",	--2186
		x"36",	--2187
		x"37",	--2188
		x"39",	--2189
		x"3a",	--2190
		x"3b",	--2191
		x"30",	--2192
		x"0e",	--2193
		x"0f",	--2194
		x"b0",	--2195
		x"62",	--2196
		x"06",	--2197
		x"07",	--2198
		x"89",	--2199
		x"14",	--2200
		x"89",	--2201
		x"16",	--2202
		x"0c",	--2203
		x"0d",	--2204
		x"0e",	--2205
		x"0f",	--2206
		x"b0",	--2207
		x"76",	--2208
		x"0f",	--2209
		x"01",	--2210
		x"a4",	--2211
		x"0a",	--2212
		x"0b",	--2213
		x"a5",	--2214
		x"0b",	--2215
		x"0a",	--2216
		x"21",	--2217
		x"0a",	--2218
		x"0b",	--2219
		x"30",	--2220
		x"79",	--2221
		x"b0",	--2222
		x"94",	--2223
		x"21",	--2224
		x"3a",	--2225
		x"03",	--2226
		x"1b",	--2227
		x"0e",	--2228
		x"1f",	--2229
		x"02",	--2230
		x"b0",	--2231
		x"b8",	--2232
		x"0a",	--2233
		x"0e",	--2234
		x"1f",	--2235
		x"04",	--2236
		x"b0",	--2237
		x"b8",	--2238
		x"0b",	--2239
		x"0f",	--2240
		x"0a",	--2241
		x"30",	--2242
		x"c1",	--2243
		x"b0",	--2244
		x"94",	--2245
		x"31",	--2246
		x"06",	--2247
		x"8a",	--2248
		x"00",	--2249
		x"0f",	--2250
		x"21",	--2251
		x"3a",	--2252
		x"3b",	--2253
		x"30",	--2254
		x"30",	--2255
		x"81",	--2256
		x"b0",	--2257
		x"94",	--2258
		x"b1",	--2259
		x"9b",	--2260
		x"00",	--2261
		x"b0",	--2262
		x"94",	--2263
		x"a1",	--2264
		x"00",	--2265
		x"30",	--2266
		x"ac",	--2267
		x"b0",	--2268
		x"94",	--2269
		x"21",	--2270
		x"3f",	--2271
		x"ea",	--2272
		x"0b",	--2273
		x"21",	--2274
		x"0b",	--2275
		x"1f",	--2276
		x"17",	--2277
		x"16",	--2278
		x"30",	--2279
		x"dc",	--2280
		x"b0",	--2281
		x"94",	--2282
		x"21",	--2283
		x"0e",	--2284
		x"1f",	--2285
		x"02",	--2286
		x"b0",	--2287
		x"b8",	--2288
		x"2f",	--2289
		x"0f",	--2290
		x"30",	--2291
		x"c1",	--2292
		x"b0",	--2293
		x"94",	--2294
		x"31",	--2295
		x"06",	--2296
		x"0f",	--2297
		x"21",	--2298
		x"3b",	--2299
		x"30",	--2300
		x"30",	--2301
		x"81",	--2302
		x"b0",	--2303
		x"94",	--2304
		x"b1",	--2305
		x"9b",	--2306
		x"00",	--2307
		x"b0",	--2308
		x"94",	--2309
		x"a1",	--2310
		x"00",	--2311
		x"30",	--2312
		x"cd",	--2313
		x"b0",	--2314
		x"94",	--2315
		x"21",	--2316
		x"3f",	--2317
		x"eb",	--2318
		x"0b",	--2319
		x"0a",	--2320
		x"09",	--2321
		x"08",	--2322
		x"07",	--2323
		x"06",	--2324
		x"06",	--2325
		x"07",	--2326
		x"08",	--2327
		x"09",	--2328
		x"b0",	--2329
		x"16",	--2330
		x"0a",	--2331
		x"0b",	--2332
		x"3c",	--2333
		x"db",	--2334
		x"3d",	--2335
		x"49",	--2336
		x"b0",	--2337
		x"66",	--2338
		x"0f",	--2339
		x"20",	--2340
		x"1f",	--2341
		x"3c",	--2342
		x"db",	--2343
		x"3d",	--2344
		x"49",	--2345
		x"0e",	--2346
		x"0f",	--2347
		x"b0",	--2348
		x"76",	--2349
		x"0f",	--2350
		x"01",	--2351
		x"09",	--2352
		x"0e",	--2353
		x"0f",	--2354
		x"36",	--2355
		x"37",	--2356
		x"38",	--2357
		x"39",	--2358
		x"3a",	--2359
		x"3b",	--2360
		x"30",	--2361
		x"3c",	--2362
		x"db",	--2363
		x"3d",	--2364
		x"c9",	--2365
		x"0e",	--2366
		x"0f",	--2367
		x"b0",	--2368
		x"62",	--2369
		x"0a",	--2370
		x"0b",	--2371
		x"ec",	--2372
		x"3c",	--2373
		x"db",	--2374
		x"3d",	--2375
		x"c9",	--2376
		x"0e",	--2377
		x"0f",	--2378
		x"b0",	--2379
		x"16",	--2380
		x"0c",	--2381
		x"0d",	--2382
		x"b0",	--2383
		x"16",	--2384
		x"0a",	--2385
		x"0b",	--2386
		x"dd",	--2387
		x"0b",	--2388
		x"0b",	--2389
		x"8f",	--2390
		x"0a",	--2391
		x"8f",	--2392
		x"0c",	--2393
		x"8f",	--2394
		x"0e",	--2395
		x"8f",	--2396
		x"10",	--2397
		x"8f",	--2398
		x"12",	--2399
		x"8f",	--2400
		x"14",	--2401
		x"8f",	--2402
		x"00",	--2403
		x"8f",	--2404
		x"02",	--2405
		x"9f",	--2406
		x"04",	--2407
		x"04",	--2408
		x"9f",	--2409
		x"06",	--2410
		x"06",	--2411
		x"9f",	--2412
		x"08",	--2413
		x"08",	--2414
		x"8f",	--2415
		x"16",	--2416
		x"8f",	--2417
		x"18",	--2418
		x"8f",	--2419
		x"1a",	--2420
		x"8f",	--2421
		x"1c",	--2422
		x"0e",	--2423
		x"3f",	--2424
		x"84",	--2425
		x"b0",	--2426
		x"5e",	--2427
		x"8b",	--2428
		x"22",	--2429
		x"3b",	--2430
		x"30",	--2431
		x"8f",	--2432
		x"20",	--2433
		x"8f",	--2434
		x"1e",	--2435
		x"30",	--2436
		x"0b",	--2437
		x"0a",	--2438
		x"09",	--2439
		x"08",	--2440
		x"07",	--2441
		x"05",	--2442
		x"04",	--2443
		x"31",	--2444
		x"f4",	--2445
		x"07",	--2446
		x"81",	--2447
		x"04",	--2448
		x"81",	--2449
		x"06",	--2450
		x"3c",	--2451
		x"db",	--2452
		x"3d",	--2453
		x"c9",	--2454
		x"2e",	--2455
		x"1f",	--2456
		x"02",	--2457
		x"b0",	--2458
		x"b2",	--2459
		x"0a",	--2460
		x"0b",	--2461
		x"1e",	--2462
		x"08",	--2463
		x"0f",	--2464
		x"8f",	--2465
		x"8f",	--2466
		x"8f",	--2467
		x"8f",	--2468
		x"b0",	--2469
		x"b6",	--2470
		x"0c",	--2471
		x"0d",	--2472
		x"0e",	--2473
		x"0f",	--2474
		x"b0",	--2475
		x"d6",	--2476
		x"0a",	--2477
		x"0b",	--2478
		x"18",	--2479
		x"04",	--2480
		x"19",	--2481
		x"06",	--2482
		x"18",	--2483
		x"16",	--2484
		x"19",	--2485
		x"18",	--2486
		x"14",	--2487
		x"1c",	--2488
		x"15",	--2489
		x"1e",	--2490
		x"14",	--2491
		x"1a",	--2492
		x"15",	--2493
		x"1c",	--2494
		x"0e",	--2495
		x"0f",	--2496
		x"b0",	--2497
		x"b6",	--2498
		x"0c",	--2499
		x"0d",	--2500
		x"b0",	--2501
		x"b2",	--2502
		x"81",	--2503
		x"00",	--2504
		x"81",	--2505
		x"02",	--2506
		x"0e",	--2507
		x"0f",	--2508
		x"b0",	--2509
		x"b6",	--2510
		x"0c",	--2511
		x"0d",	--2512
		x"b0",	--2513
		x"b2",	--2514
		x"0a",	--2515
		x"0b",	--2516
		x"0c",	--2517
		x"0d",	--2518
		x"2e",	--2519
		x"1f",	--2520
		x"02",	--2521
		x"b0",	--2522
		x"16",	--2523
		x"81",	--2524
		x"08",	--2525
		x"81",	--2526
		x"0a",	--2527
		x"08",	--2528
		x"a0",	--2529
		x"09",	--2530
		x"9e",	--2531
		x"04",	--2532
		x"02",	--2533
		x"30",	--2534
		x"7c",	--2535
		x"18",	--2536
		x"04",	--2537
		x"19",	--2538
		x"06",	--2539
		x"2c",	--2540
		x"1d",	--2541
		x"02",	--2542
		x"0e",	--2543
		x"0f",	--2544
		x"b0",	--2545
		x"62",	--2546
		x"0a",	--2547
		x"0b",	--2548
		x"0c",	--2549
		x"0d",	--2550
		x"1e",	--2551
		x"08",	--2552
		x"1f",	--2553
		x"0a",	--2554
		x"b0",	--2555
		x"b2",	--2556
		x"0c",	--2557
		x"0d",	--2558
		x"b0",	--2559
		x"d6",	--2560
		x"04",	--2561
		x"05",	--2562
		x"0c",	--2563
		x"0d",	--2564
		x"0e",	--2565
		x"0f",	--2566
		x"b0",	--2567
		x"16",	--2568
		x"0c",	--2569
		x"0d",	--2570
		x"0e",	--2571
		x"0f",	--2572
		x"b0",	--2573
		x"d6",	--2574
		x"b0",	--2575
		x"98",	--2576
		x"81",	--2577
		x"00",	--2578
		x"81",	--2579
		x"02",	--2580
		x"1a",	--2581
		x"12",	--2582
		x"1b",	--2583
		x"14",	--2584
		x"0e",	--2585
		x"0f",	--2586
		x"b0",	--2587
		x"3e",	--2588
		x"0c",	--2589
		x"0d",	--2590
		x"b0",	--2591
		x"b2",	--2592
		x"0c",	--2593
		x"0d",	--2594
		x"1e",	--2595
		x"0a",	--2596
		x"1f",	--2597
		x"0c",	--2598
		x"b0",	--2599
		x"62",	--2600
		x"81",	--2601
		x"08",	--2602
		x"81",	--2603
		x"0a",	--2604
		x"0e",	--2605
		x"0f",	--2606
		x"b0",	--2607
		x"18",	--2608
		x"0c",	--2609
		x"0d",	--2610
		x"b0",	--2611
		x"b2",	--2612
		x"1c",	--2613
		x"0e",	--2614
		x"1d",	--2615
		x"10",	--2616
		x"b0",	--2617
		x"16",	--2618
		x"08",	--2619
		x"09",	--2620
		x"2c",	--2621
		x"1d",	--2622
		x"02",	--2623
		x"0e",	--2624
		x"0f",	--2625
		x"b0",	--2626
		x"1e",	--2627
		x"0a",	--2628
		x"0b",	--2629
		x"87",	--2630
		x"12",	--2631
		x"87",	--2632
		x"14",	--2633
		x"b0",	--2634
		x"3e",	--2635
		x"0c",	--2636
		x"0d",	--2637
		x"b0",	--2638
		x"b2",	--2639
		x"1c",	--2640
		x"08",	--2641
		x"1d",	--2642
		x"0a",	--2643
		x"b0",	--2644
		x"16",	--2645
		x"87",	--2646
		x"0a",	--2647
		x"87",	--2648
		x"0c",	--2649
		x"0e",	--2650
		x"0f",	--2651
		x"b0",	--2652
		x"18",	--2653
		x"0c",	--2654
		x"0d",	--2655
		x"b0",	--2656
		x"b2",	--2657
		x"0c",	--2658
		x"0d",	--2659
		x"0e",	--2660
		x"0f",	--2661
		x"b0",	--2662
		x"62",	--2663
		x"87",	--2664
		x"0e",	--2665
		x"87",	--2666
		x"10",	--2667
		x"97",	--2668
		x"04",	--2669
		x"16",	--2670
		x"97",	--2671
		x"06",	--2672
		x"18",	--2673
		x"97",	--2674
		x"1c",	--2675
		x"1a",	--2676
		x"97",	--2677
		x"1e",	--2678
		x"1c",	--2679
		x"31",	--2680
		x"0c",	--2681
		x"34",	--2682
		x"35",	--2683
		x"37",	--2684
		x"38",	--2685
		x"39",	--2686
		x"3a",	--2687
		x"3b",	--2688
		x"30",	--2689
		x"08",	--2690
		x"64",	--2691
		x"09",	--2692
		x"62",	--2693
		x"0c",	--2694
		x"3d",	--2695
		x"00",	--2696
		x"1e",	--2697
		x"08",	--2698
		x"1f",	--2699
		x"0a",	--2700
		x"b0",	--2701
		x"b2",	--2702
		x"0a",	--2703
		x"0b",	--2704
		x"18",	--2705
		x"12",	--2706
		x"19",	--2707
		x"14",	--2708
		x"0e",	--2709
		x"0f",	--2710
		x"b0",	--2711
		x"18",	--2712
		x"0c",	--2713
		x"0d",	--2714
		x"b0",	--2715
		x"b2",	--2716
		x"0c",	--2717
		x"0d",	--2718
		x"1e",	--2719
		x"0a",	--2720
		x"1f",	--2721
		x"0c",	--2722
		x"b0",	--2723
		x"16",	--2724
		x"87",	--2725
		x"0a",	--2726
		x"87",	--2727
		x"0c",	--2728
		x"0e",	--2729
		x"0f",	--2730
		x"b0",	--2731
		x"3e",	--2732
		x"0c",	--2733
		x"0d",	--2734
		x"b0",	--2735
		x"b2",	--2736
		x"0c",	--2737
		x"0d",	--2738
		x"1e",	--2739
		x"0e",	--2740
		x"1f",	--2741
		x"10",	--2742
		x"b0",	--2743
		x"16",	--2744
		x"87",	--2745
		x"0e",	--2746
		x"87",	--2747
		x"10",	--2748
		x"ae",	--2749
		x"05",	--2750
		x"ac",	--2751
		x"30",	--2752
		x"d0",	--2753
		x"0b",	--2754
		x"0a",	--2755
		x"09",	--2756
		x"09",	--2757
		x"1f",	--2758
		x"20",	--2759
		x"b0",	--2760
		x"7e",	--2761
		x"0a",	--2762
		x"0b",	--2763
		x"1f",	--2764
		x"1e",	--2765
		x"b0",	--2766
		x"7e",	--2767
		x"0c",	--2768
		x"0d",	--2769
		x"3c",	--2770
		x"3d",	--2771
		x"1c",	--2772
		x"0d",	--2773
		x"0d",	--2774
		x"0c",	--2775
		x"0d",	--2776
		x"0e",	--2777
		x"0f",	--2778
		x"b0",	--2779
		x"0a",	--2780
		x"21",	--2781
		x"39",	--2782
		x"3a",	--2783
		x"3b",	--2784
		x"30",	--2785
		x"0d",	--2786
		x"1f",	--2787
		x"22",	--2788
		x"b0",	--2789
		x"a2",	--2790
		x"30",	--2791
		x"1f",	--2792
		x"22",	--2793
		x"b0",	--2794
		x"ca",	--2795
		x"30",	--2796
		x"0b",	--2797
		x"0a",	--2798
		x"0b",	--2799
		x"0a",	--2800
		x"8f",	--2801
		x"00",	--2802
		x"8f",	--2803
		x"02",	--2804
		x"8f",	--2805
		x"04",	--2806
		x"0c",	--2807
		x"0d",	--2808
		x"3e",	--2809
		x"00",	--2810
		x"3f",	--2811
		x"6e",	--2812
		x"b0",	--2813
		x"52",	--2814
		x"8b",	--2815
		x"02",	--2816
		x"02",	--2817
		x"32",	--2818
		x"03",	--2819
		x"82",	--2820
		x"32",	--2821
		x"b2",	--2822
		x"18",	--2823
		x"38",	--2824
		x"9b",	--2825
		x"3a",	--2826
		x"06",	--2827
		x"32",	--2828
		x"0f",	--2829
		x"3a",	--2830
		x"3b",	--2831
		x"30",	--2832
		x"0b",	--2833
		x"09",	--2834
		x"08",	--2835
		x"8f",	--2836
		x"06",	--2837
		x"bf",	--2838
		x"00",	--2839
		x"08",	--2840
		x"2b",	--2841
		x"1e",	--2842
		x"02",	--2843
		x"0f",	--2844
		x"b0",	--2845
		x"ec",	--2846
		x"0c",	--2847
		x"3d",	--2848
		x"00",	--2849
		x"b0",	--2850
		x"b2",	--2851
		x"08",	--2852
		x"09",	--2853
		x"1e",	--2854
		x"06",	--2855
		x"0f",	--2856
		x"b0",	--2857
		x"ec",	--2858
		x"0c",	--2859
		x"0d",	--2860
		x"0e",	--2861
		x"0f",	--2862
		x"b0",	--2863
		x"62",	--2864
		x"b0",	--2865
		x"42",	--2866
		x"8b",	--2867
		x"04",	--2868
		x"9b",	--2869
		x"00",	--2870
		x"38",	--2871
		x"39",	--2872
		x"3b",	--2873
		x"30",	--2874
		x"0b",	--2875
		x"0a",	--2876
		x"09",	--2877
		x"0a",	--2878
		x"0b",	--2879
		x"8f",	--2880
		x"06",	--2881
		x"8f",	--2882
		x"08",	--2883
		x"29",	--2884
		x"1e",	--2885
		x"02",	--2886
		x"0f",	--2887
		x"b0",	--2888
		x"ec",	--2889
		x"0c",	--2890
		x"0d",	--2891
		x"0e",	--2892
		x"0f",	--2893
		x"b0",	--2894
		x"b2",	--2895
		x"0a",	--2896
		x"0b",	--2897
		x"1e",	--2898
		x"06",	--2899
		x"0f",	--2900
		x"b0",	--2901
		x"ec",	--2902
		x"0c",	--2903
		x"0d",	--2904
		x"0e",	--2905
		x"0f",	--2906
		x"b0",	--2907
		x"62",	--2908
		x"b0",	--2909
		x"42",	--2910
		x"89",	--2911
		x"04",	--2912
		x"39",	--2913
		x"3a",	--2914
		x"3b",	--2915
		x"30",	--2916
		x"2f",	--2917
		x"8f",	--2918
		x"04",	--2919
		x"30",	--2920
		x"0b",	--2921
		x"0a",	--2922
		x"92",	--2923
		x"2a",	--2924
		x"14",	--2925
		x"3b",	--2926
		x"8e",	--2927
		x"0a",	--2928
		x"2b",	--2929
		x"5f",	--2930
		x"fc",	--2931
		x"8f",	--2932
		x"0f",	--2933
		x"30",	--2934
		x"e3",	--2935
		x"b0",	--2936
		x"94",	--2937
		x"31",	--2938
		x"06",	--2939
		x"1a",	--2940
		x"3b",	--2941
		x"06",	--2942
		x"1a",	--2943
		x"2a",	--2944
		x"ef",	--2945
		x"0f",	--2946
		x"3a",	--2947
		x"3b",	--2948
		x"30",	--2949
		x"1e",	--2950
		x"2a",	--2951
		x"3e",	--2952
		x"20",	--2953
		x"12",	--2954
		x"0f",	--2955
		x"0f",	--2956
		x"0f",	--2957
		x"0f",	--2958
		x"3f",	--2959
		x"8a",	--2960
		x"ff",	--2961
		x"68",	--2962
		x"00",	--2963
		x"bf",	--2964
		x"d2",	--2965
		x"02",	--2966
		x"bf",	--2967
		x"12",	--2968
		x"04",	--2969
		x"1e",	--2970
		x"82",	--2971
		x"2a",	--2972
		x"30",	--2973
		x"0b",	--2974
		x"1b",	--2975
		x"2a",	--2976
		x"3b",	--2977
		x"20",	--2978
		x"12",	--2979
		x"0c",	--2980
		x"0c",	--2981
		x"0c",	--2982
		x"0c",	--2983
		x"3c",	--2984
		x"8a",	--2985
		x"cc",	--2986
		x"00",	--2987
		x"8c",	--2988
		x"02",	--2989
		x"8c",	--2990
		x"04",	--2991
		x"1b",	--2992
		x"82",	--2993
		x"2a",	--2994
		x"0f",	--2995
		x"3b",	--2996
		x"30",	--2997
		x"3f",	--2998
		x"fc",	--2999
		x"0b",	--3000
		x"31",	--3001
		x"f0",	--3002
		x"1b",	--3003
		x"2a",	--3004
		x"1b",	--3005
		x"0f",	--3006
		x"5f",	--3007
		x"8a",	--3008
		x"16",	--3009
		x"3d",	--3010
		x"90",	--3011
		x"0c",	--3012
		x"05",	--3013
		x"3d",	--3014
		x"06",	--3015
		x"cd",	--3016
		x"fa",	--3017
		x"0e",	--3018
		x"1c",	--3019
		x"0c",	--3020
		x"f8",	--3021
		x"30",	--3022
		x"eb",	--3023
		x"b0",	--3024
		x"94",	--3025
		x"21",	--3026
		x"3f",	--3027
		x"31",	--3028
		x"10",	--3029
		x"3b",	--3030
		x"30",	--3031
		x"0c",	--3032
		x"81",	--3033
		x"00",	--3034
		x"6d",	--3035
		x"4d",	--3036
		x"24",	--3037
		x"1e",	--3038
		x"1f",	--3039
		x"06",	--3040
		x"6d",	--3041
		x"4d",	--3042
		x"11",	--3043
		x"1e",	--3044
		x"3f",	--3045
		x"0e",	--3046
		x"7d",	--3047
		x"20",	--3048
		x"f7",	--3049
		x"ce",	--3050
		x"ff",	--3051
		x"0d",	--3052
		x"0d",	--3053
		x"0d",	--3054
		x"8d",	--3055
		x"00",	--3056
		x"1f",	--3057
		x"6d",	--3058
		x"4d",	--3059
		x"ef",	--3060
		x"0e",	--3061
		x"0e",	--3062
		x"0c",	--3063
		x"0c",	--3064
		x"3c",	--3065
		x"8a",	--3066
		x"0e",	--3067
		x"9c",	--3068
		x"02",	--3069
		x"31",	--3070
		x"10",	--3071
		x"3b",	--3072
		x"30",	--3073
		x"1f",	--3074
		x"f1",	--3075
		x"8f",	--3076
		x"00",	--3077
		x"0f",	--3078
		x"30",	--3079
		x"0e",	--3080
		x"2e",	--3081
		x"2f",	--3082
		x"30",	--3083
		x"0b",	--3084
		x"0a",	--3085
		x"0e",	--3086
		x"2e",	--3087
		x"2c",	--3088
		x"0d",	--3089
		x"0e",	--3090
		x"0f",	--3091
		x"0e",	--3092
		x"0f",	--3093
		x"0a",	--3094
		x"0b",	--3095
		x"0a",	--3096
		x"0b",	--3097
		x"0a",	--3098
		x"0b",	--3099
		x"3c",	--3100
		x"3a",	--3101
		x"0d",	--3102
		x"0e",	--3103
		x"0f",	--3104
		x"b0",	--3105
		x"12",	--3106
		x"0f",	--3107
		x"3a",	--3108
		x"3b",	--3109
		x"30",	--3110
		x"b2",	--3111
		x"d2",	--3112
		x"60",	--3113
		x"b2",	--3114
		x"b8",	--3115
		x"72",	--3116
		x"0f",	--3117
		x"30",	--3118
		x"0b",	--3119
		x"0b",	--3120
		x"1f",	--3121
		x"2c",	--3122
		x"3f",	--3123
		x"20",	--3124
		x"19",	--3125
		x"0c",	--3126
		x"0c",	--3127
		x"0d",	--3128
		x"0d",	--3129
		x"0d",	--3130
		x"0d",	--3131
		x"0d",	--3132
		x"3d",	--3133
		x"4a",	--3134
		x"8d",	--3135
		x"00",	--3136
		x"8d",	--3137
		x"02",	--3138
		x"8d",	--3139
		x"08",	--3140
		x"8d",	--3141
		x"0a",	--3142
		x"8d",	--3143
		x"0c",	--3144
		x"0e",	--3145
		x"1e",	--3146
		x"82",	--3147
		x"2c",	--3148
		x"3b",	--3149
		x"30",	--3150
		x"3f",	--3151
		x"fc",	--3152
		x"0f",	--3153
		x"0c",	--3154
		x"0c",	--3155
		x"0c",	--3156
		x"0c",	--3157
		x"0c",	--3158
		x"3c",	--3159
		x"4a",	--3160
		x"8c",	--3161
		x"02",	--3162
		x"8c",	--3163
		x"04",	--3164
		x"8c",	--3165
		x"06",	--3166
		x"8c",	--3167
		x"08",	--3168
		x"9c",	--3169
		x"00",	--3170
		x"0f",	--3171
		x"30",	--3172
		x"0f",	--3173
		x"0e",	--3174
		x"0e",	--3175
		x"0e",	--3176
		x"0e",	--3177
		x"0e",	--3178
		x"8e",	--3179
		x"4a",	--3180
		x"0f",	--3181
		x"30",	--3182
		x"0f",	--3183
		x"0e",	--3184
		x"0d",	--3185
		x"0c",	--3186
		x"0b",	--3187
		x"0a",	--3188
		x"09",	--3189
		x"08",	--3190
		x"07",	--3191
		x"92",	--3192
		x"2c",	--3193
		x"33",	--3194
		x"3a",	--3195
		x"4a",	--3196
		x"0b",	--3197
		x"2b",	--3198
		x"08",	--3199
		x"38",	--3200
		x"07",	--3201
		x"37",	--3202
		x"06",	--3203
		x"09",	--3204
		x"0f",	--3205
		x"1f",	--3206
		x"8b",	--3207
		x"00",	--3208
		x"19",	--3209
		x"3a",	--3210
		x"0e",	--3211
		x"3b",	--3212
		x"0e",	--3213
		x"38",	--3214
		x"0e",	--3215
		x"37",	--3216
		x"0e",	--3217
		x"19",	--3218
		x"2c",	--3219
		x"19",	--3220
		x"8a",	--3221
		x"00",	--3222
		x"f1",	--3223
		x"2f",	--3224
		x"1f",	--3225
		x"02",	--3226
		x"ea",	--3227
		x"8b",	--3228
		x"00",	--3229
		x"1f",	--3230
		x"0a",	--3231
		x"9b",	--3232
		x"08",	--3233
		x"88",	--3234
		x"00",	--3235
		x"e4",	--3236
		x"2f",	--3237
		x"1f",	--3238
		x"87",	--3239
		x"00",	--3240
		x"2f",	--3241
		x"de",	--3242
		x"8a",	--3243
		x"00",	--3244
		x"db",	--3245
		x"b2",	--3246
		x"fe",	--3247
		x"60",	--3248
		x"37",	--3249
		x"38",	--3250
		x"39",	--3251
		x"3a",	--3252
		x"3b",	--3253
		x"3c",	--3254
		x"3d",	--3255
		x"3e",	--3256
		x"3f",	--3257
		x"00",	--3258
		x"8f",	--3259
		x"00",	--3260
		x"0f",	--3261
		x"30",	--3262
		x"2f",	--3263
		x"2e",	--3264
		x"1f",	--3265
		x"02",	--3266
		x"30",	--3267
		x"8f",	--3268
		x"00",	--3269
		x"30",	--3270
		x"8f",	--3271
		x"00",	--3272
		x"3f",	--3273
		x"88",	--3274
		x"b0",	--3275
		x"5e",	--3276
		x"82",	--3277
		x"18",	--3278
		x"0f",	--3279
		x"30",	--3280
		x"0c",	--3281
		x"2f",	--3282
		x"8f",	--3283
		x"00",	--3284
		x"1d",	--3285
		x"0e",	--3286
		x"1f",	--3287
		x"18",	--3288
		x"b0",	--3289
		x"a2",	--3290
		x"30",	--3291
		x"5e",	--3292
		x"81",	--3293
		x"3e",	--3294
		x"fc",	--3295
		x"c2",	--3296
		x"84",	--3297
		x"0f",	--3298
		x"30",	--3299
		x"3f",	--3300
		x"0f",	--3301
		x"5f",	--3302
		x"aa",	--3303
		x"8f",	--3304
		x"b0",	--3305
		x"b8",	--3306
		x"30",	--3307
		x"0b",	--3308
		x"0b",	--3309
		x"0e",	--3310
		x"0e",	--3311
		x"0e",	--3312
		x"0e",	--3313
		x"0e",	--3314
		x"0f",	--3315
		x"b0",	--3316
		x"c8",	--3317
		x"0f",	--3318
		x"b0",	--3319
		x"c8",	--3320
		x"3b",	--3321
		x"30",	--3322
		x"0b",	--3323
		x"0a",	--3324
		x"0a",	--3325
		x"3b",	--3326
		x"07",	--3327
		x"0e",	--3328
		x"4d",	--3329
		x"7d",	--3330
		x"0f",	--3331
		x"03",	--3332
		x"0e",	--3333
		x"7d",	--3334
		x"fd",	--3335
		x"1e",	--3336
		x"0a",	--3337
		x"3f",	--3338
		x"31",	--3339
		x"b0",	--3340
		x"b8",	--3341
		x"3b",	--3342
		x"3b",	--3343
		x"ef",	--3344
		x"3a",	--3345
		x"3b",	--3346
		x"30",	--3347
		x"3f",	--3348
		x"30",	--3349
		x"f5",	--3350
		x"0b",	--3351
		x"0b",	--3352
		x"0e",	--3353
		x"8e",	--3354
		x"8e",	--3355
		x"0f",	--3356
		x"b0",	--3357
		x"d8",	--3358
		x"0f",	--3359
		x"b0",	--3360
		x"d8",	--3361
		x"3b",	--3362
		x"30",	--3363
		x"0b",	--3364
		x"0a",	--3365
		x"0a",	--3366
		x"0b",	--3367
		x"0d",	--3368
		x"8d",	--3369
		x"8d",	--3370
		x"0f",	--3371
		x"b0",	--3372
		x"d8",	--3373
		x"0f",	--3374
		x"b0",	--3375
		x"d8",	--3376
		x"0c",	--3377
		x"0d",	--3378
		x"8d",	--3379
		x"8c",	--3380
		x"4d",	--3381
		x"0d",	--3382
		x"0f",	--3383
		x"b0",	--3384
		x"d8",	--3385
		x"0f",	--3386
		x"b0",	--3387
		x"d8",	--3388
		x"3a",	--3389
		x"3b",	--3390
		x"30",	--3391
		x"0b",	--3392
		x"0a",	--3393
		x"09",	--3394
		x"0a",	--3395
		x"0e",	--3396
		x"19",	--3397
		x"09",	--3398
		x"39",	--3399
		x"0b",	--3400
		x"0d",	--3401
		x"0d",	--3402
		x"6f",	--3403
		x"8f",	--3404
		x"b0",	--3405
		x"d8",	--3406
		x"0b",	--3407
		x"0e",	--3408
		x"1b",	--3409
		x"3b",	--3410
		x"07",	--3411
		x"05",	--3412
		x"3f",	--3413
		x"20",	--3414
		x"b0",	--3415
		x"b8",	--3416
		x"ef",	--3417
		x"3f",	--3418
		x"3a",	--3419
		x"b0",	--3420
		x"b8",	--3421
		x"ea",	--3422
		x"39",	--3423
		x"3a",	--3424
		x"3b",	--3425
		x"30",	--3426
		x"0b",	--3427
		x"0a",	--3428
		x"09",	--3429
		x"0a",	--3430
		x"0e",	--3431
		x"17",	--3432
		x"09",	--3433
		x"39",	--3434
		x"0b",	--3435
		x"6f",	--3436
		x"8f",	--3437
		x"b0",	--3438
		x"c8",	--3439
		x"0b",	--3440
		x"0e",	--3441
		x"1b",	--3442
		x"3b",	--3443
		x"07",	--3444
		x"f6",	--3445
		x"3f",	--3446
		x"20",	--3447
		x"b0",	--3448
		x"b8",	--3449
		x"6f",	--3450
		x"8f",	--3451
		x"b0",	--3452
		x"c8",	--3453
		x"0b",	--3454
		x"f2",	--3455
		x"39",	--3456
		x"3a",	--3457
		x"3b",	--3458
		x"30",	--3459
		x"0b",	--3460
		x"0a",	--3461
		x"09",	--3462
		x"31",	--3463
		x"ec",	--3464
		x"0b",	--3465
		x"0f",	--3466
		x"34",	--3467
		x"3b",	--3468
		x"0a",	--3469
		x"38",	--3470
		x"09",	--3471
		x"0a",	--3472
		x"0a",	--3473
		x"3e",	--3474
		x"0a",	--3475
		x"0f",	--3476
		x"b0",	--3477
		x"0a",	--3478
		x"7f",	--3479
		x"30",	--3480
		x"ca",	--3481
		x"00",	--3482
		x"19",	--3483
		x"3e",	--3484
		x"0a",	--3485
		x"0f",	--3486
		x"b0",	--3487
		x"d8",	--3488
		x"0b",	--3489
		x"3f",	--3490
		x"0a",	--3491
		x"eb",	--3492
		x"0a",	--3493
		x"1a",	--3494
		x"09",	--3495
		x"3e",	--3496
		x"0a",	--3497
		x"0f",	--3498
		x"b0",	--3499
		x"0a",	--3500
		x"7f",	--3501
		x"30",	--3502
		x"c9",	--3503
		x"00",	--3504
		x"3a",	--3505
		x"0f",	--3506
		x"0f",	--3507
		x"6f",	--3508
		x"8f",	--3509
		x"b0",	--3510
		x"b8",	--3511
		x"0a",	--3512
		x"f7",	--3513
		x"31",	--3514
		x"14",	--3515
		x"39",	--3516
		x"3a",	--3517
		x"3b",	--3518
		x"30",	--3519
		x"3f",	--3520
		x"2d",	--3521
		x"b0",	--3522
		x"b8",	--3523
		x"3b",	--3524
		x"1b",	--3525
		x"c5",	--3526
		x"1a",	--3527
		x"09",	--3528
		x"dd",	--3529
		x"0b",	--3530
		x"0a",	--3531
		x"09",	--3532
		x"0b",	--3533
		x"3b",	--3534
		x"39",	--3535
		x"6f",	--3536
		x"4f",	--3537
		x"0b",	--3538
		x"1a",	--3539
		x"8f",	--3540
		x"b0",	--3541
		x"b8",	--3542
		x"0a",	--3543
		x"09",	--3544
		x"19",	--3545
		x"5f",	--3546
		x"01",	--3547
		x"4f",	--3548
		x"10",	--3549
		x"7f",	--3550
		x"25",	--3551
		x"f3",	--3552
		x"0a",	--3553
		x"1a",	--3554
		x"5f",	--3555
		x"01",	--3556
		x"7f",	--3557
		x"db",	--3558
		x"7f",	--3559
		x"54",	--3560
		x"ee",	--3561
		x"4f",	--3562
		x"0f",	--3563
		x"10",	--3564
		x"02",	--3565
		x"39",	--3566
		x"3a",	--3567
		x"3b",	--3568
		x"30",	--3569
		x"09",	--3570
		x"29",	--3571
		x"1e",	--3572
		x"02",	--3573
		x"2f",	--3574
		x"b0",	--3575
		x"80",	--3576
		x"0b",	--3577
		x"dd",	--3578
		x"09",	--3579
		x"29",	--3580
		x"2f",	--3581
		x"b0",	--3582
		x"2e",	--3583
		x"0b",	--3584
		x"d6",	--3585
		x"0f",	--3586
		x"2b",	--3587
		x"29",	--3588
		x"6f",	--3589
		x"4f",	--3590
		x"d0",	--3591
		x"19",	--3592
		x"8f",	--3593
		x"b0",	--3594
		x"b8",	--3595
		x"7f",	--3596
		x"4f",	--3597
		x"fa",	--3598
		x"c8",	--3599
		x"09",	--3600
		x"29",	--3601
		x"1e",	--3602
		x"02",	--3603
		x"2f",	--3604
		x"b0",	--3605
		x"c6",	--3606
		x"0b",	--3607
		x"bf",	--3608
		x"09",	--3609
		x"29",	--3610
		x"2e",	--3611
		x"0f",	--3612
		x"8f",	--3613
		x"8f",	--3614
		x"8f",	--3615
		x"8f",	--3616
		x"b0",	--3617
		x"48",	--3618
		x"0b",	--3619
		x"b3",	--3620
		x"09",	--3621
		x"29",	--3622
		x"2f",	--3623
		x"b0",	--3624
		x"08",	--3625
		x"0b",	--3626
		x"ac",	--3627
		x"09",	--3628
		x"29",	--3629
		x"2f",	--3630
		x"b0",	--3631
		x"b8",	--3632
		x"0b",	--3633
		x"a5",	--3634
		x"09",	--3635
		x"29",	--3636
		x"2f",	--3637
		x"b0",	--3638
		x"d8",	--3639
		x"0b",	--3640
		x"9e",	--3641
		x"09",	--3642
		x"29",	--3643
		x"2f",	--3644
		x"b0",	--3645
		x"f6",	--3646
		x"0b",	--3647
		x"97",	--3648
		x"3f",	--3649
		x"25",	--3650
		x"b0",	--3651
		x"b8",	--3652
		x"92",	--3653
		x"0f",	--3654
		x"0e",	--3655
		x"1f",	--3656
		x"2e",	--3657
		x"df",	--3658
		x"85",	--3659
		x"0a",	--3660
		x"1f",	--3661
		x"2e",	--3662
		x"3f",	--3663
		x"3f",	--3664
		x"13",	--3665
		x"92",	--3666
		x"2e",	--3667
		x"1e",	--3668
		x"2e",	--3669
		x"1f",	--3670
		x"30",	--3671
		x"0e",	--3672
		x"02",	--3673
		x"92",	--3674
		x"30",	--3675
		x"f2",	--3676
		x"10",	--3677
		x"81",	--3678
		x"3e",	--3679
		x"3f",	--3680
		x"b1",	--3681
		x"f0",	--3682
		x"00",	--3683
		x"00",	--3684
		x"82",	--3685
		x"2e",	--3686
		x"ec",	--3687
		x"0c",	--3688
		x"0d",	--3689
		x"3e",	--3690
		x"00",	--3691
		x"3f",	--3692
		x"6e",	--3693
		x"b0",	--3694
		x"12",	--3695
		x"3e",	--3696
		x"82",	--3697
		x"82",	--3698
		x"f2",	--3699
		x"11",	--3700
		x"80",	--3701
		x"30",	--3702
		x"1e",	--3703
		x"2e",	--3704
		x"1f",	--3705
		x"30",	--3706
		x"0e",	--3707
		x"05",	--3708
		x"1f",	--3709
		x"2e",	--3710
		x"1f",	--3711
		x"30",	--3712
		x"30",	--3713
		x"1d",	--3714
		x"2e",	--3715
		x"1e",	--3716
		x"30",	--3717
		x"3f",	--3718
		x"40",	--3719
		x"0f",	--3720
		x"0f",	--3721
		x"30",	--3722
		x"1f",	--3723
		x"30",	--3724
		x"5f",	--3725
		x"0a",	--3726
		x"1d",	--3727
		x"30",	--3728
		x"1e",	--3729
		x"2e",	--3730
		x"0d",	--3731
		x"0b",	--3732
		x"1e",	--3733
		x"30",	--3734
		x"3e",	--3735
		x"3f",	--3736
		x"03",	--3737
		x"82",	--3738
		x"30",	--3739
		x"30",	--3740
		x"92",	--3741
		x"30",	--3742
		x"30",	--3743
		x"4f",	--3744
		x"30",	--3745
		x"0b",	--3746
		x"0a",	--3747
		x"09",	--3748
		x"08",	--3749
		x"07",	--3750
		x"06",	--3751
		x"05",	--3752
		x"04",	--3753
		x"31",	--3754
		x"04",	--3755
		x"05",	--3756
		x"81",	--3757
		x"00",	--3758
		x"81",	--3759
		x"02",	--3760
		x"08",	--3761
		x"09",	--3762
		x"38",	--3763
		x"39",	--3764
		x"ff",	--3765
		x"39",	--3766
		x"80",	--3767
		x"1f",	--3768
		x"39",	--3769
		x"80",	--3770
		x"0b",	--3771
		x"02",	--3772
		x"18",	--3773
		x"08",	--3774
		x"0c",	--3775
		x"0d",	--3776
		x"0e",	--3777
		x"0f",	--3778
		x"b0",	--3779
		x"16",	--3780
		x"30",	--3781
		x"18",	--3782
		x"81",	--3783
		x"02",	--3784
		x"02",	--3785
		x"30",	--3786
		x"78",	--3787
		x"05",	--3788
		x"91",	--3789
		x"00",	--3790
		x"02",	--3791
		x"30",	--3792
		x"78",	--3793
		x"34",	--3794
		x"db",	--3795
		x"35",	--3796
		x"c9",	--3797
		x"30",	--3798
		x"80",	--3799
		x"39",	--3800
		x"e0",	--3801
		x"08",	--3802
		x"0a",	--3803
		x"0b",	--3804
		x"3b",	--3805
		x"ff",	--3806
		x"39",	--3807
		x"98",	--3808
		x"1b",	--3809
		x"16",	--3810
		x"39",	--3811
		x"00",	--3812
		x"10",	--3813
		x"3c",	--3814
		x"ca",	--3815
		x"3d",	--3816
		x"49",	--3817
		x"b0",	--3818
		x"16",	--3819
		x"0c",	--3820
		x"3d",	--3821
		x"80",	--3822
		x"b0",	--3823
		x"76",	--3824
		x"0f",	--3825
		x"03",	--3826
		x"02",	--3827
		x"30",	--3828
		x"80",	--3829
		x"36",	--3830
		x"37",	--3831
		x"6d",	--3832
		x"39",	--3833
		x"1c",	--3834
		x"4b",	--3835
		x"3d",	--3836
		x"39",	--3837
		x"30",	--3838
		x"1b",	--3839
		x"0c",	--3840
		x"3d",	--3841
		x"80",	--3842
		x"0e",	--3843
		x"0f",	--3844
		x"b0",	--3845
		x"62",	--3846
		x"08",	--3847
		x"09",	--3848
		x"0c",	--3849
		x"3d",	--3850
		x"80",	--3851
		x"0e",	--3852
		x"0f",	--3853
		x"b0",	--3854
		x"16",	--3855
		x"0c",	--3856
		x"0d",	--3857
		x"0e",	--3858
		x"0f",	--3859
		x"b0",	--3860
		x"d6",	--3861
		x"04",	--3862
		x"05",	--3863
		x"16",	--3864
		x"07",	--3865
		x"4b",	--3866
		x"0c",	--3867
		x"0d",	--3868
		x"0e",	--3869
		x"0f",	--3870
		x"b0",	--3871
		x"16",	--3872
		x"0c",	--3873
		x"3d",	--3874
		x"80",	--3875
		x"b0",	--3876
		x"62",	--3877
		x"08",	--3878
		x"09",	--3879
		x"0c",	--3880
		x"3d",	--3881
		x"00",	--3882
		x"0e",	--3883
		x"0f",	--3884
		x"b0",	--3885
		x"16",	--3886
		x"0c",	--3887
		x"0d",	--3888
		x"0e",	--3889
		x"0f",	--3890
		x"b0",	--3891
		x"d6",	--3892
		x"04",	--3893
		x"05",	--3894
		x"06",	--3895
		x"07",	--3896
		x"2c",	--3897
		x"0c",	--3898
		x"0d",	--3899
		x"0e",	--3900
		x"3f",	--3901
		x"80",	--3902
		x"b0",	--3903
		x"d6",	--3904
		x"04",	--3905
		x"05",	--3906
		x"36",	--3907
		x"03",	--3908
		x"07",	--3909
		x"1f",	--3910
		x"0c",	--3911
		x"3d",	--3912
		x"c0",	--3913
		x"0e",	--3914
		x"0f",	--3915
		x"b0",	--3916
		x"62",	--3917
		x"08",	--3918
		x"09",	--3919
		x"0c",	--3920
		x"3d",	--3921
		x"c0",	--3922
		x"0e",	--3923
		x"0f",	--3924
		x"b0",	--3925
		x"b2",	--3926
		x"0c",	--3927
		x"3d",	--3928
		x"80",	--3929
		x"b0",	--3930
		x"16",	--3931
		x"0c",	--3932
		x"0d",	--3933
		x"0e",	--3934
		x"0f",	--3935
		x"b0",	--3936
		x"d6",	--3937
		x"04",	--3938
		x"05",	--3939
		x"26",	--3940
		x"07",	--3941
		x"0c",	--3942
		x"0d",	--3943
		x"0e",	--3944
		x"0f",	--3945
		x"b0",	--3946
		x"b2",	--3947
		x"08",	--3948
		x"09",	--3949
		x"0c",	--3950
		x"0d",	--3951
		x"b0",	--3952
		x"b2",	--3953
		x"0a",	--3954
		x"0b",	--3955
		x"3c",	--3956
		x"d7",	--3957
		x"3d",	--3958
		x"85",	--3959
		x"b0",	--3960
		x"b2",	--3961
		x"3c",	--3962
		x"59",	--3963
		x"3d",	--3964
		x"4b",	--3965
		x"b0",	--3966
		x"16",	--3967
		x"0c",	--3968
		x"0d",	--3969
		x"0e",	--3970
		x"0f",	--3971
		x"b0",	--3972
		x"b2",	--3973
		x"3c",	--3974
		x"35",	--3975
		x"3d",	--3976
		x"88",	--3977
		x"b0",	--3978
		x"16",	--3979
		x"0c",	--3980
		x"0d",	--3981
		x"0e",	--3982
		x"0f",	--3983
		x"b0",	--3984
		x"b2",	--3985
		x"3c",	--3986
		x"6e",	--3987
		x"3d",	--3988
		x"ba",	--3989
		x"b0",	--3990
		x"16",	--3991
		x"0c",	--3992
		x"0d",	--3993
		x"0e",	--3994
		x"0f",	--3995
		x"b0",	--3996
		x"b2",	--3997
		x"3c",	--3998
		x"25",	--3999
		x"3d",	--4000
		x"12",	--4001
		x"b0",	--4002
		x"16",	--4003
		x"0c",	--4004
		x"0d",	--4005
		x"0e",	--4006
		x"0f",	--4007
		x"b0",	--4008
		x"b2",	--4009
		x"3c",	--4010
		x"ab",	--4011
		x"3d",	--4012
		x"aa",	--4013
		x"b0",	--4014
		x"16",	--4015
		x"0c",	--4016
		x"0d",	--4017
		x"0e",	--4018
		x"0f",	--4019
		x"b0",	--4020
		x"b2",	--4021
		x"81",	--4022
		x"04",	--4023
		x"81",	--4024
		x"06",	--4025
		x"3c",	--4026
		x"21",	--4027
		x"3d",	--4028
		x"15",	--4029
		x"0e",	--4030
		x"0f",	--4031
		x"b0",	--4032
		x"b2",	--4033
		x"3c",	--4034
		x"6b",	--4035
		x"3d",	--4036
		x"6e",	--4037
		x"b0",	--4038
		x"62",	--4039
		x"0c",	--4040
		x"0d",	--4041
		x"0e",	--4042
		x"0f",	--4043
		x"b0",	--4044
		x"b2",	--4045
		x"3c",	--4046
		x"95",	--4047
		x"3d",	--4048
		x"9d",	--4049
		x"b0",	--4050
		x"62",	--4051
		x"0c",	--4052
		x"0d",	--4053
		x"0e",	--4054
		x"0f",	--4055
		x"b0",	--4056
		x"b2",	--4057
		x"3c",	--4058
		x"38",	--4059
		x"3d",	--4060
		x"e3",	--4061
		x"b0",	--4062
		x"62",	--4063
		x"0c",	--4064
		x"0d",	--4065
		x"0e",	--4066
		x"0f",	--4067
		x"b0",	--4068
		x"b2",	--4069
		x"3c",	--4070
		x"cd",	--4071
		x"3d",	--4072
		x"4c",	--4073
		x"b0",	--4074
		x"62",	--4075
		x"0c",	--4076
		x"0d",	--4077
		x"0e",	--4078
		x"0f",	--4079
		x"b0",	--4080
		x"b2",	--4081
		x"08",	--4082
		x"09",	--4083
		x"36",	--4084
		x"19",	--4085
		x"37",	--4086
		x"17",	--4087
		x"0c",	--4088
		x"0d",	--4089
		x"1e",	--4090
		x"04",	--4091
		x"1f",	--4092
		x"06",	--4093
		x"b0",	--4094
		x"16",	--4095
		x"0c",	--4096
		x"0d",	--4097
		x"0e",	--4098
		x"0f",	--4099
		x"b0",	--4100
		x"b2",	--4101
		x"0c",	--4102
		x"0d",	--4103
		x"0e",	--4104
		x"0f",	--4105
		x"b0",	--4106
		x"62",	--4107
		x"04",	--4108
		x"05",	--4109
		x"31",	--4110
		x"0b",	--4111
		x"0b",	--4112
		x"0b",	--4113
		x"07",	--4114
		x"37",	--4115
		x"bc",	--4116
		x"0c",	--4117
		x"0d",	--4118
		x"1e",	--4119
		x"04",	--4120
		x"1f",	--4121
		x"06",	--4122
		x"b0",	--4123
		x"16",	--4124
		x"0c",	--4125
		x"0d",	--4126
		x"0e",	--4127
		x"0f",	--4128
		x"b0",	--4129
		x"b2",	--4130
		x"1c",	--4131
		x"cc",	--4132
		x"1d",	--4133
		x"ce",	--4134
		x"b0",	--4135
		x"62",	--4136
		x"0c",	--4137
		x"0d",	--4138
		x"b0",	--4139
		x"62",	--4140
		x"0c",	--4141
		x"0d",	--4142
		x"2e",	--4143
		x"1f",	--4144
		x"02",	--4145
		x"b0",	--4146
		x"62",	--4147
		x"04",	--4148
		x"05",	--4149
		x"81",	--4150
		x"02",	--4151
		x"07",	--4152
		x"35",	--4153
		x"00",	--4154
		x"04",	--4155
		x"34",	--4156
		x"db",	--4157
		x"35",	--4158
		x"c9",	--4159
		x"0e",	--4160
		x"0f",	--4161
		x"31",	--4162
		x"34",	--4163
		x"35",	--4164
		x"36",	--4165
		x"37",	--4166
		x"38",	--4167
		x"39",	--4168
		x"3a",	--4169
		x"3b",	--4170
		x"30",	--4171
		x"b0",	--4172
		x"44",	--4173
		x"30",	--4174
		x"0b",	--4175
		x"0a",	--4176
		x"31",	--4177
		x"0c",	--4178
		x"0d",	--4179
		x"3c",	--4180
		x"3d",	--4181
		x"ff",	--4182
		x"3d",	--4183
		x"49",	--4184
		x"06",	--4185
		x"3d",	--4186
		x"4a",	--4187
		x"07",	--4188
		x"3c",	--4189
		x"d9",	--4190
		x"04",	--4191
		x"03",	--4192
		x"0c",	--4193
		x"0d",	--4194
		x"27",	--4195
		x"3d",	--4196
		x"80",	--4197
		x"05",	--4198
		x"0c",	--4199
		x"0d",	--4200
		x"b0",	--4201
		x"62",	--4202
		x"2f",	--4203
		x"0d",	--4204
		x"b0",	--4205
		x"28",	--4206
		x"0a",	--4207
		x"0b",	--4208
		x"3a",	--4209
		x"03",	--4210
		x"0b",	--4211
		x"1c",	--4212
		x"04",	--4213
		x"1d",	--4214
		x"06",	--4215
		x"2e",	--4216
		x"1f",	--4217
		x"02",	--4218
		x"1a",	--4219
		x"02",	--4220
		x"0b",	--4221
		x"10",	--4222
		x"2a",	--4223
		x"02",	--4224
		x"0b",	--4225
		x"0f",	--4226
		x"2e",	--4227
		x"1f",	--4228
		x"02",	--4229
		x"0a",	--4230
		x"0f",	--4231
		x"0b",	--4232
		x"0d",	--4233
		x"13",	--4234
		x"b0",	--4235
		x"1e",	--4236
		x"21",	--4237
		x"0c",	--4238
		x"b0",	--4239
		x"44",	--4240
		x"09",	--4241
		x"13",	--4242
		x"b0",	--4243
		x"1e",	--4244
		x"21",	--4245
		x"02",	--4246
		x"b0",	--4247
		x"44",	--4248
		x"3f",	--4249
		x"00",	--4250
		x"31",	--4251
		x"3a",	--4252
		x"3b",	--4253
		x"30",	--4254
		x"b0",	--4255
		x"9e",	--4256
		x"30",	--4257
		x"0b",	--4258
		x"0a",	--4259
		x"09",	--4260
		x"08",	--4261
		x"07",	--4262
		x"06",	--4263
		x"05",	--4264
		x"04",	--4265
		x"31",	--4266
		x"06",	--4267
		x"07",	--4268
		x"04",	--4269
		x"05",	--4270
		x"0a",	--4271
		x"0b",	--4272
		x"3a",	--4273
		x"3b",	--4274
		x"ff",	--4275
		x"3b",	--4276
		x"00",	--4277
		x"04",	--4278
		x"b0",	--4279
		x"5c",	--4280
		x"0e",	--4281
		x"cc",	--4282
		x"0c",	--4283
		x"0d",	--4284
		x"0e",	--4285
		x"0f",	--4286
		x"b0",	--4287
		x"b2",	--4288
		x"08",	--4289
		x"09",	--4290
		x"3c",	--4291
		x"4e",	--4292
		x"3d",	--4293
		x"47",	--4294
		x"b0",	--4295
		x"b2",	--4296
		x"3c",	--4297
		x"f6",	--4298
		x"3d",	--4299
		x"0f",	--4300
		x"b0",	--4301
		x"16",	--4302
		x"0c",	--4303
		x"0d",	--4304
		x"0e",	--4305
		x"0f",	--4306
		x"b0",	--4307
		x"b2",	--4308
		x"3c",	--4309
		x"7c",	--4310
		x"3d",	--4311
		x"93",	--4312
		x"b0",	--4313
		x"62",	--4314
		x"0c",	--4315
		x"0d",	--4316
		x"0e",	--4317
		x"0f",	--4318
		x"b0",	--4319
		x"b2",	--4320
		x"3c",	--4321
		x"01",	--4322
		x"3d",	--4323
		x"d0",	--4324
		x"b0",	--4325
		x"16",	--4326
		x"0c",	--4327
		x"0d",	--4328
		x"0e",	--4329
		x"0f",	--4330
		x"b0",	--4331
		x"b2",	--4332
		x"3c",	--4333
		x"61",	--4334
		x"3d",	--4335
		x"b6",	--4336
		x"b0",	--4337
		x"62",	--4338
		x"0c",	--4339
		x"0d",	--4340
		x"0e",	--4341
		x"0f",	--4342
		x"b0",	--4343
		x"b2",	--4344
		x"3c",	--4345
		x"ab",	--4346
		x"3d",	--4347
		x"2a",	--4348
		x"b0",	--4349
		x"16",	--4350
		x"0c",	--4351
		x"0d",	--4352
		x"0e",	--4353
		x"0f",	--4354
		x"b0",	--4355
		x"b2",	--4356
		x"81",	--4357
		x"00",	--4358
		x"81",	--4359
		x"02",	--4360
		x"3b",	--4361
		x"99",	--4362
		x"06",	--4363
		x"3b",	--4364
		x"9a",	--4365
		x"2d",	--4366
		x"3a",	--4367
		x"9a",	--4368
		x"2a",	--4369
		x"0c",	--4370
		x"3d",	--4371
		x"00",	--4372
		x"0e",	--4373
		x"0f",	--4374
		x"b0",	--4375
		x"b2",	--4376
		x"0a",	--4377
		x"0b",	--4378
		x"2c",	--4379
		x"1d",	--4380
		x"02",	--4381
		x"0e",	--4382
		x"0f",	--4383
		x"b0",	--4384
		x"b2",	--4385
		x"08",	--4386
		x"09",	--4387
		x"0c",	--4388
		x"0d",	--4389
		x"0e",	--4390
		x"0f",	--4391
		x"b0",	--4392
		x"b2",	--4393
		x"0c",	--4394
		x"0d",	--4395
		x"0e",	--4396
		x"0f",	--4397
		x"b0",	--4398
		x"62",	--4399
		x"0c",	--4400
		x"0d",	--4401
		x"0e",	--4402
		x"0f",	--4403
		x"b0",	--4404
		x"62",	--4405
		x"0c",	--4406
		x"0d",	--4407
		x"0e",	--4408
		x"3f",	--4409
		x"80",	--4410
		x"48",	--4411
		x"3b",	--4412
		x"48",	--4413
		x"05",	--4414
		x"3b",	--4415
		x"49",	--4416
		x"06",	--4417
		x"1a",	--4418
		x"04",	--4419
		x"0a",	--4420
		x"3b",	--4421
		x"00",	--4422
		x"03",	--4423
		x"0a",	--4424
		x"3b",	--4425
		x"90",	--4426
		x"0c",	--4427
		x"0d",	--4428
		x"0e",	--4429
		x"3f",	--4430
		x"80",	--4431
		x"b0",	--4432
		x"62",	--4433
		x"81",	--4434
		x"04",	--4435
		x"81",	--4436
		x"06",	--4437
		x"0c",	--4438
		x"3d",	--4439
		x"00",	--4440
		x"0e",	--4441
		x"0f",	--4442
		x"b0",	--4443
		x"b2",	--4444
		x"0c",	--4445
		x"0d",	--4446
		x"b0",	--4447
		x"62",	--4448
		x"0a",	--4449
		x"0b",	--4450
		x"2c",	--4451
		x"1d",	--4452
		x"02",	--4453
		x"0e",	--4454
		x"0f",	--4455
		x"b0",	--4456
		x"b2",	--4457
		x"08",	--4458
		x"09",	--4459
		x"0c",	--4460
		x"0d",	--4461
		x"0e",	--4462
		x"0f",	--4463
		x"b0",	--4464
		x"b2",	--4465
		x"0c",	--4466
		x"0d",	--4467
		x"0e",	--4468
		x"0f",	--4469
		x"b0",	--4470
		x"62",	--4471
		x"0c",	--4472
		x"0d",	--4473
		x"0e",	--4474
		x"0f",	--4475
		x"b0",	--4476
		x"62",	--4477
		x"0c",	--4478
		x"0d",	--4479
		x"1e",	--4480
		x"04",	--4481
		x"1f",	--4482
		x"06",	--4483
		x"b0",	--4484
		x"62",	--4485
		x"03",	--4486
		x"0e",	--4487
		x"3f",	--4488
		x"80",	--4489
		x"31",	--4490
		x"34",	--4491
		x"35",	--4492
		x"36",	--4493
		x"37",	--4494
		x"38",	--4495
		x"39",	--4496
		x"3a",	--4497
		x"3b",	--4498
		x"30",	--4499
		x"0b",	--4500
		x"0a",	--4501
		x"09",	--4502
		x"08",	--4503
		x"07",	--4504
		x"06",	--4505
		x"05",	--4506
		x"04",	--4507
		x"31",	--4508
		x"de",	--4509
		x"81",	--4510
		x"0c",	--4511
		x"81",	--4512
		x"12",	--4513
		x"81",	--4514
		x"14",	--4515
		x"0a",	--4516
		x"0b",	--4517
		x"3a",	--4518
		x"3b",	--4519
		x"ff",	--4520
		x"3b",	--4521
		x"49",	--4522
		x"06",	--4523
		x"3b",	--4524
		x"4a",	--4525
		x"0f",	--4526
		x"3a",	--4527
		x"d9",	--4528
		x"0c",	--4529
		x"1d",	--4530
		x"0c",	--4531
		x"8d",	--4532
		x"00",	--4533
		x"8d",	--4534
		x"02",	--4535
		x"8d",	--4536
		x"04",	--4537
		x"8d",	--4538
		x"06",	--4539
		x"30",	--4540
		x"f4",	--4541
		x"3b",	--4542
		x"16",	--4543
		x"06",	--4544
		x"3b",	--4545
		x"17",	--4546
		x"b2",	--4547
		x"3a",	--4548
		x"e4",	--4549
		x"af",	--4550
		x"81",	--4551
		x"14",	--4552
		x"58",	--4553
		x"03",	--4554
		x"91",	--4555
		x"12",	--4556
		x"54",	--4557
		x"3c",	--4558
		x"80",	--4559
		x"3d",	--4560
		x"c9",	--4561
		x"b0",	--4562
		x"62",	--4563
		x"08",	--4564
		x"09",	--4565
		x"3a",	--4566
		x"f0",	--4567
		x"3b",	--4568
		x"3a",	--4569
		x"d0",	--4570
		x"03",	--4571
		x"3b",	--4572
		x"c9",	--4573
		x"19",	--4574
		x"3c",	--4575
		x"43",	--4576
		x"3d",	--4577
		x"35",	--4578
		x"0e",	--4579
		x"0f",	--4580
		x"b0",	--4581
		x"62",	--4582
		x"0c",	--4583
		x"0d",	--4584
		x"1f",	--4585
		x"0c",	--4586
		x"8f",	--4587
		x"00",	--4588
		x"8f",	--4589
		x"02",	--4590
		x"0e",	--4591
		x"0f",	--4592
		x"b0",	--4593
		x"62",	--4594
		x"3c",	--4595
		x"43",	--4596
		x"3d",	--4597
		x"35",	--4598
		x"1e",	--4599
		x"3c",	--4600
		x"00",	--4601
		x"3d",	--4602
		x"35",	--4603
		x"b0",	--4604
		x"62",	--4605
		x"0a",	--4606
		x"0b",	--4607
		x"3c",	--4608
		x"08",	--4609
		x"3d",	--4610
		x"85",	--4611
		x"b0",	--4612
		x"62",	--4613
		x"0c",	--4614
		x"0d",	--4615
		x"1e",	--4616
		x"0c",	--4617
		x"8e",	--4618
		x"00",	--4619
		x"8e",	--4620
		x"02",	--4621
		x"0e",	--4622
		x"0f",	--4623
		x"b0",	--4624
		x"62",	--4625
		x"3c",	--4626
		x"08",	--4627
		x"3d",	--4628
		x"85",	--4629
		x"b0",	--4630
		x"62",	--4631
		x"1d",	--4632
		x"0c",	--4633
		x"8d",	--4634
		x"04",	--4635
		x"8d",	--4636
		x"06",	--4637
		x"16",	--4638
		x"07",	--4639
		x"30",	--4640
		x"ee",	--4641
		x"3c",	--4642
		x"80",	--4643
		x"3d",	--4644
		x"c9",	--4645
		x"b0",	--4646
		x"16",	--4647
		x"08",	--4648
		x"09",	--4649
		x"3a",	--4650
		x"f0",	--4651
		x"3b",	--4652
		x"3a",	--4653
		x"d0",	--4654
		x"03",	--4655
		x"3b",	--4656
		x"c9",	--4657
		x"19",	--4658
		x"3c",	--4659
		x"43",	--4660
		x"3d",	--4661
		x"35",	--4662
		x"0e",	--4663
		x"0f",	--4664
		x"b0",	--4665
		x"16",	--4666
		x"0c",	--4667
		x"0d",	--4668
		x"1e",	--4669
		x"0c",	--4670
		x"8e",	--4671
		x"00",	--4672
		x"8e",	--4673
		x"02",	--4674
		x"0e",	--4675
		x"0f",	--4676
		x"b0",	--4677
		x"62",	--4678
		x"3c",	--4679
		x"43",	--4680
		x"3d",	--4681
		x"35",	--4682
		x"1e",	--4683
		x"3c",	--4684
		x"00",	--4685
		x"3d",	--4686
		x"35",	--4687
		x"b0",	--4688
		x"16",	--4689
		x"0a",	--4690
		x"0b",	--4691
		x"3c",	--4692
		x"08",	--4693
		x"3d",	--4694
		x"85",	--4695
		x"b0",	--4696
		x"16",	--4697
		x"0c",	--4698
		x"0d",	--4699
		x"1e",	--4700
		x"0c",	--4701
		x"8e",	--4702
		x"00",	--4703
		x"8e",	--4704
		x"02",	--4705
		x"0e",	--4706
		x"0f",	--4707
		x"b0",	--4708
		x"62",	--4709
		x"3c",	--4710
		x"08",	--4711
		x"3d",	--4712
		x"85",	--4713
		x"b0",	--4714
		x"16",	--4715
		x"1d",	--4716
		x"0c",	--4717
		x"8d",	--4718
		x"04",	--4719
		x"8d",	--4720
		x"06",	--4721
		x"36",	--4722
		x"37",	--4723
		x"30",	--4724
		x"ee",	--4725
		x"3b",	--4726
		x"49",	--4727
		x"0a",	--4728
		x"3b",	--4729
		x"4a",	--4730
		x"02",	--4731
		x"30",	--4732
		x"d2",	--4733
		x"3a",	--4734
		x"81",	--4735
		x"02",	--4736
		x"30",	--4737
		x"d2",	--4738
		x"08",	--4739
		x"09",	--4740
		x"39",	--4741
		x"ff",	--4742
		x"3c",	--4743
		x"84",	--4744
		x"3d",	--4745
		x"22",	--4746
		x"0e",	--4747
		x"0f",	--4748
		x"b0",	--4749
		x"b2",	--4750
		x"0c",	--4751
		x"3d",	--4752
		x"00",	--4753
		x"b0",	--4754
		x"16",	--4755
		x"b0",	--4756
		x"5c",	--4757
		x"06",	--4758
		x"07",	--4759
		x"b0",	--4760
		x"b6",	--4761
		x"81",	--4762
		x"1a",	--4763
		x"81",	--4764
		x"1c",	--4765
		x"3c",	--4766
		x"80",	--4767
		x"3d",	--4768
		x"c9",	--4769
		x"b0",	--4770
		x"b2",	--4771
		x"0c",	--4772
		x"0d",	--4773
		x"0e",	--4774
		x"0f",	--4775
		x"b0",	--4776
		x"62",	--4777
		x"04",	--4778
		x"05",	--4779
		x"3c",	--4780
		x"43",	--4781
		x"3d",	--4782
		x"35",	--4783
		x"1e",	--4784
		x"1a",	--4785
		x"1f",	--4786
		x"1c",	--4787
		x"b0",	--4788
		x"b2",	--4789
		x"81",	--4790
		x"0e",	--4791
		x"81",	--4792
		x"10",	--4793
		x"07",	--4794
		x"05",	--4795
		x"17",	--4796
		x"19",	--4797
		x"36",	--4798
		x"20",	--4799
		x"16",	--4800
		x"08",	--4801
		x"09",	--4802
		x"38",	--4803
		x"00",	--4804
		x"39",	--4805
		x"0f",	--4806
		x"3f",	--4807
		x"0f",	--4808
		x"0f",	--4809
		x"3f",	--4810
		x"dc",	--4811
		x"28",	--4812
		x"03",	--4813
		x"19",	--4814
		x"02",	--4815
		x"06",	--4816
		x"1c",	--4817
		x"0e",	--4818
		x"1d",	--4819
		x"10",	--4820
		x"30",	--4821
		x"5a",	--4822
		x"1c",	--4823
		x"0e",	--4824
		x"1d",	--4825
		x"10",	--4826
		x"0e",	--4827
		x"0f",	--4828
		x"b0",	--4829
		x"62",	--4830
		x"08",	--4831
		x"09",	--4832
		x"1e",	--4833
		x"0c",	--4834
		x"8e",	--4835
		x"00",	--4836
		x"8e",	--4837
		x"02",	--4838
		x"81",	--4839
		x"16",	--4840
		x"0d",	--4841
		x"8d",	--4842
		x"8d",	--4843
		x"8d",	--4844
		x"8d",	--4845
		x"81",	--4846
		x"18",	--4847
		x"7d",	--4848
		x"07",	--4849
		x"0c",	--4850
		x"1e",	--4851
		x"16",	--4852
		x"1f",	--4853
		x"18",	--4854
		x"0f",	--4855
		x"0e",	--4856
		x"7d",	--4857
		x"fc",	--4858
		x"81",	--4859
		x"16",	--4860
		x"81",	--4861
		x"18",	--4862
		x"0a",	--4863
		x"0b",	--4864
		x"7f",	--4865
		x"07",	--4866
		x"12",	--4867
		x"0b",	--4868
		x"0a",	--4869
		x"7f",	--4870
		x"fb",	--4871
		x"3a",	--4872
		x"ff",	--4873
		x"0b",	--4874
		x"18",	--4875
		x"16",	--4876
		x"19",	--4877
		x"18",	--4878
		x"08",	--4879
		x"09",	--4880
		x"09",	--4881
		x"a9",	--4882
		x"03",	--4883
		x"38",	--4884
		x"09",	--4885
		x"a5",	--4886
		x"3c",	--4887
		x"00",	--4888
		x"3d",	--4889
		x"35",	--4890
		x"1e",	--4891
		x"1a",	--4892
		x"1f",	--4893
		x"1c",	--4894
		x"b0",	--4895
		x"b2",	--4896
		x"08",	--4897
		x"09",	--4898
		x"0c",	--4899
		x"0d",	--4900
		x"0e",	--4901
		x"0f",	--4902
		x"b0",	--4903
		x"62",	--4904
		x"81",	--4905
		x"1e",	--4906
		x"81",	--4907
		x"20",	--4908
		x"0c",	--4909
		x"0d",	--4910
		x"0e",	--4911
		x"0f",	--4912
		x"b0",	--4913
		x"62",	--4914
		x"0c",	--4915
		x"0d",	--4916
		x"b0",	--4917
		x"62",	--4918
		x"08",	--4919
		x"09",	--4920
		x"3c",	--4921
		x"08",	--4922
		x"3d",	--4923
		x"85",	--4924
		x"1e",	--4925
		x"1a",	--4926
		x"1f",	--4927
		x"1c",	--4928
		x"b0",	--4929
		x"b2",	--4930
		x"0c",	--4931
		x"0d",	--4932
		x"b0",	--4933
		x"62",	--4934
		x"81",	--4935
		x"0e",	--4936
		x"81",	--4937
		x"10",	--4938
		x"0c",	--4939
		x"0d",	--4940
		x"1e",	--4941
		x"1e",	--4942
		x"1f",	--4943
		x"20",	--4944
		x"b0",	--4945
		x"62",	--4946
		x"0a",	--4947
		x"0b",	--4948
		x"1e",	--4949
		x"0c",	--4950
		x"8e",	--4951
		x"00",	--4952
		x"8e",	--4953
		x"02",	--4954
		x"0a",	--4955
		x"0b",	--4956
		x"7f",	--4957
		x"07",	--4958
		x"12",	--4959
		x"0b",	--4960
		x"0a",	--4961
		x"7f",	--4962
		x"fb",	--4963
		x"3a",	--4964
		x"ff",	--4965
		x"0b",	--4966
		x"1d",	--4967
		x"16",	--4968
		x"1e",	--4969
		x"18",	--4970
		x"0d",	--4971
		x"0e",	--4972
		x"0a",	--4973
		x"0b",	--4974
		x"0b",	--4975
		x"47",	--4976
		x"03",	--4977
		x"3d",	--4978
		x"1a",	--4979
		x"43",	--4980
		x"3c",	--4981
		x"00",	--4982
		x"3d",	--4983
		x"85",	--4984
		x"1e",	--4985
		x"1a",	--4986
		x"1f",	--4987
		x"1c",	--4988
		x"b0",	--4989
		x"b2",	--4990
		x"0a",	--4991
		x"0b",	--4992
		x"0c",	--4993
		x"0d",	--4994
		x"1e",	--4995
		x"1e",	--4996
		x"1f",	--4997
		x"20",	--4998
		x"b0",	--4999
		x"62",	--5000
		x"04",	--5001
		x"05",	--5002
		x"0c",	--5003
		x"0d",	--5004
		x"1e",	--5005
		x"1e",	--5006
		x"1f",	--5007
		x"20",	--5008
		x"b0",	--5009
		x"62",	--5010
		x"0c",	--5011
		x"0d",	--5012
		x"b0",	--5013
		x"62",	--5014
		x"0a",	--5015
		x"0b",	--5016
		x"3c",	--5017
		x"32",	--5018
		x"3d",	--5019
		x"8d",	--5020
		x"1e",	--5021
		x"1a",	--5022
		x"1f",	--5023
		x"1c",	--5024
		x"b0",	--5025
		x"b2",	--5026
		x"0c",	--5027
		x"0d",	--5028
		x"b0",	--5029
		x"62",	--5030
		x"81",	--5031
		x"0e",	--5032
		x"81",	--5033
		x"10",	--5034
		x"0c",	--5035
		x"0d",	--5036
		x"0e",	--5037
		x"0f",	--5038
		x"b0",	--5039
		x"62",	--5040
		x"1d",	--5041
		x"0c",	--5042
		x"8d",	--5043
		x"00",	--5044
		x"8d",	--5045
		x"02",	--5046
		x"04",	--5047
		x"14",	--5048
		x"1e",	--5049
		x"15",	--5050
		x"20",	--5051
		x"1e",	--5052
		x"0c",	--5053
		x"28",	--5054
		x"19",	--5055
		x"02",	--5056
		x"0c",	--5057
		x"0d",	--5058
		x"0e",	--5059
		x"0f",	--5060
		x"b0",	--5061
		x"62",	--5062
		x"1c",	--5063
		x"0e",	--5064
		x"1d",	--5065
		x"10",	--5066
		x"b0",	--5067
		x"62",	--5068
		x"0a",	--5069
		x"0b",	--5070
		x"1f",	--5071
		x"0c",	--5072
		x"8f",	--5073
		x"04",	--5074
		x"8f",	--5075
		x"06",	--5076
		x"81",	--5077
		x"14",	--5078
		x"9f",	--5079
		x"0d",	--5080
		x"0e",	--5081
		x"3e",	--5082
		x"00",	--5083
		x"8f",	--5084
		x"00",	--5085
		x"8f",	--5086
		x"02",	--5087
		x"0d",	--5088
		x"0e",	--5089
		x"3e",	--5090
		x"00",	--5091
		x"8f",	--5092
		x"04",	--5093
		x"8f",	--5094
		x"06",	--5095
		x"8a",	--5096
		x"3b",	--5097
		x"80",	--5098
		x"11",	--5099
		x"0c",	--5100
		x"0d",	--5101
		x"b0",	--5102
		x"62",	--5103
		x"1d",	--5104
		x"0c",	--5105
		x"8d",	--5106
		x"04",	--5107
		x"8d",	--5108
		x"06",	--5109
		x"8d",	--5110
		x"00",	--5111
		x"8d",	--5112
		x"02",	--5113
		x"06",	--5114
		x"07",	--5115
		x"7a",	--5116
		x"0c",	--5117
		x"0d",	--5118
		x"8d",	--5119
		x"8d",	--5120
		x"8d",	--5121
		x"8d",	--5122
		x"7f",	--5123
		x"07",	--5124
		x"0d",	--5125
		x"0c",	--5126
		x"7f",	--5127
		x"fc",	--5128
		x"09",	--5129
		x"39",	--5130
		x"7a",	--5131
		x"0c",	--5132
		x"0d",	--5133
		x"0d",	--5134
		x"7f",	--5135
		x"07",	--5136
		x"0c",	--5137
		x"0d",	--5138
		x"7f",	--5139
		x"fc",	--5140
		x"0a",	--5141
		x"0b",	--5142
		x"0e",	--5143
		x"0f",	--5144
		x"b0",	--5145
		x"5c",	--5146
		x"b0",	--5147
		x"b6",	--5148
		x"0c",	--5149
		x"0d",	--5150
		x"81",	--5151
		x"00",	--5152
		x"81",	--5153
		x"02",	--5154
		x"0e",	--5155
		x"0f",	--5156
		x"b0",	--5157
		x"62",	--5158
		x"0c",	--5159
		x"3d",	--5160
		x"80",	--5161
		x"b0",	--5162
		x"b2",	--5163
		x"0a",	--5164
		x"0b",	--5165
		x"b0",	--5166
		x"5c",	--5167
		x"b0",	--5168
		x"b6",	--5169
		x"0c",	--5170
		x"0d",	--5171
		x"81",	--5172
		x"04",	--5173
		x"81",	--5174
		x"06",	--5175
		x"0e",	--5176
		x"0f",	--5177
		x"b0",	--5178
		x"62",	--5179
		x"0c",	--5180
		x"3d",	--5181
		x"80",	--5182
		x"b0",	--5183
		x"b2",	--5184
		x"81",	--5185
		x"08",	--5186
		x"81",	--5187
		x"0a",	--5188
		x"08",	--5189
		x"38",	--5190
		x"3a",	--5191
		x"03",	--5192
		x"01",	--5193
		x"3a",	--5194
		x"28",	--5195
		x"0c",	--5196
		x"0d",	--5197
		x"1e",	--5198
		x"04",	--5199
		x"1f",	--5200
		x"06",	--5201
		x"b0",	--5202
		x"26",	--5203
		x"0f",	--5204
		x"f4",	--5205
		x"30",	--5206
		x"5c",	--5207
		x"23",	--5208
		x"0c",	--5209
		x"0d",	--5210
		x"1e",	--5211
		x"10",	--5212
		x"0f",	--5213
		x"2f",	--5214
		x"b0",	--5215
		x"08",	--5216
		x"21",	--5217
		x"06",	--5218
		x"8f",	--5219
		x"8f",	--5220
		x"8f",	--5221
		x"8f",	--5222
		x"07",	--5223
		x"81",	--5224
		x"14",	--5225
		x"0c",	--5226
		x"1e",	--5227
		x"0c",	--5228
		x"be",	--5229
		x"00",	--5230
		x"02",	--5231
		x"be",	--5232
		x"00",	--5233
		x"06",	--5234
		x"36",	--5235
		x"37",	--5236
		x"16",	--5237
		x"07",	--5238
		x"0e",	--5239
		x"0f",	--5240
		x"31",	--5241
		x"22",	--5242
		x"34",	--5243
		x"35",	--5244
		x"36",	--5245
		x"37",	--5246
		x"38",	--5247
		x"39",	--5248
		x"3a",	--5249
		x"3b",	--5250
		x"30",	--5251
		x"0b",	--5252
		x"0a",	--5253
		x"09",	--5254
		x"08",	--5255
		x"07",	--5256
		x"06",	--5257
		x"05",	--5258
		x"04",	--5259
		x"31",	--5260
		x"8c",	--5261
		x"81",	--5262
		x"66",	--5263
		x"81",	--5264
		x"60",	--5265
		x"81",	--5266
		x"48",	--5267
		x"1a",	--5268
		x"86",	--5269
		x"0a",	--5270
		x"81",	--5271
		x"4c",	--5272
		x"81",	--5273
		x"4e",	--5274
		x"91",	--5275
		x"74",	--5276
		x"4c",	--5277
		x"1a",	--5278
		x"4c",	--5279
		x"8a",	--5280
		x"8a",	--5281
		x"8a",	--5282
		x"8a",	--5283
		x"81",	--5284
		x"4e",	--5285
		x"0a",	--5286
		x"3a",	--5287
		x"81",	--5288
		x"50",	--5289
		x"8a",	--5290
		x"8a",	--5291
		x"8a",	--5292
		x"8a",	--5293
		x"81",	--5294
		x"52",	--5295
		x"0a",	--5296
		x"3a",	--5297
		x"fd",	--5298
		x"0a",	--5299
		x"02",	--5300
		x"3a",	--5301
		x"07",	--5302
		x"0a",	--5303
		x"0a",	--5304
		x"0a",	--5305
		x"08",	--5306
		x"88",	--5307
		x"88",	--5308
		x"88",	--5309
		x"88",	--5310
		x"81",	--5311
		x"54",	--5312
		x"81",	--5313
		x"56",	--5314
		x"04",	--5315
		x"81",	--5316
		x"54",	--5317
		x"81",	--5318
		x"56",	--5319
		x"08",	--5320
		x"8d",	--5321
		x"8d",	--5322
		x"8d",	--5323
		x"8d",	--5324
		x"09",	--5325
		x"1a",	--5326
		x"54",	--5327
		x"1b",	--5328
		x"56",	--5329
		x"3a",	--5330
		x"3b",	--5331
		x"0a",	--5332
		x"0b",	--5333
		x"0a",	--5334
		x"0b",	--5335
		x"0a",	--5336
		x"0b",	--5337
		x"0d",	--5338
		x"0e",	--5339
		x"0d",	--5340
		x"0e",	--5341
		x"81",	--5342
		x"44",	--5343
		x"81",	--5344
		x"46",	--5345
		x"18",	--5346
		x"54",	--5347
		x"19",	--5348
		x"56",	--5349
		x"18",	--5350
		x"50",	--5351
		x"19",	--5352
		x"52",	--5353
		x"81",	--5354
		x"40",	--5355
		x"81",	--5356
		x"42",	--5357
		x"14",	--5358
		x"50",	--5359
		x"15",	--5360
		x"52",	--5361
		x"14",	--5362
		x"4c",	--5363
		x"15",	--5364
		x"4e",	--5365
		x"09",	--5366
		x"06",	--5367
		x"07",	--5368
		x"22",	--5369
		x"1e",	--5370
		x"40",	--5371
		x"1f",	--5372
		x"42",	--5373
		x"0e",	--5374
		x"0f",	--5375
		x"0f",	--5376
		x"0d",	--5377
		x"1f",	--5378
		x"40",	--5379
		x"0f",	--5380
		x"0f",	--5381
		x"1f",	--5382
		x"88",	--5383
		x"0f",	--5384
		x"2e",	--5385
		x"1f",	--5386
		x"02",	--5387
		x"b0",	--5388
		x"b6",	--5389
		x"02",	--5390
		x"0e",	--5391
		x"0f",	--5392
		x"3d",	--5393
		x"a0",	--5394
		x"0d",	--5395
		x"0d",	--5396
		x"8d",	--5397
		x"00",	--5398
		x"8d",	--5399
		x"02",	--5400
		x"16",	--5401
		x"07",	--5402
		x"29",	--5403
		x"05",	--5404
		x"04",	--5405
		x"07",	--5406
		x"da",	--5407
		x"04",	--5408
		x"d8",	--5409
		x"81",	--5410
		x"40",	--5411
		x"81",	--5412
		x"42",	--5413
		x"04",	--5414
		x"2d",	--5415
		x"1f",	--5416
		x"48",	--5417
		x"3f",	--5418
		x"0f",	--5419
		x"0f",	--5420
		x"3f",	--5421
		x"a0",	--5422
		x"0f",	--5423
		x"0f",	--5424
		x"2c",	--5425
		x"1d",	--5426
		x"02",	--5427
		x"3e",	--5428
		x"3f",	--5429
		x"b0",	--5430
		x"b2",	--5431
		x"0c",	--5432
		x"0d",	--5433
		x"0e",	--5434
		x"0f",	--5435
		x"b0",	--5436
		x"16",	--5437
		x"0a",	--5438
		x"0b",	--5439
		x"18",	--5440
		x"09",	--5441
		x"25",	--5442
		x"81",	--5443
		x"52",	--5444
		x"06",	--5445
		x"19",	--5446
		x"52",	--5447
		x"df",	--5448
		x"81",	--5449
		x"50",	--5450
		x"dc",	--5451
		x"84",	--5452
		x"00",	--5453
		x"84",	--5454
		x"02",	--5455
		x"91",	--5456
		x"40",	--5457
		x"81",	--5458
		x"42",	--5459
		x"24",	--5460
		x"91",	--5461
		x"42",	--5462
		x"4e",	--5463
		x"08",	--5464
		x"91",	--5465
		x"4e",	--5466
		x"42",	--5467
		x"15",	--5468
		x"91",	--5469
		x"40",	--5470
		x"4c",	--5471
		x"11",	--5472
		x"91",	--5473
		x"4c",	--5474
		x"40",	--5475
		x"91",	--5476
		x"4e",	--5477
		x"42",	--5478
		x"19",	--5479
		x"4c",	--5480
		x"1a",	--5481
		x"4e",	--5482
		x"39",	--5483
		x"3a",	--5484
		x"81",	--5485
		x"70",	--5486
		x"81",	--5487
		x"72",	--5488
		x"08",	--5489
		x"17",	--5490
		x"66",	--5491
		x"05",	--5492
		x"0a",	--5493
		x"0b",	--5494
		x"08",	--5495
		x"09",	--5496
		x"c9",	--5497
		x"1f",	--5498
		x"40",	--5499
		x"0f",	--5500
		x"0f",	--5501
		x"0f",	--5502
		x"28",	--5503
		x"19",	--5504
		x"02",	--5505
		x"0a",	--5506
		x"3a",	--5507
		x"f0",	--5508
		x"81",	--5509
		x"62",	--5510
		x"16",	--5511
		x"40",	--5512
		x"17",	--5513
		x"42",	--5514
		x"81",	--5515
		x"48",	--5516
		x"04",	--5517
		x"05",	--5518
		x"34",	--5519
		x"35",	--5520
		x"81",	--5521
		x"58",	--5522
		x"81",	--5523
		x"5a",	--5524
		x"05",	--5525
		x"32",	--5526
		x"0c",	--5527
		x"3d",	--5528
		x"80",	--5529
		x"0e",	--5530
		x"0f",	--5531
		x"b0",	--5532
		x"b2",	--5533
		x"b0",	--5534
		x"5c",	--5535
		x"b0",	--5536
		x"b6",	--5537
		x"0a",	--5538
		x"0b",	--5539
		x"0c",	--5540
		x"3d",	--5541
		x"80",	--5542
		x"b0",	--5543
		x"b2",	--5544
		x"0c",	--5545
		x"0d",	--5546
		x"0e",	--5547
		x"0f",	--5548
		x"b0",	--5549
		x"62",	--5550
		x"b0",	--5551
		x"5c",	--5552
		x"85",	--5553
		x"00",	--5554
		x"85",	--5555
		x"02",	--5556
		x"1f",	--5557
		x"58",	--5558
		x"0f",	--5559
		x"0f",	--5560
		x"0f",	--5561
		x"1f",	--5562
		x"48",	--5563
		x"1c",	--5564
		x"04",	--5565
		x"1d",	--5566
		x"06",	--5567
		x"0e",	--5568
		x"0f",	--5569
		x"b0",	--5570
		x"16",	--5571
		x"08",	--5572
		x"09",	--5573
		x"36",	--5574
		x"37",	--5575
		x"25",	--5576
		x"a1",	--5577
		x"48",	--5578
		x"07",	--5579
		x"04",	--5580
		x"17",	--5581
		x"c8",	--5582
		x"16",	--5583
		x"c6",	--5584
		x"91",	--5585
		x"44",	--5586
		x"5c",	--5587
		x"1d",	--5588
		x"44",	--5589
		x"0e",	--5590
		x"0f",	--5591
		x"b0",	--5592
		x"a2",	--5593
		x"0a",	--5594
		x"0b",	--5595
		x"0c",	--5596
		x"3d",	--5597
		x"00",	--5598
		x"b0",	--5599
		x"b2",	--5600
		x"b0",	--5601
		x"26",	--5602
		x"0c",	--5603
		x"3d",	--5604
		x"00",	--5605
		x"b0",	--5606
		x"b2",	--5607
		x"0c",	--5608
		x"0d",	--5609
		x"0e",	--5610
		x"0f",	--5611
		x"b0",	--5612
		x"62",	--5613
		x"0a",	--5614
		x"0b",	--5615
		x"b0",	--5616
		x"5c",	--5617
		x"81",	--5618
		x"58",	--5619
		x"81",	--5620
		x"5a",	--5621
		x"b0",	--5622
		x"b6",	--5623
		x"0c",	--5624
		x"0d",	--5625
		x"0e",	--5626
		x"0f",	--5627
		x"b0",	--5628
		x"62",	--5629
		x"81",	--5630
		x"48",	--5631
		x"81",	--5632
		x"4a",	--5633
		x"81",	--5634
		x"46",	--5635
		x"46",	--5636
		x"03",	--5637
		x"91",	--5638
		x"44",	--5639
		x"42",	--5640
		x"1c",	--5641
		x"40",	--5642
		x"1d",	--5643
		x"42",	--5644
		x"3c",	--5645
		x"3d",	--5646
		x"0b",	--5647
		x"0b",	--5648
		x"0b",	--5649
		x"0b",	--5650
		x"16",	--5651
		x"f0",	--5652
		x"17",	--5653
		x"f2",	--5654
		x"1e",	--5655
		x"44",	--5656
		x"39",	--5657
		x"09",	--5658
		x"0a",	--5659
		x"0b",	--5660
		x"48",	--5661
		x"78",	--5662
		x"1f",	--5663
		x"48",	--5664
		x"04",	--5665
		x"0b",	--5666
		x"0a",	--5667
		x"78",	--5668
		x"fa",	--5669
		x"81",	--5670
		x"58",	--5671
		x"81",	--5672
		x"5a",	--5673
		x"79",	--5674
		x"1f",	--5675
		x"49",	--5676
		x"04",	--5677
		x"0a",	--5678
		x"0b",	--5679
		x"79",	--5680
		x"fa",	--5681
		x"08",	--5682
		x"09",	--5683
		x"08",	--5684
		x"09",	--5685
		x"0f",	--5686
		x"0f",	--5687
		x"0f",	--5688
		x"0f",	--5689
		x"8f",	--5690
		x"f0",	--5691
		x"8f",	--5692
		x"f2",	--5693
		x"06",	--5694
		x"07",	--5695
		x"3f",	--5696
		x"07",	--5697
		x"4f",	--5698
		x"7f",	--5699
		x"1f",	--5700
		x"4f",	--5701
		x"28",	--5702
		x"07",	--5703
		x"06",	--5704
		x"7f",	--5705
		x"fa",	--5706
		x"81",	--5707
		x"44",	--5708
		x"13",	--5709
		x"81",	--5710
		x"46",	--5711
		x"10",	--5712
		x"1f",	--5713
		x"40",	--5714
		x"3f",	--5715
		x"0f",	--5716
		x"0f",	--5717
		x"0f",	--5718
		x"16",	--5719
		x"f0",	--5720
		x"17",	--5721
		x"f2",	--5722
		x"86",	--5723
		x"87",	--5724
		x"46",	--5725
		x"06",	--5726
		x"87",	--5727
		x"0e",	--5728
		x"0c",	--5729
		x"3d",	--5730
		x"00",	--5731
		x"1e",	--5732
		x"48",	--5733
		x"1f",	--5734
		x"4a",	--5735
		x"b0",	--5736
		x"c6",	--5737
		x"0f",	--5738
		x"09",	--5739
		x"06",	--5740
		x"07",	--5741
		x"94",	--5742
		x"07",	--5743
		x"92",	--5744
		x"05",	--5745
		x"16",	--5746
		x"8f",	--5747
		x"02",	--5748
		x"26",	--5749
		x"07",	--5750
		x"91",	--5751
		x"58",	--5752
		x"81",	--5753
		x"5a",	--5754
		x"04",	--5755
		x"05",	--5756
		x"08",	--5757
		x"09",	--5758
		x"1b",	--5759
		x"62",	--5760
		x"27",	--5761
		x"2c",	--5762
		x"1d",	--5763
		x"02",	--5764
		x"08",	--5765
		x"12",	--5766
		x"09",	--5767
		x"10",	--5768
		x"0c",	--5769
		x"02",	--5770
		x"0d",	--5771
		x"19",	--5772
		x"3e",	--5773
		x"00",	--5774
		x"0f",	--5775
		x"09",	--5776
		x"0a",	--5777
		x"09",	--5778
		x"0a",	--5779
		x"8b",	--5780
		x"00",	--5781
		x"8b",	--5782
		x"02",	--5783
		x"0b",	--5784
		x"3e",	--5785
		x"ff",	--5786
		x"0f",	--5787
		x"08",	--5788
		x"09",	--5789
		x"08",	--5790
		x"09",	--5791
		x"8b",	--5792
		x"00",	--5793
		x"8b",	--5794
		x"02",	--5795
		x"18",	--5796
		x"09",	--5797
		x"14",	--5798
		x"05",	--5799
		x"2b",	--5800
		x"15",	--5801
		x"42",	--5802
		x"d6",	--5803
		x"03",	--5804
		x"14",	--5805
		x"40",	--5806
		x"d2",	--5807
		x"81",	--5808
		x"46",	--5809
		x"28",	--5810
		x"03",	--5811
		x"91",	--5812
		x"44",	--5813
		x"24",	--5814
		x"91",	--5815
		x"44",	--5816
		x"03",	--5817
		x"81",	--5818
		x"46",	--5819
		x"07",	--5820
		x"a1",	--5821
		x"44",	--5822
		x"1b",	--5823
		x"81",	--5824
		x"46",	--5825
		x"0d",	--5826
		x"17",	--5827
		x"1f",	--5828
		x"40",	--5829
		x"3f",	--5830
		x"0f",	--5831
		x"0f",	--5832
		x"0f",	--5833
		x"bf",	--5834
		x"7f",	--5835
		x"f0",	--5836
		x"8f",	--5837
		x"f2",	--5838
		x"0b",	--5839
		x"1f",	--5840
		x"40",	--5841
		x"3f",	--5842
		x"0f",	--5843
		x"0f",	--5844
		x"0f",	--5845
		x"bf",	--5846
		x"3f",	--5847
		x"f0",	--5848
		x"8f",	--5849
		x"f2",	--5850
		x"26",	--5851
		x"26",	--5852
		x"07",	--5853
		x"24",	--5854
		x"1c",	--5855
		x"48",	--5856
		x"1d",	--5857
		x"4a",	--5858
		x"0e",	--5859
		x"3f",	--5860
		x"80",	--5861
		x"b0",	--5862
		x"62",	--5863
		x"81",	--5864
		x"48",	--5865
		x"81",	--5866
		x"4a",	--5867
		x"08",	--5868
		x"02",	--5869
		x"09",	--5870
		x"13",	--5871
		x"1d",	--5872
		x"5c",	--5873
		x"0e",	--5874
		x"3f",	--5875
		x"80",	--5876
		x"b0",	--5877
		x"a2",	--5878
		x"0c",	--5879
		x"0d",	--5880
		x"1e",	--5881
		x"48",	--5882
		x"1f",	--5883
		x"4a",	--5884
		x"b0",	--5885
		x"62",	--5886
		x"81",	--5887
		x"48",	--5888
		x"81",	--5889
		x"4a",	--5890
		x"0c",	--5891
		x"0d",	--5892
		x"1e",	--5893
		x"48",	--5894
		x"1f",	--5895
		x"4a",	--5896
		x"b0",	--5897
		x"26",	--5898
		x"0f",	--5899
		x"d7",	--5900
		x"1a",	--5901
		x"40",	--5902
		x"1b",	--5903
		x"42",	--5904
		x"3a",	--5905
		x"3b",	--5906
		x"1c",	--5907
		x"40",	--5908
		x"1d",	--5909
		x"42",	--5910
		x"09",	--5911
		x"81",	--5912
		x"5c",	--5913
		x"81",	--5914
		x"5e",	--5915
		x"0e",	--5916
		x"0f",	--5917
		x"0f",	--5918
		x"0f",	--5919
		x"3e",	--5920
		x"f0",	--5921
		x"0e",	--5922
		x"0f",	--5923
		x"0f",	--5924
		x"91",	--5925
		x"04",	--5926
		x"5c",	--5927
		x"91",	--5928
		x"06",	--5929
		x"5e",	--5930
		x"3c",	--5931
		x"3d",	--5932
		x"29",	--5933
		x"1d",	--5934
		x"4e",	--5935
		x"06",	--5936
		x"81",	--5937
		x"4e",	--5938
		x"e9",	--5939
		x"1c",	--5940
		x"4c",	--5941
		x"e6",	--5942
		x"81",	--5943
		x"5c",	--5944
		x"c3",	--5945
		x"81",	--5946
		x"5e",	--5947
		x"06",	--5948
		x"bf",	--5949
		x"91",	--5950
		x"62",	--5951
		x"81",	--5952
		x"64",	--5953
		x"05",	--5954
		x"0e",	--5955
		x"91",	--5956
		x"62",	--5957
		x"81",	--5958
		x"64",	--5959
		x"2e",	--5960
		x"1f",	--5961
		x"70",	--5962
		x"0f",	--5963
		x"0f",	--5964
		x"38",	--5965
		x"f0",	--5966
		x"08",	--5967
		x"0f",	--5968
		x"0f",	--5969
		x"8f",	--5970
		x"04",	--5971
		x"03",	--5972
		x"8f",	--5973
		x"06",	--5974
		x"e6",	--5975
		x"19",	--5976
		x"40",	--5977
		x"1a",	--5978
		x"42",	--5979
		x"19",	--5980
		x"0a",	--5981
		x"81",	--5982
		x"48",	--5983
		x"81",	--5984
		x"4a",	--5985
		x"81",	--5986
		x"58",	--5987
		x"04",	--5988
		x"81",	--5989
		x"68",	--5990
		x"1d",	--5991
		x"50",	--5992
		x"1e",	--5993
		x"52",	--5994
		x"0d",	--5995
		x"0e",	--5996
		x"81",	--5997
		x"6a",	--5998
		x"81",	--5999
		x"6c",	--6000
		x"08",	--6001
		x"18",	--6002
		x"54",	--6003
		x"81",	--6004
		x"6e",	--6005
		x"06",	--6006
		x"55",	--6007
		x"a1",	--6008
		x"58",	--6009
		x"1f",	--6010
		x"6a",	--6011
		x"0f",	--6012
		x"0f",	--6013
		x"04",	--6014
		x"34",	--6015
		x"a0",	--6016
		x"04",	--6017
		x"1b",	--6018
		x"58",	--6019
		x"0b",	--6020
		x"1f",	--6021
		x"6e",	--6022
		x"0f",	--6023
		x"0f",	--6024
		x"1f",	--6025
		x"88",	--6026
		x"0f",	--6027
		x"2e",	--6028
		x"1f",	--6029
		x"02",	--6030
		x"b0",	--6031
		x"b6",	--6032
		x"8b",	--6033
		x"fc",	--6034
		x"8b",	--6035
		x"fe",	--6036
		x"17",	--6037
		x"66",	--6038
		x"1a",	--6039
		x"5c",	--6040
		x"1b",	--6041
		x"5e",	--6042
		x"05",	--6043
		x"08",	--6044
		x"09",	--6045
		x"04",	--6046
		x"14",	--6047
		x"0f",	--6048
		x"0f",	--6049
		x"2c",	--6050
		x"1d",	--6051
		x"02",	--6052
		x"3e",	--6053
		x"3f",	--6054
		x"b0",	--6055
		x"b2",	--6056
		x"0c",	--6057
		x"0d",	--6058
		x"0e",	--6059
		x"0f",	--6060
		x"b0",	--6061
		x"16",	--6062
		x"08",	--6063
		x"09",	--6064
		x"1a",	--6065
		x"0b",	--6066
		x"25",	--6067
		x"81",	--6068
		x"52",	--6069
		x"06",	--6070
		x"1b",	--6071
		x"52",	--6072
		x"e6",	--6073
		x"81",	--6074
		x"50",	--6075
		x"e3",	--6076
		x"1f",	--6077
		x"68",	--6078
		x"0f",	--6079
		x"0f",	--6080
		x"0f",	--6081
		x"1f",	--6082
		x"58",	--6083
		x"8f",	--6084
		x"fc",	--6085
		x"8f",	--6086
		x"fe",	--6087
		x"91",	--6088
		x"48",	--6089
		x"81",	--6090
		x"4a",	--6091
		x"26",	--6092
		x"1e",	--6093
		x"40",	--6094
		x"1f",	--6095
		x"42",	--6096
		x"1e",	--6097
		x"62",	--6098
		x"1f",	--6099
		x"64",	--6100
		x"1f",	--6101
		x"4a",	--6102
		x"06",	--6103
		x"81",	--6104
		x"4a",	--6105
		x"9d",	--6106
		x"1e",	--6107
		x"48",	--6108
		x"9a",	--6109
		x"81",	--6110
		x"40",	--6111
		x"81",	--6112
		x"42",	--6113
		x"30",	--6114
		x"f4",	--6115
		x"81",	--6116
		x"50",	--6117
		x"81",	--6118
		x"52",	--6119
		x"17",	--6120
		x"5c",	--6121
		x"37",	--6122
		x"0d",	--6123
		x"1d",	--6124
		x"1e",	--6125
		x"48",	--6126
		x"1f",	--6127
		x"4a",	--6128
		x"b0",	--6129
		x"a2",	--6130
		x"06",	--6131
		x"07",	--6132
		x"0c",	--6133
		x"3d",	--6134
		x"80",	--6135
		x"b0",	--6136
		x"c6",	--6137
		x"0f",	--6138
		x"2d",	--6139
		x"6b",	--6140
		x"81",	--6141
		x"50",	--6142
		x"81",	--6143
		x"52",	--6144
		x"16",	--6145
		x"40",	--6146
		x"17",	--6147
		x"42",	--6148
		x"36",	--6149
		x"37",	--6150
		x"b1",	--6151
		x"44",	--6152
		x"81",	--6153
		x"46",	--6154
		x"81",	--6155
		x"40",	--6156
		x"81",	--6157
		x"42",	--6158
		x"0d",	--6159
		x"08",	--6160
		x"b1",	--6161
		x"40",	--6162
		x"b1",	--6163
		x"42",	--6164
		x"b1",	--6165
		x"44",	--6166
		x"81",	--6167
		x"46",	--6168
		x"2d",	--6169
		x"0f",	--6170
		x"0f",	--6171
		x"0f",	--6172
		x"39",	--6173
		x"f0",	--6174
		x"09",	--6175
		x"0f",	--6176
		x"0f",	--6177
		x"8f",	--6178
		x"04",	--6179
		x"53",	--6180
		x"8f",	--6181
		x"06",	--6182
		x"e9",	--6183
		x"4f",	--6184
		x"0c",	--6185
		x"3d",	--6186
		x"80",	--6187
		x"0e",	--6188
		x"0f",	--6189
		x"b0",	--6190
		x"b2",	--6191
		x"b0",	--6192
		x"5c",	--6193
		x"b0",	--6194
		x"b6",	--6195
		x"04",	--6196
		x"05",	--6197
		x"1c",	--6198
		x"40",	--6199
		x"0c",	--6200
		x"0c",	--6201
		x"0b",	--6202
		x"0b",	--6203
		x"3b",	--6204
		x"f0",	--6205
		x"0c",	--6206
		x"3d",	--6207
		x"80",	--6208
		x"b0",	--6209
		x"b2",	--6210
		x"0c",	--6211
		x"0d",	--6212
		x"0e",	--6213
		x"0f",	--6214
		x"b0",	--6215
		x"62",	--6216
		x"b0",	--6217
		x"5c",	--6218
		x"8b",	--6219
		x"00",	--6220
		x"8b",	--6221
		x"02",	--6222
		x"91",	--6223
		x"40",	--6224
		x"81",	--6225
		x"42",	--6226
		x"b1",	--6227
		x"44",	--6228
		x"81",	--6229
		x"46",	--6230
		x"1c",	--6231
		x"40",	--6232
		x"0c",	--6233
		x"0c",	--6234
		x"07",	--6235
		x"07",	--6236
		x"37",	--6237
		x"f0",	--6238
		x"0e",	--6239
		x"0f",	--6240
		x"b0",	--6241
		x"5c",	--6242
		x"87",	--6243
		x"00",	--6244
		x"87",	--6245
		x"02",	--6246
		x"10",	--6247
		x"1c",	--6248
		x"40",	--6249
		x"0c",	--6250
		x"0c",	--6251
		x"05",	--6252
		x"05",	--6253
		x"35",	--6254
		x"f0",	--6255
		x"0e",	--6256
		x"0f",	--6257
		x"b0",	--6258
		x"5c",	--6259
		x"85",	--6260
		x"00",	--6261
		x"85",	--6262
		x"02",	--6263
		x"1d",	--6264
		x"44",	--6265
		x"0e",	--6266
		x"3f",	--6267
		x"80",	--6268
		x"b0",	--6269
		x"a2",	--6270
		x"06",	--6271
		x"07",	--6272
		x"14",	--6273
		x"40",	--6274
		x"15",	--6275
		x"42",	--6276
		x"0b",	--6277
		x"05",	--6278
		x"28",	--6279
		x"1f",	--6280
		x"40",	--6281
		x"0f",	--6282
		x"0f",	--6283
		x"0a",	--6284
		x"0a",	--6285
		x"0a",	--6286
		x"3d",	--6287
		x"f0",	--6288
		x"0d",	--6289
		x"0f",	--6290
		x"0f",	--6291
		x"2e",	--6292
		x"1f",	--6293
		x"02",	--6294
		x"b0",	--6295
		x"b6",	--6296
		x"0c",	--6297
		x"0d",	--6298
		x"0e",	--6299
		x"0f",	--6300
		x"b0",	--6301
		x"b2",	--6302
		x"8a",	--6303
		x"00",	--6304
		x"8a",	--6305
		x"02",	--6306
		x"0c",	--6307
		x"3d",	--6308
		x"80",	--6309
		x"0e",	--6310
		x"0f",	--6311
		x"b0",	--6312
		x"b2",	--6313
		x"06",	--6314
		x"07",	--6315
		x"34",	--6316
		x"35",	--6317
		x"2b",	--6318
		x"d6",	--6319
		x"91",	--6320
		x"40",	--6321
		x"44",	--6322
		x"91",	--6323
		x"42",	--6324
		x"46",	--6325
		x"04",	--6326
		x"05",	--6327
		x"07",	--6328
		x"37",	--6329
		x"1f",	--6330
		x"40",	--6331
		x"0f",	--6332
		x"0f",	--6333
		x"0f",	--6334
		x"0f",	--6335
		x"0f",	--6336
		x"2c",	--6337
		x"1d",	--6338
		x"02",	--6339
		x"1e",	--6340
		x"7a",	--6341
		x"1f",	--6342
		x"7c",	--6343
		x"b0",	--6344
		x"b2",	--6345
		x"0c",	--6346
		x"0d",	--6347
		x"0e",	--6348
		x"0f",	--6349
		x"b0",	--6350
		x"16",	--6351
		x"08",	--6352
		x"09",	--6353
		x"1a",	--6354
		x"0b",	--6355
		x"26",	--6356
		x"81",	--6357
		x"4e",	--6358
		x"0a",	--6359
		x"03",	--6360
		x"81",	--6361
		x"4c",	--6362
		x"06",	--6363
		x"05",	--6364
		x"04",	--6365
		x"0b",	--6366
		x"da",	--6367
		x"04",	--6368
		x"d8",	--6369
		x"3f",	--6370
		x"50",	--6371
		x"0f",	--6372
		x"0f",	--6373
		x"8f",	--6374
		x"00",	--6375
		x"8f",	--6376
		x"02",	--6377
		x"b1",	--6378
		x"44",	--6379
		x"b1",	--6380
		x"46",	--6381
		x"27",	--6382
		x"14",	--6383
		x"05",	--6384
		x"81",	--6385
		x"46",	--6386
		x"06",	--6387
		x"06",	--6388
		x"08",	--6389
		x"09",	--6390
		x"0a",	--6391
		x"0b",	--6392
		x"db",	--6393
		x"b1",	--6394
		x"03",	--6395
		x"86",	--6396
		x"08",	--6397
		x"91",	--6398
		x"86",	--6399
		x"3b",	--6400
		x"81",	--6401
		x"86",	--6402
		x"09",	--6403
		x"30",	--6404
		x"5c",	--6405
		x"b1",	--6406
		x"03",	--6407
		x"86",	--6408
		x"02",	--6409
		x"30",	--6410
		x"5c",	--6411
		x"cf",	--6412
		x"16",	--6413
		x"40",	--6414
		x"17",	--6415
		x"42",	--6416
		x"05",	--6417
		x"0a",	--6418
		x"0b",	--6419
		x"07",	--6420
		x"16",	--6421
		x"1f",	--6422
		x"40",	--6423
		x"0f",	--6424
		x"0f",	--6425
		x"3e",	--6426
		x"50",	--6427
		x"0e",	--6428
		x"0f",	--6429
		x"0f",	--6430
		x"2c",	--6431
		x"1d",	--6432
		x"02",	--6433
		x"0e",	--6434
		x"0f",	--6435
		x"b0",	--6436
		x"16",	--6437
		x"0a",	--6438
		x"0b",	--6439
		x"36",	--6440
		x"37",	--6441
		x"25",	--6442
		x"e8",	--6443
		x"81",	--6444
		x"50",	--6445
		x"03",	--6446
		x"81",	--6447
		x"52",	--6448
		x"02",	--6449
		x"3b",	--6450
		x"00",	--6451
		x"18",	--6452
		x"60",	--6453
		x"88",	--6454
		x"00",	--6455
		x"88",	--6456
		x"02",	--6457
		x"30",	--6458
		x"5c",	--6459
		x"16",	--6460
		x"40",	--6461
		x"17",	--6462
		x"42",	--6463
		x"05",	--6464
		x"0a",	--6465
		x"0b",	--6466
		x"07",	--6467
		x"16",	--6468
		x"1f",	--6469
		x"40",	--6470
		x"0f",	--6471
		x"0f",	--6472
		x"39",	--6473
		x"50",	--6474
		x"09",	--6475
		x"0f",	--6476
		x"0f",	--6477
		x"2c",	--6478
		x"1d",	--6479
		x"02",	--6480
		x"0e",	--6481
		x"0f",	--6482
		x"b0",	--6483
		x"16",	--6484
		x"0a",	--6485
		x"0b",	--6486
		x"36",	--6487
		x"37",	--6488
		x"25",	--6489
		x"e8",	--6490
		x"0c",	--6491
		x"0d",	--6492
		x"81",	--6493
		x"50",	--6494
		x"03",	--6495
		x"81",	--6496
		x"52",	--6497
		x"02",	--6498
		x"3b",	--6499
		x"00",	--6500
		x"18",	--6501
		x"60",	--6502
		x"88",	--6503
		x"00",	--6504
		x"88",	--6505
		x"02",	--6506
		x"1e",	--6507
		x"50",	--6508
		x"1f",	--6509
		x"52",	--6510
		x"b0",	--6511
		x"62",	--6512
		x"05",	--6513
		x"35",	--6514
		x"54",	--6515
		x"16",	--6516
		x"07",	--6517
		x"06",	--6518
		x"3c",	--6519
		x"3d",	--6520
		x"b0",	--6521
		x"16",	--6522
		x"16",	--6523
		x"07",	--6524
		x"81",	--6525
		x"42",	--6526
		x"06",	--6527
		x"17",	--6528
		x"42",	--6529
		x"f4",	--6530
		x"81",	--6531
		x"40",	--6532
		x"f1",	--6533
		x"0a",	--6534
		x"0b",	--6535
		x"81",	--6536
		x"50",	--6537
		x"03",	--6538
		x"81",	--6539
		x"52",	--6540
		x"02",	--6541
		x"3b",	--6542
		x"00",	--6543
		x"19",	--6544
		x"60",	--6545
		x"89",	--6546
		x"04",	--6547
		x"89",	--6548
		x"06",	--6549
		x"30",	--6550
		x"5c",	--6551
		x"1f",	--6552
		x"5c",	--6553
		x"0f",	--6554
		x"0f",	--6555
		x"3a",	--6556
		x"50",	--6557
		x"0a",	--6558
		x"0a",	--6559
		x"1a",	--6560
		x"48",	--6561
		x"81",	--6562
		x"44",	--6563
		x"16",	--6564
		x"04",	--6565
		x"17",	--6566
		x"06",	--6567
		x"1f",	--6568
		x"40",	--6569
		x"0f",	--6570
		x"0f",	--6571
		x"39",	--6572
		x"50",	--6573
		x"09",	--6574
		x"09",	--6575
		x"19",	--6576
		x"54",	--6577
		x"81",	--6578
		x"4c",	--6579
		x"28",	--6580
		x"19",	--6581
		x"02",	--6582
		x"0c",	--6583
		x"0d",	--6584
		x"0e",	--6585
		x"0f",	--6586
		x"b0",	--6587
		x"16",	--6588
		x"0a",	--6589
		x"0b",	--6590
		x"0c",	--6591
		x"0d",	--6592
		x"0e",	--6593
		x"0f",	--6594
		x"b0",	--6595
		x"62",	--6596
		x"0c",	--6597
		x"0d",	--6598
		x"0e",	--6599
		x"0f",	--6600
		x"b0",	--6601
		x"16",	--6602
		x"18",	--6603
		x"4c",	--6604
		x"88",	--6605
		x"00",	--6606
		x"88",	--6607
		x"02",	--6608
		x"19",	--6609
		x"44",	--6610
		x"89",	--6611
		x"04",	--6612
		x"89",	--6613
		x"06",	--6614
		x"34",	--6615
		x"35",	--6616
		x"a1",	--6617
		x"54",	--6618
		x"12",	--6619
		x"1c",	--6620
		x"40",	--6621
		x"1d",	--6622
		x"42",	--6623
		x"81",	--6624
		x"54",	--6625
		x"81",	--6626
		x"48",	--6627
		x"08",	--6628
		x"09",	--6629
		x"38",	--6630
		x"39",	--6631
		x"81",	--6632
		x"5c",	--6633
		x"81",	--6634
		x"5e",	--6635
		x"04",	--6636
		x"05",	--6637
		x"a1",	--6638
		x"48",	--6639
		x"05",	--6640
		x"04",	--6641
		x"15",	--6642
		x"a4",	--6643
		x"14",	--6644
		x"a2",	--6645
		x"1c",	--6646
		x"40",	--6647
		x"1d",	--6648
		x"42",	--6649
		x"81",	--6650
		x"54",	--6651
		x"81",	--6652
		x"48",	--6653
		x"09",	--6654
		x"0a",	--6655
		x"39",	--6656
		x"3a",	--6657
		x"81",	--6658
		x"5c",	--6659
		x"81",	--6660
		x"5e",	--6661
		x"04",	--6662
		x"05",	--6663
		x"43",	--6664
		x"1f",	--6665
		x"5c",	--6666
		x"0f",	--6667
		x"0f",	--6668
		x"3a",	--6669
		x"50",	--6670
		x"0a",	--6671
		x"0a",	--6672
		x"1a",	--6673
		x"48",	--6674
		x"81",	--6675
		x"44",	--6676
		x"16",	--6677
		x"04",	--6678
		x"17",	--6679
		x"06",	--6680
		x"1f",	--6681
		x"40",	--6682
		x"0f",	--6683
		x"0f",	--6684
		x"39",	--6685
		x"50",	--6686
		x"09",	--6687
		x"09",	--6688
		x"19",	--6689
		x"54",	--6690
		x"81",	--6691
		x"4c",	--6692
		x"28",	--6693
		x"19",	--6694
		x"02",	--6695
		x"0c",	--6696
		x"0d",	--6697
		x"0e",	--6698
		x"0f",	--6699
		x"b0",	--6700
		x"16",	--6701
		x"0a",	--6702
		x"0b",	--6703
		x"0c",	--6704
		x"0d",	--6705
		x"0e",	--6706
		x"0f",	--6707
		x"b0",	--6708
		x"62",	--6709
		x"0c",	--6710
		x"0d",	--6711
		x"0e",	--6712
		x"0f",	--6713
		x"b0",	--6714
		x"16",	--6715
		x"18",	--6716
		x"4c",	--6717
		x"88",	--6718
		x"00",	--6719
		x"88",	--6720
		x"02",	--6721
		x"19",	--6722
		x"44",	--6723
		x"89",	--6724
		x"04",	--6725
		x"89",	--6726
		x"06",	--6727
		x"34",	--6728
		x"35",	--6729
		x"a1",	--6730
		x"54",	--6731
		x"a1",	--6732
		x"48",	--6733
		x"05",	--6734
		x"04",	--6735
		x"15",	--6736
		x"b7",	--6737
		x"24",	--6738
		x"b5",	--6739
		x"16",	--6740
		x"40",	--6741
		x"17",	--6742
		x"42",	--6743
		x"05",	--6744
		x"0a",	--6745
		x"0b",	--6746
		x"15",	--6747
		x"1f",	--6748
		x"40",	--6749
		x"0f",	--6750
		x"0f",	--6751
		x"3d",	--6752
		x"50",	--6753
		x"0d",	--6754
		x"0f",	--6755
		x"0f",	--6756
		x"2c",	--6757
		x"1d",	--6758
		x"02",	--6759
		x"0e",	--6760
		x"0f",	--6761
		x"b0",	--6762
		x"16",	--6763
		x"0a",	--6764
		x"0b",	--6765
		x"36",	--6766
		x"37",	--6767
		x"25",	--6768
		x"07",	--6769
		x"04",	--6770
		x"17",	--6771
		x"e7",	--6772
		x"26",	--6773
		x"e5",	--6774
		x"81",	--6775
		x"50",	--6776
		x"16",	--6777
		x"81",	--6778
		x"52",	--6779
		x"13",	--6780
		x"18",	--6781
		x"60",	--6782
		x"98",	--6783
		x"50",	--6784
		x"00",	--6785
		x"98",	--6786
		x"52",	--6787
		x"02",	--6788
		x"98",	--6789
		x"54",	--6790
		x"04",	--6791
		x"98",	--6792
		x"56",	--6793
		x"06",	--6794
		x"88",	--6795
		x"08",	--6796
		x"88",	--6797
		x"0a",	--6798
		x"1e",	--6799
		x"1d",	--6800
		x"50",	--6801
		x"1e",	--6802
		x"52",	--6803
		x"3e",	--6804
		x"00",	--6805
		x"18",	--6806
		x"60",	--6807
		x"88",	--6808
		x"00",	--6809
		x"88",	--6810
		x"02",	--6811
		x"1d",	--6812
		x"54",	--6813
		x"1e",	--6814
		x"56",	--6815
		x"3e",	--6816
		x"00",	--6817
		x"88",	--6818
		x"04",	--6819
		x"88",	--6820
		x"06",	--6821
		x"0d",	--6822
		x"0e",	--6823
		x"3e",	--6824
		x"00",	--6825
		x"88",	--6826
		x"08",	--6827
		x"88",	--6828
		x"0a",	--6829
		x"1f",	--6830
		x"58",	--6831
		x"3f",	--6832
		x"07",	--6833
		x"31",	--6834
		x"74",	--6835
		x"34",	--6836
		x"35",	--6837
		x"36",	--6838
		x"37",	--6839
		x"38",	--6840
		x"39",	--6841
		x"3a",	--6842
		x"3b",	--6843
		x"30",	--6844
		x"0b",	--6845
		x"0a",	--6846
		x"31",	--6847
		x"0c",	--6848
		x"0d",	--6849
		x"3c",	--6850
		x"3d",	--6851
		x"ff",	--6852
		x"3d",	--6853
		x"49",	--6854
		x"06",	--6855
		x"3d",	--6856
		x"4a",	--6857
		x"06",	--6858
		x"3c",	--6859
		x"d9",	--6860
		x"03",	--6861
		x"0c",	--6862
		x"0d",	--6863
		x"26",	--6864
		x"3d",	--6865
		x"80",	--6866
		x"05",	--6867
		x"0c",	--6868
		x"0d",	--6869
		x"b0",	--6870
		x"62",	--6871
		x"2f",	--6872
		x"0d",	--6873
		x"b0",	--6874
		x"28",	--6875
		x"0a",	--6876
		x"0b",	--6877
		x"3a",	--6878
		x"03",	--6879
		x"0b",	--6880
		x"1c",	--6881
		x"04",	--6882
		x"1d",	--6883
		x"06",	--6884
		x"2e",	--6885
		x"1f",	--6886
		x"02",	--6887
		x"1a",	--6888
		x"02",	--6889
		x"0b",	--6890
		x"0e",	--6891
		x"2a",	--6892
		x"02",	--6893
		x"0b",	--6894
		x"0f",	--6895
		x"2e",	--6896
		x"1f",	--6897
		x"02",	--6898
		x"0a",	--6899
		x"0f",	--6900
		x"0b",	--6901
		x"0d",	--6902
		x"b0",	--6903
		x"44",	--6904
		x"0e",	--6905
		x"13",	--6906
		x"b0",	--6907
		x"1e",	--6908
		x"21",	--6909
		x"02",	--6910
		x"b0",	--6911
		x"44",	--6912
		x"3f",	--6913
		x"00",	--6914
		x"04",	--6915
		x"13",	--6916
		x"b0",	--6917
		x"1e",	--6918
		x"21",	--6919
		x"31",	--6920
		x"3a",	--6921
		x"3b",	--6922
		x"30",	--6923
		x"b0",	--6924
		x"7a",	--6925
		x"30",	--6926
		x"0b",	--6927
		x"0a",	--6928
		x"09",	--6929
		x"08",	--6930
		x"07",	--6931
		x"06",	--6932
		x"05",	--6933
		x"04",	--6934
		x"31",	--6935
		x"08",	--6936
		x"09",	--6937
		x"81",	--6938
		x"00",	--6939
		x"81",	--6940
		x"02",	--6941
		x"0a",	--6942
		x"0b",	--6943
		x"3a",	--6944
		x"3b",	--6945
		x"ff",	--6946
		x"3b",	--6947
		x"00",	--6948
		x"04",	--6949
		x"b0",	--6950
		x"5c",	--6951
		x"0e",	--6952
		x"9b",	--6953
		x"0c",	--6954
		x"0d",	--6955
		x"0e",	--6956
		x"0f",	--6957
		x"b0",	--6958
		x"b2",	--6959
		x"0a",	--6960
		x"0b",	--6961
		x"0c",	--6962
		x"0d",	--6963
		x"b0",	--6964
		x"b2",	--6965
		x"06",	--6966
		x"07",	--6967
		x"3c",	--6968
		x"d3",	--6969
		x"3d",	--6970
		x"2e",	--6971
		x"0e",	--6972
		x"0f",	--6973
		x"b0",	--6974
		x"b2",	--6975
		x"3c",	--6976
		x"34",	--6977
		x"3d",	--6978
		x"d7",	--6979
		x"b0",	--6980
		x"62",	--6981
		x"0c",	--6982
		x"0d",	--6983
		x"0e",	--6984
		x"0f",	--6985
		x"b0",	--6986
		x"b2",	--6987
		x"3c",	--6988
		x"1b",	--6989
		x"3d",	--6990
		x"38",	--6991
		x"b0",	--6992
		x"16",	--6993
		x"0c",	--6994
		x"0d",	--6995
		x"0e",	--6996
		x"0f",	--6997
		x"b0",	--6998
		x"b2",	--6999
		x"3c",	--7000
		x"01",	--7001
		x"3d",	--7002
		x"50",	--7003
		x"b0",	--7004
		x"62",	--7005
		x"0c",	--7006
		x"0d",	--7007
		x"0e",	--7008
		x"0f",	--7009
		x"b0",	--7010
		x"b2",	--7011
		x"3c",	--7012
		x"89",	--7013
		x"3d",	--7014
		x"08",	--7015
		x"b0",	--7016
		x"16",	--7017
		x"04",	--7018
		x"05",	--7019
		x"81",	--7020
		x"1a",	--7021
		x"19",	--7022
		x"0c",	--7023
		x"0d",	--7024
		x"0e",	--7025
		x"0f",	--7026
		x"b0",	--7027
		x"b2",	--7028
		x"3c",	--7029
		x"ab",	--7030
		x"3d",	--7031
		x"2a",	--7032
		x"b0",	--7033
		x"62",	--7034
		x"0c",	--7035
		x"0d",	--7036
		x"0e",	--7037
		x"0f",	--7038
		x"b0",	--7039
		x"b2",	--7040
		x"0c",	--7041
		x"0d",	--7042
		x"0e",	--7043
		x"0f",	--7044
		x"b0",	--7045
		x"16",	--7046
		x"3b",	--7047
		x"0c",	--7048
		x"3d",	--7049
		x"00",	--7050
		x"2e",	--7051
		x"1f",	--7052
		x"02",	--7053
		x"b0",	--7054
		x"b2",	--7055
		x"81",	--7056
		x"04",	--7057
		x"81",	--7058
		x"06",	--7059
		x"0c",	--7060
		x"0d",	--7061
		x"0e",	--7062
		x"0f",	--7063
		x"b0",	--7064
		x"b2",	--7065
		x"0c",	--7066
		x"0d",	--7067
		x"1e",	--7068
		x"04",	--7069
		x"1f",	--7070
		x"06",	--7071
		x"b0",	--7072
		x"62",	--7073
		x"0c",	--7074
		x"0d",	--7075
		x"0e",	--7076
		x"0f",	--7077
		x"b0",	--7078
		x"b2",	--7079
		x"2c",	--7080
		x"1d",	--7081
		x"02",	--7082
		x"b0",	--7083
		x"62",	--7084
		x"0a",	--7085
		x"0b",	--7086
		x"3c",	--7087
		x"ab",	--7088
		x"3d",	--7089
		x"2a",	--7090
		x"0e",	--7091
		x"0f",	--7092
		x"b0",	--7093
		x"b2",	--7094
		x"0c",	--7095
		x"0d",	--7096
		x"0e",	--7097
		x"0f",	--7098
		x"b0",	--7099
		x"16",	--7100
		x"0c",	--7101
		x"0d",	--7102
		x"0e",	--7103
		x"0f",	--7104
		x"b0",	--7105
		x"62",	--7106
		x"08",	--7107
		x"09",	--7108
		x"0e",	--7109
		x"0f",	--7110
		x"31",	--7111
		x"34",	--7112
		x"35",	--7113
		x"36",	--7114
		x"37",	--7115
		x"38",	--7116
		x"39",	--7117
		x"3a",	--7118
		x"3b",	--7119
		x"30",	--7120
		x"0b",	--7121
		x"0a",	--7122
		x"09",	--7123
		x"08",	--7124
		x"07",	--7125
		x"07",	--7126
		x"08",	--7127
		x"09",	--7128
		x"0c",	--7129
		x"0d",	--7130
		x"3c",	--7131
		x"3d",	--7132
		x"ff",	--7133
		x"0c",	--7134
		x"02",	--7135
		x"0d",	--7136
		x"a8",	--7137
		x"3d",	--7138
		x"80",	--7139
		x"05",	--7140
		x"0c",	--7141
		x"0d",	--7142
		x"b0",	--7143
		x"16",	--7144
		x"a0",	--7145
		x"3d",	--7146
		x"80",	--7147
		x"0a",	--7148
		x"0c",	--7149
		x"0d",	--7150
		x"7e",	--7151
		x"07",	--7152
		x"12",	--7153
		x"0d",	--7154
		x"0c",	--7155
		x"7e",	--7156
		x"fb",	--7157
		x"1b",	--7158
		x"0c",	--7159
		x"3d",	--7160
		x"00",	--7161
		x"b0",	--7162
		x"b2",	--7163
		x"08",	--7164
		x"09",	--7165
		x"0a",	--7166
		x"0b",	--7167
		x"0a",	--7168
		x"3b",	--7169
		x"80",	--7170
		x"0c",	--7171
		x"0d",	--7172
		x"8d",	--7173
		x"8d",	--7174
		x"8d",	--7175
		x"8d",	--7176
		x"7e",	--7177
		x"07",	--7178
		x"0d",	--7179
		x"0c",	--7180
		x"7e",	--7181
		x"fc",	--7182
		x"3c",	--7183
		x"e7",	--7184
		x"3d",	--7185
		x"0a",	--7186
		x"0e",	--7187
		x"8e",	--7188
		x"8e",	--7189
		x"8e",	--7190
		x"8e",	--7191
		x"0b",	--7192
		x"0c",	--7193
		x"0d",	--7194
		x"0d",	--7195
		x"15",	--7196
		x"03",	--7197
		x"3c",	--7198
		x"ff",	--7199
		x"11",	--7200
		x"3a",	--7201
		x"ca",	--7202
		x"3b",	--7203
		x"49",	--7204
		x"0f",	--7205
		x"04",	--7206
		x"3a",	--7207
		x"ca",	--7208
		x"3b",	--7209
		x"49",	--7210
		x"3c",	--7211
		x"ca",	--7212
		x"3d",	--7213
		x"49",	--7214
		x"0e",	--7215
		x"0f",	--7216
		x"56",	--7217
		x"0d",	--7218
		x"14",	--7219
		x"02",	--7220
		x"1c",	--7221
		x"11",	--7222
		x"0a",	--7223
		x"0b",	--7224
		x"0b",	--7225
		x"7f",	--7226
		x"07",	--7227
		x"0a",	--7228
		x"0b",	--7229
		x"7f",	--7230
		x"fc",	--7231
		x"38",	--7232
		x"39",	--7233
		x"7f",	--7234
		x"08",	--7235
		x"09",	--7236
		x"0e",	--7237
		x"0f",	--7238
		x"42",	--7239
		x"3d",	--7240
		x"05",	--7241
		x"0d",	--7242
		x"27",	--7243
		x"3c",	--7244
		x"ea",	--7245
		x"24",	--7246
		x"0d",	--7247
		x"3d",	--7248
		x"00",	--7249
		x"37",	--7250
		x"31",	--7251
		x"0f",	--7252
		x"3e",	--7253
		x"ca",	--7254
		x"3f",	--7255
		x"49",	--7256
		x"0d",	--7257
		x"04",	--7258
		x"3e",	--7259
		x"ca",	--7260
		x"3f",	--7261
		x"49",	--7262
		x"3c",	--7263
		x"ca",	--7264
		x"3d",	--7265
		x"49",	--7266
		x"24",	--7267
		x"3e",	--7268
		x"60",	--7269
		x"3f",	--7270
		x"a2",	--7271
		x"0d",	--7272
		x"04",	--7273
		x"3e",	--7274
		x"60",	--7275
		x"3f",	--7276
		x"a2",	--7277
		x"3c",	--7278
		x"60",	--7279
		x"3d",	--7280
		x"a2",	--7281
		x"15",	--7282
		x"0a",	--7283
		x"0b",	--7284
		x"0b",	--7285
		x"3b",	--7286
		x"19",	--7287
		x"7f",	--7288
		x"07",	--7289
		x"0a",	--7290
		x"0b",	--7291
		x"7f",	--7292
		x"fc",	--7293
		x"0e",	--7294
		x"0f",	--7295
		x"3e",	--7296
		x"3f",	--7297
		x"7f",	--7298
		x"0e",	--7299
		x"0f",	--7300
		x"0c",	--7301
		x"3d",	--7302
		x"00",	--7303
		x"b0",	--7304
		x"b2",	--7305
		x"37",	--7306
		x"38",	--7307
		x"39",	--7308
		x"3a",	--7309
		x"3b",	--7310
		x"30",	--7311
		x"b0",	--7312
		x"a2",	--7313
		x"30",	--7314
		x"0b",	--7315
		x"0a",	--7316
		x"09",	--7317
		x"08",	--7318
		x"07",	--7319
		x"06",	--7320
		x"05",	--7321
		x"04",	--7322
		x"21",	--7323
		x"06",	--7324
		x"07",	--7325
		x"08",	--7326
		x"09",	--7327
		x"38",	--7328
		x"39",	--7329
		x"ff",	--7330
		x"0c",	--7331
		x"0d",	--7332
		x"7a",	--7333
		x"07",	--7334
		x"12",	--7335
		x"0d",	--7336
		x"0c",	--7337
		x"7a",	--7338
		x"fb",	--7339
		x"3c",	--7340
		x"81",	--7341
		x"3d",	--7342
		x"0d",	--7343
		x"05",	--7344
		x"1d",	--7345
		x"57",	--7346
		x"3c",	--7347
		x"17",	--7348
		x"54",	--7349
		x"0a",	--7350
		x"0b",	--7351
		x"0d",	--7352
		x"09",	--7353
		x"81",	--7354
		x"00",	--7355
		x"38",	--7356
		x"39",	--7357
		x"7f",	--7358
		x"6d",	--7359
		x"7d",	--7360
		x"1f",	--7361
		x"1d",	--7362
		x"3c",	--7363
		x"ca",	--7364
		x"3d",	--7365
		x"49",	--7366
		x"b0",	--7367
		x"16",	--7368
		x"0c",	--7369
		x"0d",	--7370
		x"b0",	--7371
		x"76",	--7372
		x"0f",	--7373
		x"43",	--7374
		x"42",	--7375
		x"0b",	--7376
		x"03",	--7377
		x"0a",	--7378
		x"0b",	--7379
		x"3d",	--7380
		x"08",	--7381
		x"02",	--7382
		x"09",	--7383
		x"39",	--7384
		x"0a",	--7385
		x"3b",	--7386
		x"80",	--7387
		x"35",	--7388
		x"09",	--7389
		x"08",	--7390
		x"7d",	--7391
		x"4d",	--7392
		x"fb",	--7393
		x"04",	--7394
		x"05",	--7395
		x"04",	--7396
		x"05",	--7397
		x"04",	--7398
		x"02",	--7399
		x"05",	--7400
		x"2a",	--7401
		x"3c",	--7402
		x"ca",	--7403
		x"3d",	--7404
		x"49",	--7405
		x"b0",	--7406
		x"16",	--7407
		x"0c",	--7408
		x"0d",	--7409
		x"b0",	--7410
		x"76",	--7411
		x"0f",	--7412
		x"1c",	--7413
		x"1b",	--7414
		x"07",	--7415
		x"0e",	--7416
		x"0a",	--7417
		x"3b",	--7418
		x"80",	--7419
		x"6c",	--7420
		x"7c",	--7421
		x"1f",	--7422
		x"4c",	--7423
		x"04",	--7424
		x"0b",	--7425
		x"0a",	--7426
		x"7c",	--7427
		x"fa",	--7428
		x"0a",	--7429
		x"0b",	--7430
		x"0a",	--7431
		x"0b",	--7432
		x"08",	--7433
		x"39",	--7434
		x"80",	--7435
		x"07",	--7436
		x"0c",	--7437
		x"0d",	--7438
		x"b0",	--7439
		x"16",	--7440
		x"02",	--7441
		x"0e",	--7442
		x"0f",	--7443
		x"21",	--7444
		x"34",	--7445
		x"35",	--7446
		x"36",	--7447
		x"37",	--7448
		x"38",	--7449
		x"39",	--7450
		x"3a",	--7451
		x"3b",	--7452
		x"30",	--7453
		x"b0",	--7454
		x"26",	--7455
		x"30",	--7456
		x"0b",	--7457
		x"0a",	--7458
		x"0a",	--7459
		x"0b",	--7460
		x"0c",	--7461
		x"3d",	--7462
		x"00",	--7463
		x"b0",	--7464
		x"c6",	--7465
		x"0f",	--7466
		x"07",	--7467
		x"0e",	--7468
		x"0f",	--7469
		x"b0",	--7470
		x"5c",	--7471
		x"3a",	--7472
		x"3b",	--7473
		x"30",	--7474
		x"0c",	--7475
		x"3d",	--7476
		x"00",	--7477
		x"0e",	--7478
		x"0f",	--7479
		x"b0",	--7480
		x"62",	--7481
		x"b0",	--7482
		x"5c",	--7483
		x"0e",	--7484
		x"3f",	--7485
		x"00",	--7486
		x"3a",	--7487
		x"3b",	--7488
		x"30",	--7489
		x"0b",	--7490
		x"0a",	--7491
		x"09",	--7492
		x"08",	--7493
		x"07",	--7494
		x"06",	--7495
		x"05",	--7496
		x"04",	--7497
		x"31",	--7498
		x"fa",	--7499
		x"08",	--7500
		x"6b",	--7501
		x"6b",	--7502
		x"67",	--7503
		x"6c",	--7504
		x"6c",	--7505
		x"e9",	--7506
		x"6b",	--7507
		x"02",	--7508
		x"30",	--7509
		x"04",	--7510
		x"6c",	--7511
		x"e3",	--7512
		x"6c",	--7513
		x"bb",	--7514
		x"6b",	--7515
		x"df",	--7516
		x"91",	--7517
		x"02",	--7518
		x"00",	--7519
		x"1b",	--7520
		x"02",	--7521
		x"14",	--7522
		x"04",	--7523
		x"15",	--7524
		x"06",	--7525
		x"16",	--7526
		x"04",	--7527
		x"17",	--7528
		x"06",	--7529
		x"2c",	--7530
		x"0c",	--7531
		x"09",	--7532
		x"0c",	--7533
		x"bf",	--7534
		x"39",	--7535
		x"20",	--7536
		x"50",	--7537
		x"1c",	--7538
		x"d7",	--7539
		x"81",	--7540
		x"02",	--7541
		x"81",	--7542
		x"04",	--7543
		x"4c",	--7544
		x"7c",	--7545
		x"1f",	--7546
		x"0b",	--7547
		x"0a",	--7548
		x"0b",	--7549
		x"12",	--7550
		x"0b",	--7551
		x"0a",	--7552
		x"7c",	--7553
		x"fb",	--7554
		x"81",	--7555
		x"02",	--7556
		x"81",	--7557
		x"04",	--7558
		x"1c",	--7559
		x"0d",	--7560
		x"79",	--7561
		x"1f",	--7562
		x"04",	--7563
		x"0c",	--7564
		x"0d",	--7565
		x"79",	--7566
		x"fc",	--7567
		x"3c",	--7568
		x"3d",	--7569
		x"0c",	--7570
		x"0d",	--7571
		x"1a",	--7572
		x"0b",	--7573
		x"0c",	--7574
		x"02",	--7575
		x"0d",	--7576
		x"e5",	--7577
		x"16",	--7578
		x"02",	--7579
		x"17",	--7580
		x"04",	--7581
		x"06",	--7582
		x"07",	--7583
		x"5f",	--7584
		x"01",	--7585
		x"5f",	--7586
		x"01",	--7587
		x"28",	--7588
		x"c8",	--7589
		x"01",	--7590
		x"a8",	--7591
		x"02",	--7592
		x"0e",	--7593
		x"0f",	--7594
		x"0e",	--7595
		x"0f",	--7596
		x"88",	--7597
		x"04",	--7598
		x"88",	--7599
		x"06",	--7600
		x"f8",	--7601
		x"03",	--7602
		x"00",	--7603
		x"0f",	--7604
		x"4d",	--7605
		x"0f",	--7606
		x"31",	--7607
		x"06",	--7608
		x"34",	--7609
		x"35",	--7610
		x"36",	--7611
		x"37",	--7612
		x"38",	--7613
		x"39",	--7614
		x"3a",	--7615
		x"3b",	--7616
		x"30",	--7617
		x"2b",	--7618
		x"67",	--7619
		x"81",	--7620
		x"00",	--7621
		x"04",	--7622
		x"05",	--7623
		x"5f",	--7624
		x"01",	--7625
		x"5f",	--7626
		x"01",	--7627
		x"d8",	--7628
		x"4f",	--7629
		x"68",	--7630
		x"0e",	--7631
		x"0f",	--7632
		x"0e",	--7633
		x"0f",	--7634
		x"0f",	--7635
		x"69",	--7636
		x"c8",	--7637
		x"01",	--7638
		x"a8",	--7639
		x"02",	--7640
		x"88",	--7641
		x"04",	--7642
		x"88",	--7643
		x"06",	--7644
		x"0c",	--7645
		x"0d",	--7646
		x"3c",	--7647
		x"3d",	--7648
		x"3d",	--7649
		x"ff",	--7650
		x"05",	--7651
		x"3d",	--7652
		x"00",	--7653
		x"17",	--7654
		x"3c",	--7655
		x"15",	--7656
		x"1b",	--7657
		x"02",	--7658
		x"3b",	--7659
		x"0e",	--7660
		x"0f",	--7661
		x"0a",	--7662
		x"3b",	--7663
		x"0c",	--7664
		x"0d",	--7665
		x"3c",	--7666
		x"3d",	--7667
		x"3d",	--7668
		x"ff",	--7669
		x"f5",	--7670
		x"3c",	--7671
		x"88",	--7672
		x"04",	--7673
		x"88",	--7674
		x"06",	--7675
		x"88",	--7676
		x"02",	--7677
		x"f8",	--7678
		x"03",	--7679
		x"00",	--7680
		x"0f",	--7681
		x"b3",	--7682
		x"0c",	--7683
		x"0d",	--7684
		x"1c",	--7685
		x"0d",	--7686
		x"12",	--7687
		x"0f",	--7688
		x"0e",	--7689
		x"0a",	--7690
		x"0b",	--7691
		x"0a",	--7692
		x"0b",	--7693
		x"88",	--7694
		x"04",	--7695
		x"88",	--7696
		x"06",	--7697
		x"98",	--7698
		x"02",	--7699
		x"0f",	--7700
		x"a1",	--7701
		x"6b",	--7702
		x"9f",	--7703
		x"ad",	--7704
		x"00",	--7705
		x"9d",	--7706
		x"02",	--7707
		x"02",	--7708
		x"9d",	--7709
		x"04",	--7710
		x"04",	--7711
		x"9d",	--7712
		x"06",	--7713
		x"06",	--7714
		x"5e",	--7715
		x"01",	--7716
		x"5e",	--7717
		x"01",	--7718
		x"cd",	--7719
		x"01",	--7720
		x"0f",	--7721
		x"8c",	--7722
		x"06",	--7723
		x"07",	--7724
		x"9a",	--7725
		x"39",	--7726
		x"19",	--7727
		x"39",	--7728
		x"20",	--7729
		x"8f",	--7730
		x"3e",	--7731
		x"3c",	--7732
		x"b6",	--7733
		x"c1",	--7734
		x"0e",	--7735
		x"0f",	--7736
		x"0e",	--7737
		x"0f",	--7738
		x"97",	--7739
		x"0f",	--7740
		x"79",	--7741
		x"d8",	--7742
		x"01",	--7743
		x"a8",	--7744
		x"02",	--7745
		x"3e",	--7746
		x"3f",	--7747
		x"1e",	--7748
		x"0f",	--7749
		x"88",	--7750
		x"04",	--7751
		x"88",	--7752
		x"06",	--7753
		x"92",	--7754
		x"0c",	--7755
		x"7b",	--7756
		x"81",	--7757
		x"00",	--7758
		x"81",	--7759
		x"02",	--7760
		x"81",	--7761
		x"04",	--7762
		x"4d",	--7763
		x"7d",	--7764
		x"1f",	--7765
		x"0c",	--7766
		x"4b",	--7767
		x"0c",	--7768
		x"0d",	--7769
		x"12",	--7770
		x"0d",	--7771
		x"0c",	--7772
		x"7b",	--7773
		x"fb",	--7774
		x"81",	--7775
		x"02",	--7776
		x"81",	--7777
		x"04",	--7778
		x"1c",	--7779
		x"0d",	--7780
		x"79",	--7781
		x"1f",	--7782
		x"04",	--7783
		x"0c",	--7784
		x"0d",	--7785
		x"79",	--7786
		x"fc",	--7787
		x"3c",	--7788
		x"3d",	--7789
		x"0c",	--7790
		x"0d",	--7791
		x"1a",	--7792
		x"0b",	--7793
		x"0c",	--7794
		x"04",	--7795
		x"0d",	--7796
		x"02",	--7797
		x"0a",	--7798
		x"0b",	--7799
		x"14",	--7800
		x"02",	--7801
		x"15",	--7802
		x"04",	--7803
		x"04",	--7804
		x"05",	--7805
		x"49",	--7806
		x"0a",	--7807
		x"0b",	--7808
		x"18",	--7809
		x"6c",	--7810
		x"33",	--7811
		x"df",	--7812
		x"01",	--7813
		x"01",	--7814
		x"2f",	--7815
		x"3f",	--7816
		x"a6",	--7817
		x"2c",	--7818
		x"31",	--7819
		x"e0",	--7820
		x"81",	--7821
		x"04",	--7822
		x"81",	--7823
		x"06",	--7824
		x"81",	--7825
		x"00",	--7826
		x"81",	--7827
		x"02",	--7828
		x"0e",	--7829
		x"3e",	--7830
		x"18",	--7831
		x"0f",	--7832
		x"2f",	--7833
		x"b0",	--7834
		x"1e",	--7835
		x"0e",	--7836
		x"3e",	--7837
		x"10",	--7838
		x"0f",	--7839
		x"b0",	--7840
		x"1e",	--7841
		x"0d",	--7842
		x"3d",	--7843
		x"0e",	--7844
		x"3e",	--7845
		x"10",	--7846
		x"0f",	--7847
		x"3f",	--7848
		x"18",	--7849
		x"b0",	--7850
		x"84",	--7851
		x"b0",	--7852
		x"40",	--7853
		x"31",	--7854
		x"20",	--7855
		x"30",	--7856
		x"31",	--7857
		x"e0",	--7858
		x"81",	--7859
		x"04",	--7860
		x"81",	--7861
		x"06",	--7862
		x"81",	--7863
		x"00",	--7864
		x"81",	--7865
		x"02",	--7866
		x"0e",	--7867
		x"3e",	--7868
		x"18",	--7869
		x"0f",	--7870
		x"2f",	--7871
		x"b0",	--7872
		x"1e",	--7873
		x"0e",	--7874
		x"3e",	--7875
		x"10",	--7876
		x"0f",	--7877
		x"b0",	--7878
		x"1e",	--7879
		x"d1",	--7880
		x"11",	--7881
		x"0d",	--7882
		x"3d",	--7883
		x"0e",	--7884
		x"3e",	--7885
		x"10",	--7886
		x"0f",	--7887
		x"3f",	--7888
		x"18",	--7889
		x"b0",	--7890
		x"84",	--7891
		x"b0",	--7892
		x"40",	--7893
		x"31",	--7894
		x"20",	--7895
		x"30",	--7896
		x"0b",	--7897
		x"0a",	--7898
		x"09",	--7899
		x"08",	--7900
		x"07",	--7901
		x"06",	--7902
		x"05",	--7903
		x"04",	--7904
		x"31",	--7905
		x"dc",	--7906
		x"81",	--7907
		x"04",	--7908
		x"81",	--7909
		x"06",	--7910
		x"81",	--7911
		x"00",	--7912
		x"81",	--7913
		x"02",	--7914
		x"0e",	--7915
		x"3e",	--7916
		x"18",	--7917
		x"0f",	--7918
		x"2f",	--7919
		x"b0",	--7920
		x"1e",	--7921
		x"0e",	--7922
		x"3e",	--7923
		x"10",	--7924
		x"0f",	--7925
		x"b0",	--7926
		x"1e",	--7927
		x"5f",	--7928
		x"18",	--7929
		x"6f",	--7930
		x"b6",	--7931
		x"5e",	--7932
		x"10",	--7933
		x"6e",	--7934
		x"d9",	--7935
		x"6f",	--7936
		x"ae",	--7937
		x"6e",	--7938
		x"e2",	--7939
		x"6f",	--7940
		x"ac",	--7941
		x"6e",	--7942
		x"d1",	--7943
		x"14",	--7944
		x"1c",	--7945
		x"15",	--7946
		x"1e",	--7947
		x"18",	--7948
		x"14",	--7949
		x"19",	--7950
		x"16",	--7951
		x"3c",	--7952
		x"20",	--7953
		x"0e",	--7954
		x"0f",	--7955
		x"06",	--7956
		x"07",	--7957
		x"81",	--7958
		x"20",	--7959
		x"81",	--7960
		x"22",	--7961
		x"0a",	--7962
		x"0b",	--7963
		x"81",	--7964
		x"20",	--7965
		x"08",	--7966
		x"08",	--7967
		x"09",	--7968
		x"12",	--7969
		x"05",	--7970
		x"04",	--7971
		x"b1",	--7972
		x"20",	--7973
		x"19",	--7974
		x"14",	--7975
		x"0d",	--7976
		x"0a",	--7977
		x"0b",	--7978
		x"0e",	--7979
		x"0f",	--7980
		x"1c",	--7981
		x"0d",	--7982
		x"0b",	--7983
		x"03",	--7984
		x"0b",	--7985
		x"0c",	--7986
		x"0d",	--7987
		x"0e",	--7988
		x"0f",	--7989
		x"06",	--7990
		x"07",	--7991
		x"09",	--7992
		x"e5",	--7993
		x"16",	--7994
		x"07",	--7995
		x"e2",	--7996
		x"0a",	--7997
		x"f5",	--7998
		x"f2",	--7999
		x"81",	--8000
		x"20",	--8001
		x"81",	--8002
		x"22",	--8003
		x"0c",	--8004
		x"1a",	--8005
		x"1a",	--8006
		x"1a",	--8007
		x"12",	--8008
		x"06",	--8009
		x"26",	--8010
		x"81",	--8011
		x"0a",	--8012
		x"5d",	--8013
		x"d1",	--8014
		x"11",	--8015
		x"19",	--8016
		x"83",	--8017
		x"c1",	--8018
		x"09",	--8019
		x"0c",	--8020
		x"3c",	--8021
		x"3f",	--8022
		x"00",	--8023
		x"18",	--8024
		x"1d",	--8025
		x"0a",	--8026
		x"3d",	--8027
		x"1a",	--8028
		x"20",	--8029
		x"1b",	--8030
		x"22",	--8031
		x"0c",	--8032
		x"0e",	--8033
		x"0f",	--8034
		x"0b",	--8035
		x"2a",	--8036
		x"0a",	--8037
		x"0b",	--8038
		x"3d",	--8039
		x"3f",	--8040
		x"00",	--8041
		x"f5",	--8042
		x"81",	--8043
		x"20",	--8044
		x"81",	--8045
		x"22",	--8046
		x"81",	--8047
		x"0a",	--8048
		x"0c",	--8049
		x"0d",	--8050
		x"3c",	--8051
		x"7f",	--8052
		x"0d",	--8053
		x"3c",	--8054
		x"40",	--8055
		x"44",	--8056
		x"81",	--8057
		x"0c",	--8058
		x"81",	--8059
		x"0e",	--8060
		x"f1",	--8061
		x"03",	--8062
		x"08",	--8063
		x"0f",	--8064
		x"3f",	--8065
		x"b0",	--8066
		x"40",	--8067
		x"31",	--8068
		x"24",	--8069
		x"34",	--8070
		x"35",	--8071
		x"36",	--8072
		x"37",	--8073
		x"38",	--8074
		x"39",	--8075
		x"3a",	--8076
		x"3b",	--8077
		x"30",	--8078
		x"1e",	--8079
		x"0f",	--8080
		x"d3",	--8081
		x"3a",	--8082
		x"03",	--8083
		x"08",	--8084
		x"1e",	--8085
		x"10",	--8086
		x"1c",	--8087
		x"20",	--8088
		x"1d",	--8089
		x"22",	--8090
		x"12",	--8091
		x"0d",	--8092
		x"0c",	--8093
		x"06",	--8094
		x"07",	--8095
		x"06",	--8096
		x"37",	--8097
		x"00",	--8098
		x"81",	--8099
		x"20",	--8100
		x"81",	--8101
		x"22",	--8102
		x"12",	--8103
		x"0f",	--8104
		x"0e",	--8105
		x"1a",	--8106
		x"0f",	--8107
		x"e7",	--8108
		x"81",	--8109
		x"0a",	--8110
		x"a6",	--8111
		x"6e",	--8112
		x"36",	--8113
		x"5f",	--8114
		x"d1",	--8115
		x"11",	--8116
		x"19",	--8117
		x"20",	--8118
		x"c1",	--8119
		x"19",	--8120
		x"0f",	--8121
		x"3f",	--8122
		x"18",	--8123
		x"c5",	--8124
		x"0d",	--8125
		x"ba",	--8126
		x"0c",	--8127
		x"0d",	--8128
		x"3c",	--8129
		x"80",	--8130
		x"0d",	--8131
		x"0c",	--8132
		x"b3",	--8133
		x"0d",	--8134
		x"b1",	--8135
		x"81",	--8136
		x"20",	--8137
		x"03",	--8138
		x"81",	--8139
		x"22",	--8140
		x"ab",	--8141
		x"3e",	--8142
		x"40",	--8143
		x"0f",	--8144
		x"3e",	--8145
		x"80",	--8146
		x"3f",	--8147
		x"a4",	--8148
		x"4d",	--8149
		x"7b",	--8150
		x"4f",	--8151
		x"de",	--8152
		x"5f",	--8153
		x"d1",	--8154
		x"11",	--8155
		x"19",	--8156
		x"06",	--8157
		x"c1",	--8158
		x"11",	--8159
		x"0f",	--8160
		x"3f",	--8161
		x"10",	--8162
		x"9e",	--8163
		x"4f",	--8164
		x"f8",	--8165
		x"6f",	--8166
		x"f1",	--8167
		x"3f",	--8168
		x"a6",	--8169
		x"97",	--8170
		x"0b",	--8171
		x"0a",	--8172
		x"09",	--8173
		x"08",	--8174
		x"07",	--8175
		x"31",	--8176
		x"e8",	--8177
		x"81",	--8178
		x"04",	--8179
		x"81",	--8180
		x"06",	--8181
		x"81",	--8182
		x"00",	--8183
		x"81",	--8184
		x"02",	--8185
		x"0e",	--8186
		x"3e",	--8187
		x"10",	--8188
		x"0f",	--8189
		x"2f",	--8190
		x"b0",	--8191
		x"1e",	--8192
		x"0e",	--8193
		x"3e",	--8194
		x"0f",	--8195
		x"b0",	--8196
		x"1e",	--8197
		x"5f",	--8198
		x"10",	--8199
		x"6f",	--8200
		x"5d",	--8201
		x"5e",	--8202
		x"08",	--8203
		x"6e",	--8204
		x"82",	--8205
		x"d1",	--8206
		x"09",	--8207
		x"11",	--8208
		x"6f",	--8209
		x"58",	--8210
		x"6f",	--8211
		x"56",	--8212
		x"6e",	--8213
		x"6f",	--8214
		x"6e",	--8215
		x"4c",	--8216
		x"1d",	--8217
		x"12",	--8218
		x"1d",	--8219
		x"0a",	--8220
		x"81",	--8221
		x"12",	--8222
		x"1e",	--8223
		x"14",	--8224
		x"1f",	--8225
		x"16",	--8226
		x"18",	--8227
		x"0c",	--8228
		x"19",	--8229
		x"0e",	--8230
		x"0f",	--8231
		x"1e",	--8232
		x"0e",	--8233
		x"0f",	--8234
		x"3d",	--8235
		x"81",	--8236
		x"12",	--8237
		x"37",	--8238
		x"1f",	--8239
		x"0c",	--8240
		x"3d",	--8241
		x"00",	--8242
		x"0a",	--8243
		x"0b",	--8244
		x"0b",	--8245
		x"0a",	--8246
		x"0b",	--8247
		x"0e",	--8248
		x"0f",	--8249
		x"12",	--8250
		x"0d",	--8251
		x"0c",	--8252
		x"0e",	--8253
		x"0f",	--8254
		x"37",	--8255
		x"0b",	--8256
		x"0f",	--8257
		x"f7",	--8258
		x"f2",	--8259
		x"0e",	--8260
		x"f4",	--8261
		x"ef",	--8262
		x"09",	--8263
		x"e5",	--8264
		x"0e",	--8265
		x"e3",	--8266
		x"dd",	--8267
		x"0c",	--8268
		x"0d",	--8269
		x"3c",	--8270
		x"7f",	--8271
		x"0d",	--8272
		x"3c",	--8273
		x"40",	--8274
		x"1c",	--8275
		x"81",	--8276
		x"14",	--8277
		x"81",	--8278
		x"16",	--8279
		x"0f",	--8280
		x"3f",	--8281
		x"10",	--8282
		x"b0",	--8283
		x"40",	--8284
		x"31",	--8285
		x"18",	--8286
		x"37",	--8287
		x"38",	--8288
		x"39",	--8289
		x"3a",	--8290
		x"3b",	--8291
		x"30",	--8292
		x"e1",	--8293
		x"10",	--8294
		x"0f",	--8295
		x"3f",	--8296
		x"10",	--8297
		x"f0",	--8298
		x"4f",	--8299
		x"fa",	--8300
		x"3f",	--8301
		x"a6",	--8302
		x"eb",	--8303
		x"0d",	--8304
		x"e2",	--8305
		x"0c",	--8306
		x"0d",	--8307
		x"3c",	--8308
		x"80",	--8309
		x"0d",	--8310
		x"0c",	--8311
		x"db",	--8312
		x"0d",	--8313
		x"d9",	--8314
		x"0e",	--8315
		x"02",	--8316
		x"0f",	--8317
		x"d5",	--8318
		x"3a",	--8319
		x"40",	--8320
		x"0b",	--8321
		x"3a",	--8322
		x"80",	--8323
		x"3b",	--8324
		x"ce",	--8325
		x"81",	--8326
		x"14",	--8327
		x"81",	--8328
		x"16",	--8329
		x"81",	--8330
		x"12",	--8331
		x"0f",	--8332
		x"3f",	--8333
		x"10",	--8334
		x"cb",	--8335
		x"0f",	--8336
		x"3f",	--8337
		x"c8",	--8338
		x"31",	--8339
		x"e8",	--8340
		x"81",	--8341
		x"04",	--8342
		x"81",	--8343
		x"06",	--8344
		x"81",	--8345
		x"00",	--8346
		x"81",	--8347
		x"02",	--8348
		x"0e",	--8349
		x"3e",	--8350
		x"10",	--8351
		x"0f",	--8352
		x"2f",	--8353
		x"b0",	--8354
		x"1e",	--8355
		x"0e",	--8356
		x"3e",	--8357
		x"0f",	--8358
		x"b0",	--8359
		x"1e",	--8360
		x"e1",	--8361
		x"10",	--8362
		x"0d",	--8363
		x"e1",	--8364
		x"08",	--8365
		x"0a",	--8366
		x"0e",	--8367
		x"3e",	--8368
		x"0f",	--8369
		x"3f",	--8370
		x"10",	--8371
		x"b0",	--8372
		x"42",	--8373
		x"31",	--8374
		x"18",	--8375
		x"30",	--8376
		x"1f",	--8377
		x"fb",	--8378
		x"31",	--8379
		x"e8",	--8380
		x"81",	--8381
		x"04",	--8382
		x"81",	--8383
		x"06",	--8384
		x"81",	--8385
		x"00",	--8386
		x"81",	--8387
		x"02",	--8388
		x"0e",	--8389
		x"3e",	--8390
		x"10",	--8391
		x"0f",	--8392
		x"2f",	--8393
		x"b0",	--8394
		x"1e",	--8395
		x"0e",	--8396
		x"3e",	--8397
		x"0f",	--8398
		x"b0",	--8399
		x"1e",	--8400
		x"e1",	--8401
		x"10",	--8402
		x"0d",	--8403
		x"e1",	--8404
		x"08",	--8405
		x"0a",	--8406
		x"0e",	--8407
		x"3e",	--8408
		x"0f",	--8409
		x"3f",	--8410
		x"10",	--8411
		x"b0",	--8412
		x"42",	--8413
		x"31",	--8414
		x"18",	--8415
		x"30",	--8416
		x"3f",	--8417
		x"fb",	--8418
		x"31",	--8419
		x"e8",	--8420
		x"81",	--8421
		x"04",	--8422
		x"81",	--8423
		x"06",	--8424
		x"81",	--8425
		x"00",	--8426
		x"81",	--8427
		x"02",	--8428
		x"0e",	--8429
		x"3e",	--8430
		x"10",	--8431
		x"0f",	--8432
		x"2f",	--8433
		x"b0",	--8434
		x"1e",	--8435
		x"0e",	--8436
		x"3e",	--8437
		x"0f",	--8438
		x"b0",	--8439
		x"1e",	--8440
		x"e1",	--8441
		x"10",	--8442
		x"0d",	--8443
		x"e1",	--8444
		x"08",	--8445
		x"0a",	--8446
		x"0e",	--8447
		x"3e",	--8448
		x"0f",	--8449
		x"3f",	--8450
		x"10",	--8451
		x"b0",	--8452
		x"42",	--8453
		x"31",	--8454
		x"18",	--8455
		x"30",	--8456
		x"3f",	--8457
		x"fb",	--8458
		x"31",	--8459
		x"e8",	--8460
		x"81",	--8461
		x"04",	--8462
		x"81",	--8463
		x"06",	--8464
		x"81",	--8465
		x"00",	--8466
		x"81",	--8467
		x"02",	--8468
		x"0e",	--8469
		x"3e",	--8470
		x"10",	--8471
		x"0f",	--8472
		x"2f",	--8473
		x"b0",	--8474
		x"1e",	--8475
		x"0e",	--8476
		x"3e",	--8477
		x"0f",	--8478
		x"b0",	--8479
		x"1e",	--8480
		x"e1",	--8481
		x"10",	--8482
		x"0d",	--8483
		x"e1",	--8484
		x"08",	--8485
		x"0a",	--8486
		x"0e",	--8487
		x"3e",	--8488
		x"0f",	--8489
		x"3f",	--8490
		x"10",	--8491
		x"b0",	--8492
		x"42",	--8493
		x"31",	--8494
		x"18",	--8495
		x"30",	--8496
		x"1f",	--8497
		x"fb",	--8498
		x"31",	--8499
		x"e8",	--8500
		x"81",	--8501
		x"04",	--8502
		x"81",	--8503
		x"06",	--8504
		x"81",	--8505
		x"00",	--8506
		x"81",	--8507
		x"02",	--8508
		x"0e",	--8509
		x"3e",	--8510
		x"10",	--8511
		x"0f",	--8512
		x"2f",	--8513
		x"b0",	--8514
		x"1e",	--8515
		x"0e",	--8516
		x"3e",	--8517
		x"0f",	--8518
		x"b0",	--8519
		x"1e",	--8520
		x"e1",	--8521
		x"10",	--8522
		x"0d",	--8523
		x"e1",	--8524
		x"08",	--8525
		x"0a",	--8526
		x"0e",	--8527
		x"3e",	--8528
		x"0f",	--8529
		x"3f",	--8530
		x"10",	--8531
		x"b0",	--8532
		x"42",	--8533
		x"31",	--8534
		x"18",	--8535
		x"30",	--8536
		x"1f",	--8537
		x"fb",	--8538
		x"0b",	--8539
		x"0a",	--8540
		x"31",	--8541
		x"f1",	--8542
		x"03",	--8543
		x"00",	--8544
		x"0d",	--8545
		x"0d",	--8546
		x"0d",	--8547
		x"0d",	--8548
		x"4c",	--8549
		x"c1",	--8550
		x"01",	--8551
		x"0e",	--8552
		x"0b",	--8553
		x"0f",	--8554
		x"09",	--8555
		x"e1",	--8556
		x"00",	--8557
		x"0f",	--8558
		x"b0",	--8559
		x"40",	--8560
		x"31",	--8561
		x"3a",	--8562
		x"3b",	--8563
		x"30",	--8564
		x"b1",	--8565
		x"1e",	--8566
		x"02",	--8567
		x"4c",	--8568
		x"1b",	--8569
		x"0a",	--8570
		x"0b",	--8571
		x"81",	--8572
		x"04",	--8573
		x"81",	--8574
		x"06",	--8575
		x"0e",	--8576
		x"0f",	--8577
		x"b0",	--8578
		x"ce",	--8579
		x"3f",	--8580
		x"1f",	--8581
		x"e7",	--8582
		x"81",	--8583
		x"04",	--8584
		x"81",	--8585
		x"06",	--8586
		x"4e",	--8587
		x"7e",	--8588
		x"1f",	--8589
		x"0f",	--8590
		x"3e",	--8591
		x"1e",	--8592
		x"0e",	--8593
		x"81",	--8594
		x"02",	--8595
		x"d9",	--8596
		x"0e",	--8597
		x"10",	--8598
		x"0a",	--8599
		x"0b",	--8600
		x"3a",	--8601
		x"3b",	--8602
		x"1a",	--8603
		x"0b",	--8604
		x"de",	--8605
		x"91",	--8606
		x"04",	--8607
		x"04",	--8608
		x"91",	--8609
		x"06",	--8610
		x"06",	--8611
		x"7e",	--8612
		x"f8",	--8613
		x"e8",	--8614
		x"3f",	--8615
		x"00",	--8616
		x"ed",	--8617
		x"0e",	--8618
		x"3f",	--8619
		x"00",	--8620
		x"c3",	--8621
		x"31",	--8622
		x"f4",	--8623
		x"81",	--8624
		x"00",	--8625
		x"81",	--8626
		x"02",	--8627
		x"0e",	--8628
		x"2e",	--8629
		x"0f",	--8630
		x"b0",	--8631
		x"1e",	--8632
		x"5f",	--8633
		x"04",	--8634
		x"6f",	--8635
		x"28",	--8636
		x"27",	--8637
		x"6f",	--8638
		x"07",	--8639
		x"1d",	--8640
		x"06",	--8641
		x"0d",	--8642
		x"21",	--8643
		x"3d",	--8644
		x"1f",	--8645
		x"09",	--8646
		x"c1",	--8647
		x"05",	--8648
		x"26",	--8649
		x"3e",	--8650
		x"3f",	--8651
		x"ff",	--8652
		x"31",	--8653
		x"0c",	--8654
		x"30",	--8655
		x"1e",	--8656
		x"08",	--8657
		x"1f",	--8658
		x"0a",	--8659
		x"3c",	--8660
		x"1e",	--8661
		x"4c",	--8662
		x"4d",	--8663
		x"7d",	--8664
		x"1f",	--8665
		x"0f",	--8666
		x"c1",	--8667
		x"05",	--8668
		x"ef",	--8669
		x"3e",	--8670
		x"3f",	--8671
		x"1e",	--8672
		x"0f",	--8673
		x"31",	--8674
		x"0c",	--8675
		x"30",	--8676
		x"0e",	--8677
		x"0f",	--8678
		x"31",	--8679
		x"0c",	--8680
		x"30",	--8681
		x"12",	--8682
		x"0f",	--8683
		x"0e",	--8684
		x"7d",	--8685
		x"fb",	--8686
		x"eb",	--8687
		x"0e",	--8688
		x"3f",	--8689
		x"00",	--8690
		x"31",	--8691
		x"0c",	--8692
		x"30",	--8693
		x"0b",	--8694
		x"0a",	--8695
		x"09",	--8696
		x"08",	--8697
		x"31",	--8698
		x"0a",	--8699
		x"0b",	--8700
		x"c1",	--8701
		x"01",	--8702
		x"0e",	--8703
		x"0d",	--8704
		x"0b",	--8705
		x"0b",	--8706
		x"e1",	--8707
		x"00",	--8708
		x"0f",	--8709
		x"b0",	--8710
		x"40",	--8711
		x"31",	--8712
		x"38",	--8713
		x"39",	--8714
		x"3a",	--8715
		x"3b",	--8716
		x"30",	--8717
		x"f1",	--8718
		x"03",	--8719
		x"00",	--8720
		x"b1",	--8721
		x"1e",	--8722
		x"02",	--8723
		x"81",	--8724
		x"04",	--8725
		x"81",	--8726
		x"06",	--8727
		x"0e",	--8728
		x"0f",	--8729
		x"b0",	--8730
		x"ce",	--8731
		x"3f",	--8732
		x"0f",	--8733
		x"18",	--8734
		x"e5",	--8735
		x"81",	--8736
		x"04",	--8737
		x"81",	--8738
		x"06",	--8739
		x"4e",	--8740
		x"7e",	--8741
		x"1f",	--8742
		x"06",	--8743
		x"3e",	--8744
		x"1e",	--8745
		x"0e",	--8746
		x"81",	--8747
		x"02",	--8748
		x"d7",	--8749
		x"91",	--8750
		x"04",	--8751
		x"04",	--8752
		x"91",	--8753
		x"06",	--8754
		x"06",	--8755
		x"7e",	--8756
		x"f8",	--8757
		x"f1",	--8758
		x"0e",	--8759
		x"3e",	--8760
		x"1e",	--8761
		x"1c",	--8762
		x"0d",	--8763
		x"48",	--8764
		x"78",	--8765
		x"1f",	--8766
		x"04",	--8767
		x"0c",	--8768
		x"0d",	--8769
		x"78",	--8770
		x"fc",	--8771
		x"3c",	--8772
		x"3d",	--8773
		x"0c",	--8774
		x"0d",	--8775
		x"18",	--8776
		x"09",	--8777
		x"0c",	--8778
		x"04",	--8779
		x"0d",	--8780
		x"02",	--8781
		x"08",	--8782
		x"09",	--8783
		x"7e",	--8784
		x"1f",	--8785
		x"0e",	--8786
		x"0d",	--8787
		x"0e",	--8788
		x"0d",	--8789
		x"0e",	--8790
		x"81",	--8791
		x"04",	--8792
		x"81",	--8793
		x"06",	--8794
		x"3e",	--8795
		x"1e",	--8796
		x"0e",	--8797
		x"81",	--8798
		x"02",	--8799
		x"a4",	--8800
		x"12",	--8801
		x"0b",	--8802
		x"0a",	--8803
		x"7e",	--8804
		x"fb",	--8805
		x"ec",	--8806
		x"0b",	--8807
		x"0a",	--8808
		x"09",	--8809
		x"1f",	--8810
		x"17",	--8811
		x"3e",	--8812
		x"00",	--8813
		x"2c",	--8814
		x"3a",	--8815
		x"18",	--8816
		x"0b",	--8817
		x"39",	--8818
		x"0c",	--8819
		x"0d",	--8820
		x"4f",	--8821
		x"4f",	--8822
		x"17",	--8823
		x"3c",	--8824
		x"ae",	--8825
		x"6e",	--8826
		x"0f",	--8827
		x"0a",	--8828
		x"0b",	--8829
		x"0f",	--8830
		x"39",	--8831
		x"3a",	--8832
		x"3b",	--8833
		x"30",	--8834
		x"3f",	--8835
		x"00",	--8836
		x"0f",	--8837
		x"3a",	--8838
		x"0b",	--8839
		x"39",	--8840
		x"18",	--8841
		x"0c",	--8842
		x"0d",	--8843
		x"4f",	--8844
		x"4f",	--8845
		x"e9",	--8846
		x"12",	--8847
		x"0d",	--8848
		x"0c",	--8849
		x"7f",	--8850
		x"fb",	--8851
		x"e3",	--8852
		x"3a",	--8853
		x"10",	--8854
		x"0b",	--8855
		x"39",	--8856
		x"10",	--8857
		x"ef",	--8858
		x"3a",	--8859
		x"20",	--8860
		x"0b",	--8861
		x"09",	--8862
		x"ea",	--8863
		x"0b",	--8864
		x"0a",	--8865
		x"09",	--8866
		x"08",	--8867
		x"07",	--8868
		x"0d",	--8869
		x"1e",	--8870
		x"04",	--8871
		x"1f",	--8872
		x"06",	--8873
		x"5a",	--8874
		x"01",	--8875
		x"6c",	--8876
		x"6c",	--8877
		x"70",	--8878
		x"6c",	--8879
		x"6a",	--8880
		x"6c",	--8881
		x"36",	--8882
		x"0e",	--8883
		x"32",	--8884
		x"1b",	--8885
		x"02",	--8886
		x"3b",	--8887
		x"82",	--8888
		x"6d",	--8889
		x"3b",	--8890
		x"80",	--8891
		x"5e",	--8892
		x"0c",	--8893
		x"0d",	--8894
		x"3c",	--8895
		x"7f",	--8896
		x"0d",	--8897
		x"3c",	--8898
		x"40",	--8899
		x"40",	--8900
		x"3e",	--8901
		x"3f",	--8902
		x"0f",	--8903
		x"0f",	--8904
		x"4a",	--8905
		x"0d",	--8906
		x"3d",	--8907
		x"7f",	--8908
		x"12",	--8909
		x"0f",	--8910
		x"0e",	--8911
		x"12",	--8912
		x"0f",	--8913
		x"0e",	--8914
		x"12",	--8915
		x"0f",	--8916
		x"0e",	--8917
		x"12",	--8918
		x"0f",	--8919
		x"0e",	--8920
		x"12",	--8921
		x"0f",	--8922
		x"0e",	--8923
		x"12",	--8924
		x"0f",	--8925
		x"0e",	--8926
		x"12",	--8927
		x"0f",	--8928
		x"0e",	--8929
		x"3e",	--8930
		x"3f",	--8931
		x"7f",	--8932
		x"4d",	--8933
		x"05",	--8934
		x"0f",	--8935
		x"cc",	--8936
		x"4d",	--8937
		x"0e",	--8938
		x"0f",	--8939
		x"4d",	--8940
		x"0d",	--8941
		x"0d",	--8942
		x"0d",	--8943
		x"0d",	--8944
		x"0d",	--8945
		x"0d",	--8946
		x"0d",	--8947
		x"0c",	--8948
		x"3c",	--8949
		x"7f",	--8950
		x"0c",	--8951
		x"4f",	--8952
		x"0f",	--8953
		x"0f",	--8954
		x"0f",	--8955
		x"0d",	--8956
		x"0d",	--8957
		x"0f",	--8958
		x"37",	--8959
		x"38",	--8960
		x"39",	--8961
		x"3a",	--8962
		x"3b",	--8963
		x"30",	--8964
		x"0d",	--8965
		x"be",	--8966
		x"0c",	--8967
		x"0d",	--8968
		x"3c",	--8969
		x"80",	--8970
		x"0d",	--8971
		x"0c",	--8972
		x"02",	--8973
		x"0d",	--8974
		x"b8",	--8975
		x"3e",	--8976
		x"40",	--8977
		x"0f",	--8978
		x"b4",	--8979
		x"12",	--8980
		x"0f",	--8981
		x"0e",	--8982
		x"0d",	--8983
		x"3d",	--8984
		x"80",	--8985
		x"b2",	--8986
		x"7d",	--8987
		x"0e",	--8988
		x"0f",	--8989
		x"cd",	--8990
		x"0e",	--8991
		x"3f",	--8992
		x"10",	--8993
		x"3e",	--8994
		x"3f",	--8995
		x"7f",	--8996
		x"7d",	--8997
		x"c5",	--8998
		x"37",	--8999
		x"82",	--9000
		x"07",	--9001
		x"37",	--9002
		x"1a",	--9003
		x"4f",	--9004
		x"0c",	--9005
		x"0d",	--9006
		x"4b",	--9007
		x"7b",	--9008
		x"1f",	--9009
		x"05",	--9010
		x"12",	--9011
		x"0d",	--9012
		x"0c",	--9013
		x"7b",	--9014
		x"fb",	--9015
		x"18",	--9016
		x"09",	--9017
		x"77",	--9018
		x"1f",	--9019
		x"04",	--9020
		x"08",	--9021
		x"09",	--9022
		x"77",	--9023
		x"fc",	--9024
		x"38",	--9025
		x"39",	--9026
		x"08",	--9027
		x"09",	--9028
		x"1e",	--9029
		x"0f",	--9030
		x"08",	--9031
		x"04",	--9032
		x"09",	--9033
		x"02",	--9034
		x"0e",	--9035
		x"0f",	--9036
		x"08",	--9037
		x"09",	--9038
		x"08",	--9039
		x"09",	--9040
		x"0e",	--9041
		x"0f",	--9042
		x"3e",	--9043
		x"7f",	--9044
		x"0f",	--9045
		x"3e",	--9046
		x"40",	--9047
		x"26",	--9048
		x"38",	--9049
		x"3f",	--9050
		x"09",	--9051
		x"0e",	--9052
		x"0f",	--9053
		x"12",	--9054
		x"0f",	--9055
		x"0e",	--9056
		x"12",	--9057
		x"0f",	--9058
		x"0e",	--9059
		x"12",	--9060
		x"0f",	--9061
		x"0e",	--9062
		x"12",	--9063
		x"0f",	--9064
		x"0e",	--9065
		x"12",	--9066
		x"0f",	--9067
		x"0e",	--9068
		x"12",	--9069
		x"0f",	--9070
		x"0e",	--9071
		x"12",	--9072
		x"0f",	--9073
		x"0e",	--9074
		x"3e",	--9075
		x"3f",	--9076
		x"7f",	--9077
		x"5d",	--9078
		x"39",	--9079
		x"00",	--9080
		x"72",	--9081
		x"4d",	--9082
		x"70",	--9083
		x"08",	--9084
		x"09",	--9085
		x"da",	--9086
		x"0f",	--9087
		x"d8",	--9088
		x"0e",	--9089
		x"0f",	--9090
		x"3e",	--9091
		x"80",	--9092
		x"0f",	--9093
		x"0e",	--9094
		x"04",	--9095
		x"38",	--9096
		x"40",	--9097
		x"09",	--9098
		x"d0",	--9099
		x"0f",	--9100
		x"ce",	--9101
		x"f9",	--9102
		x"0b",	--9103
		x"0a",	--9104
		x"2a",	--9105
		x"5b",	--9106
		x"02",	--9107
		x"3b",	--9108
		x"7f",	--9109
		x"1d",	--9110
		x"02",	--9111
		x"12",	--9112
		x"0d",	--9113
		x"12",	--9114
		x"0d",	--9115
		x"12",	--9116
		x"0d",	--9117
		x"12",	--9118
		x"0d",	--9119
		x"12",	--9120
		x"0d",	--9121
		x"12",	--9122
		x"0d",	--9123
		x"12",	--9124
		x"0d",	--9125
		x"4d",	--9126
		x"5f",	--9127
		x"03",	--9128
		x"3f",	--9129
		x"80",	--9130
		x"0f",	--9131
		x"0f",	--9132
		x"ce",	--9133
		x"01",	--9134
		x"0d",	--9135
		x"2d",	--9136
		x"0a",	--9137
		x"51",	--9138
		x"be",	--9139
		x"82",	--9140
		x"02",	--9141
		x"0c",	--9142
		x"0d",	--9143
		x"0c",	--9144
		x"0d",	--9145
		x"0c",	--9146
		x"0d",	--9147
		x"0c",	--9148
		x"0d",	--9149
		x"0c",	--9150
		x"0d",	--9151
		x"0c",	--9152
		x"0d",	--9153
		x"0c",	--9154
		x"0d",	--9155
		x"0c",	--9156
		x"0d",	--9157
		x"fe",	--9158
		x"03",	--9159
		x"00",	--9160
		x"3d",	--9161
		x"00",	--9162
		x"0b",	--9163
		x"3f",	--9164
		x"81",	--9165
		x"0c",	--9166
		x"0d",	--9167
		x"0a",	--9168
		x"3f",	--9169
		x"3d",	--9170
		x"00",	--9171
		x"f9",	--9172
		x"8e",	--9173
		x"02",	--9174
		x"8e",	--9175
		x"04",	--9176
		x"8e",	--9177
		x"06",	--9178
		x"3a",	--9179
		x"3b",	--9180
		x"30",	--9181
		x"3d",	--9182
		x"ff",	--9183
		x"2a",	--9184
		x"3d",	--9185
		x"81",	--9186
		x"8e",	--9187
		x"02",	--9188
		x"fe",	--9189
		x"03",	--9190
		x"00",	--9191
		x"0c",	--9192
		x"0d",	--9193
		x"0c",	--9194
		x"0d",	--9195
		x"0c",	--9196
		x"0d",	--9197
		x"0c",	--9198
		x"0d",	--9199
		x"0c",	--9200
		x"0d",	--9201
		x"0c",	--9202
		x"0d",	--9203
		x"0c",	--9204
		x"0d",	--9205
		x"0c",	--9206
		x"0d",	--9207
		x"0a",	--9208
		x"0b",	--9209
		x"0a",	--9210
		x"3b",	--9211
		x"00",	--9212
		x"8e",	--9213
		x"04",	--9214
		x"8e",	--9215
		x"06",	--9216
		x"3a",	--9217
		x"3b",	--9218
		x"30",	--9219
		x"0b",	--9220
		x"ad",	--9221
		x"ee",	--9222
		x"00",	--9223
		x"3a",	--9224
		x"3b",	--9225
		x"30",	--9226
		x"0a",	--9227
		x"0c",	--9228
		x"0c",	--9229
		x"0d",	--9230
		x"0c",	--9231
		x"3d",	--9232
		x"10",	--9233
		x"0c",	--9234
		x"02",	--9235
		x"0d",	--9236
		x"08",	--9237
		x"de",	--9238
		x"00",	--9239
		x"e4",	--9240
		x"0b",	--9241
		x"f2",	--9242
		x"ee",	--9243
		x"00",	--9244
		x"e3",	--9245
		x"ce",	--9246
		x"00",	--9247
		x"dc",	--9248
		x"0b",	--9249
		x"6d",	--9250
		x"6d",	--9251
		x"12",	--9252
		x"6c",	--9253
		x"6c",	--9254
		x"0f",	--9255
		x"6d",	--9256
		x"41",	--9257
		x"6c",	--9258
		x"11",	--9259
		x"6d",	--9260
		x"0d",	--9261
		x"6c",	--9262
		x"14",	--9263
		x"5d",	--9264
		x"01",	--9265
		x"5d",	--9266
		x"01",	--9267
		x"14",	--9268
		x"4d",	--9269
		x"09",	--9270
		x"1e",	--9271
		x"0f",	--9272
		x"3b",	--9273
		x"30",	--9274
		x"6c",	--9275
		x"28",	--9276
		x"ce",	--9277
		x"01",	--9278
		x"f7",	--9279
		x"3e",	--9280
		x"0f",	--9281
		x"3b",	--9282
		x"30",	--9283
		x"cf",	--9284
		x"01",	--9285
		x"f0",	--9286
		x"3e",	--9287
		x"f8",	--9288
		x"1b",	--9289
		x"02",	--9290
		x"1c",	--9291
		x"02",	--9292
		x"0c",	--9293
		x"e6",	--9294
		x"0b",	--9295
		x"16",	--9296
		x"1b",	--9297
		x"04",	--9298
		x"1f",	--9299
		x"06",	--9300
		x"1c",	--9301
		x"04",	--9302
		x"1e",	--9303
		x"06",	--9304
		x"0e",	--9305
		x"da",	--9306
		x"0f",	--9307
		x"02",	--9308
		x"0c",	--9309
		x"d6",	--9310
		x"0f",	--9311
		x"06",	--9312
		x"0e",	--9313
		x"02",	--9314
		x"0b",	--9315
		x"02",	--9316
		x"0e",	--9317
		x"d1",	--9318
		x"4d",	--9319
		x"ce",	--9320
		x"3e",	--9321
		x"d6",	--9322
		x"6c",	--9323
		x"d7",	--9324
		x"5e",	--9325
		x"01",	--9326
		x"5f",	--9327
		x"01",	--9328
		x"0e",	--9329
		x"c5",	--9330
		x"1e",	--9331
		x"34",	--9332
		x"1e",	--9333
		x"0b",	--9334
		x"1d",	--9335
		x"32",	--9336
		x"cd",	--9337
		x"00",	--9338
		x"1d",	--9339
		x"82",	--9340
		x"32",	--9341
		x"3e",	--9342
		x"82",	--9343
		x"34",	--9344
		x"30",	--9345
		x"3f",	--9346
		x"30",	--9347
		x"0b",	--9348
		x"0a",	--9349
		x"21",	--9350
		x"81",	--9351
		x"00",	--9352
		x"1a",	--9353
		x"32",	--9354
		x"1b",	--9355
		x"34",	--9356
		x"0d",	--9357
		x"0e",	--9358
		x"3f",	--9359
		x"e6",	--9360
		x"b0",	--9361
		x"3a",	--9362
		x"0f",	--9363
		x"05",	--9364
		x"0e",	--9365
		x"0e",	--9366
		x"ce",	--9367
		x"ff",	--9368
		x"04",	--9369
		x"1e",	--9370
		x"32",	--9371
		x"ce",	--9372
		x"00",	--9373
		x"21",	--9374
		x"3a",	--9375
		x"3b",	--9376
		x"30",	--9377
		x"92",	--9378
		x"02",	--9379
		x"32",	--9380
		x"b2",	--9381
		x"ff",	--9382
		x"34",	--9383
		x"0e",	--9384
		x"3e",	--9385
		x"06",	--9386
		x"1f",	--9387
		x"04",	--9388
		x"b0",	--9389
		x"08",	--9390
		x"30",	--9391
		x"92",	--9392
		x"02",	--9393
		x"32",	--9394
		x"92",	--9395
		x"04",	--9396
		x"34",	--9397
		x"0e",	--9398
		x"3e",	--9399
		x"1f",	--9400
		x"06",	--9401
		x"b0",	--9402
		x"08",	--9403
		x"30",	--9404
		x"0c",	--9405
		x"82",	--9406
		x"32",	--9407
		x"b2",	--9408
		x"ff",	--9409
		x"34",	--9410
		x"0e",	--9411
		x"0f",	--9412
		x"b0",	--9413
		x"08",	--9414
		x"30",	--9415
		x"82",	--9416
		x"32",	--9417
		x"82",	--9418
		x"34",	--9419
		x"0e",	--9420
		x"0f",	--9421
		x"b0",	--9422
		x"08",	--9423
		x"30",	--9424
		x"0b",	--9425
		x"0a",	--9426
		x"09",	--9427
		x"08",	--9428
		x"07",	--9429
		x"06",	--9430
		x"05",	--9431
		x"04",	--9432
		x"31",	--9433
		x"08",	--9434
		x"81",	--9435
		x"04",	--9436
		x"09",	--9437
		x"1f",	--9438
		x"1a",	--9439
		x"1d",	--9440
		x"1c",	--9441
		x"4c",	--9442
		x"04",	--9443
		x"84",	--9444
		x"45",	--9445
		x"4e",	--9446
		x"7e",	--9447
		x"40",	--9448
		x"11",	--9449
		x"f1",	--9450
		x"30",	--9451
		x"00",	--9452
		x"0e",	--9453
		x"8e",	--9454
		x"5e",	--9455
		x"03",	--9456
		x"7e",	--9457
		x"58",	--9458
		x"02",	--9459
		x"7e",	--9460
		x"78",	--9461
		x"c1",	--9462
		x"01",	--9463
		x"0c",	--9464
		x"2c",	--9465
		x"0f",	--9466
		x"7e",	--9467
		x"20",	--9468
		x"04",	--9469
		x"f1",	--9470
		x"30",	--9471
		x"00",	--9472
		x"04",	--9473
		x"4c",	--9474
		x"05",	--9475
		x"c1",	--9476
		x"00",	--9477
		x"0c",	--9478
		x"1c",	--9479
		x"01",	--9480
		x"0c",	--9481
		x"0a",	--9482
		x"8c",	--9483
		x"8c",	--9484
		x"8c",	--9485
		x"8c",	--9486
		x"0b",	--9487
		x"06",	--9488
		x"0c",	--9489
		x"8c",	--9490
		x"8c",	--9491
		x"8c",	--9492
		x"8c",	--9493
		x"07",	--9494
		x"0a",	--9495
		x"0b",	--9496
		x"0e",	--9497
		x"8e",	--9498
		x"c1",	--9499
		x"02",	--9500
		x"6e",	--9501
		x"02",	--9502
		x"07",	--9503
		x"01",	--9504
		x"37",	--9505
		x"4f",	--9506
		x"7f",	--9507
		x"10",	--9508
		x"3c",	--9509
		x"1d",	--9510
		x"04",	--9511
		x"3d",	--9512
		x"1d",	--9513
		x"cd",	--9514
		x"00",	--9515
		x"fc",	--9516
		x"1d",	--9517
		x"04",	--9518
		x"09",	--9519
		x"02",	--9520
		x"09",	--9521
		x"01",	--9522
		x"09",	--9523
		x"e1",	--9524
		x"02",	--9525
		x"05",	--9526
		x"09",	--9527
		x"02",	--9528
		x"09",	--9529
		x"01",	--9530
		x"09",	--9531
		x"05",	--9532
		x"07",	--9533
		x"01",	--9534
		x"05",	--9535
		x"4f",	--9536
		x"0d",	--9537
		x"f1",	--9538
		x"20",	--9539
		x"06",	--9540
		x"06",	--9541
		x"0b",	--9542
		x"0e",	--9543
		x"0f",	--9544
		x"0f",	--9545
		x"6f",	--9546
		x"8f",	--9547
		x"16",	--9548
		x"88",	--9549
		x"01",	--9550
		x"06",	--9551
		x"06",	--9552
		x"f6",	--9553
		x"0b",	--9554
		x"f1",	--9555
		x"30",	--9556
		x"06",	--9557
		x"05",	--9558
		x"05",	--9559
		x"5f",	--9560
		x"06",	--9561
		x"8f",	--9562
		x"88",	--9563
		x"1b",	--9564
		x"0f",	--9565
		x"0f",	--9566
		x"0f",	--9567
		x"f7",	--9568
		x"0a",	--9569
		x"06",	--9570
		x"0b",	--9571
		x"07",	--9572
		x"1b",	--9573
		x"0f",	--9574
		x"0f",	--9575
		x"6f",	--9576
		x"8f",	--9577
		x"16",	--9578
		x"88",	--9579
		x"06",	--9580
		x"f7",	--9581
		x"e1",	--9582
		x"02",	--9583
		x"02",	--9584
		x"4a",	--9585
		x"08",	--9586
		x"1a",	--9587
		x"04",	--9588
		x"0a",	--9589
		x"0d",	--9590
		x"3f",	--9591
		x"30",	--9592
		x"88",	--9593
		x"7a",	--9594
		x"4a",	--9595
		x"fa",	--9596
		x"44",	--9597
		x"0b",	--9598
		x"f3",	--9599
		x"37",	--9600
		x"8f",	--9601
		x"88",	--9602
		x"1b",	--9603
		x"0f",	--9604
		x"0f",	--9605
		x"6f",	--9606
		x"4f",	--9607
		x"07",	--9608
		x"07",	--9609
		x"f5",	--9610
		x"04",	--9611
		x"3f",	--9612
		x"20",	--9613
		x"88",	--9614
		x"1b",	--9615
		x"0b",	--9616
		x"fa",	--9617
		x"0f",	--9618
		x"31",	--9619
		x"34",	--9620
		x"35",	--9621
		x"36",	--9622
		x"37",	--9623
		x"38",	--9624
		x"39",	--9625
		x"3a",	--9626
		x"3b",	--9627
		x"30",	--9628
		x"0b",	--9629
		x"0a",	--9630
		x"09",	--9631
		x"08",	--9632
		x"07",	--9633
		x"06",	--9634
		x"05",	--9635
		x"04",	--9636
		x"31",	--9637
		x"b6",	--9638
		x"81",	--9639
		x"3a",	--9640
		x"06",	--9641
		x"05",	--9642
		x"81",	--9643
		x"3e",	--9644
		x"c1",	--9645
		x"2f",	--9646
		x"c1",	--9647
		x"2b",	--9648
		x"c1",	--9649
		x"2e",	--9650
		x"c1",	--9651
		x"2a",	--9652
		x"81",	--9653
		x"30",	--9654
		x"81",	--9655
		x"26",	--9656
		x"07",	--9657
		x"81",	--9658
		x"2c",	--9659
		x"0e",	--9660
		x"3e",	--9661
		x"1c",	--9662
		x"81",	--9663
		x"1c",	--9664
		x"30",	--9665
		x"b4",	--9666
		x"0f",	--9667
		x"1f",	--9668
		x"81",	--9669
		x"40",	--9670
		x"07",	--9671
		x"1e",	--9672
		x"7e",	--9673
		x"25",	--9674
		x"13",	--9675
		x"81",	--9676
		x"00",	--9677
		x"81",	--9678
		x"02",	--9679
		x"81",	--9680
		x"3e",	--9681
		x"c1",	--9682
		x"2f",	--9683
		x"c1",	--9684
		x"2b",	--9685
		x"c1",	--9686
		x"2e",	--9687
		x"c1",	--9688
		x"2a",	--9689
		x"81",	--9690
		x"30",	--9691
		x"30",	--9692
		x"aa",	--9693
		x"05",	--9694
		x"8e",	--9695
		x"0f",	--9696
		x"91",	--9697
		x"3c",	--9698
		x"91",	--9699
		x"2c",	--9700
		x"30",	--9701
		x"90",	--9702
		x"7e",	--9703
		x"63",	--9704
		x"c5",	--9705
		x"7e",	--9706
		x"64",	--9707
		x"27",	--9708
		x"7e",	--9709
		x"30",	--9710
		x"94",	--9711
		x"7e",	--9712
		x"31",	--9713
		x"1a",	--9714
		x"7e",	--9715
		x"2a",	--9716
		x"77",	--9717
		x"7e",	--9718
		x"2b",	--9719
		x"0a",	--9720
		x"7e",	--9721
		x"23",	--9722
		x"42",	--9723
		x"7e",	--9724
		x"25",	--9725
		x"e0",	--9726
		x"7e",	--9727
		x"20",	--9728
		x"32",	--9729
		x"56",	--9730
		x"7e",	--9731
		x"2d",	--9732
		x"49",	--9733
		x"7e",	--9734
		x"2e",	--9735
		x"5b",	--9736
		x"7e",	--9737
		x"2b",	--9738
		x"28",	--9739
		x"47",	--9740
		x"7e",	--9741
		x"3a",	--9742
		x"8c",	--9743
		x"7e",	--9744
		x"58",	--9745
		x"21",	--9746
		x"e9",	--9747
		x"7e",	--9748
		x"6f",	--9749
		x"24",	--9750
		x"7e",	--9751
		x"70",	--9752
		x"0a",	--9753
		x"7e",	--9754
		x"69",	--9755
		x"e3",	--9756
		x"7e",	--9757
		x"6c",	--9758
		x"22",	--9759
		x"7e",	--9760
		x"64",	--9761
		x"11",	--9762
		x"dc",	--9763
		x"7e",	--9764
		x"73",	--9765
		x"98",	--9766
		x"7e",	--9767
		x"74",	--9768
		x"04",	--9769
		x"7e",	--9770
		x"70",	--9771
		x"07",	--9772
		x"b8",	--9773
		x"7e",	--9774
		x"75",	--9775
		x"d1",	--9776
		x"7e",	--9777
		x"78",	--9778
		x"d2",	--9779
		x"19",	--9780
		x"3e",	--9781
		x"18",	--9782
		x"2c",	--9783
		x"08",	--9784
		x"30",	--9785
		x"7e",	--9786
		x"b1",	--9787
		x"28",	--9788
		x"cb",	--9789
		x"f1",	--9790
		x"00",	--9791
		x"30",	--9792
		x"ae",	--9793
		x"69",	--9794
		x"59",	--9795
		x"6e",	--9796
		x"04",	--9797
		x"7e",	--9798
		x"fe",	--9799
		x"6e",	--9800
		x"01",	--9801
		x"5e",	--9802
		x"c1",	--9803
		x"00",	--9804
		x"30",	--9805
		x"ae",	--9806
		x"f1",	--9807
		x"10",	--9808
		x"00",	--9809
		x"30",	--9810
		x"ae",	--9811
		x"f1",	--9812
		x"2b",	--9813
		x"02",	--9814
		x"30",	--9815
		x"ae",	--9816
		x"f1",	--9817
		x"2b",	--9818
		x"02",	--9819
		x"02",	--9820
		x"30",	--9821
		x"ae",	--9822
		x"f1",	--9823
		x"20",	--9824
		x"02",	--9825
		x"30",	--9826
		x"ae",	--9827
		x"c1",	--9828
		x"2a",	--9829
		x"02",	--9830
		x"30",	--9831
		x"94",	--9832
		x"d1",	--9833
		x"2e",	--9834
		x"30",	--9835
		x"ae",	--9836
		x"0e",	--9837
		x"2e",	--9838
		x"2a",	--9839
		x"0a",	--9840
		x"03",	--9841
		x"81",	--9842
		x"26",	--9843
		x"0d",	--9844
		x"c1",	--9845
		x"2e",	--9846
		x"02",	--9847
		x"30",	--9848
		x"a4",	--9849
		x"f1",	--9850
		x"10",	--9851
		x"00",	--9852
		x"3a",	--9853
		x"81",	--9854
		x"26",	--9855
		x"91",	--9856
		x"26",	--9857
		x"05",	--9858
		x"27",	--9859
		x"81",	--9860
		x"26",	--9861
		x"15",	--9862
		x"c1",	--9863
		x"2e",	--9864
		x"12",	--9865
		x"69",	--9866
		x"79",	--9867
		x"10",	--9868
		x"5e",	--9869
		x"01",	--9870
		x"4e",	--9871
		x"4e",	--9872
		x"0e",	--9873
		x"0e",	--9874
		x"4e",	--9875
		x"6a",	--9876
		x"7a",	--9877
		x"7f",	--9878
		x"4a",	--9879
		x"c1",	--9880
		x"00",	--9881
		x"30",	--9882
		x"ae",	--9883
		x"1a",	--9884
		x"26",	--9885
		x"0a",	--9886
		x"0c",	--9887
		x"0c",	--9888
		x"0c",	--9889
		x"0a",	--9890
		x"81",	--9891
		x"26",	--9892
		x"b1",	--9893
		x"d0",	--9894
		x"26",	--9895
		x"8e",	--9896
		x"81",	--9897
		x"26",	--9898
		x"d1",	--9899
		x"2a",	--9900
		x"30",	--9901
		x"ae",	--9902
		x"07",	--9903
		x"27",	--9904
		x"6e",	--9905
		x"c1",	--9906
		x"2e",	--9907
		x"03",	--9908
		x"c1",	--9909
		x"2a",	--9910
		x"26",	--9911
		x"c1",	--9912
		x"04",	--9913
		x"c1",	--9914
		x"05",	--9915
		x"0e",	--9916
		x"2e",	--9917
		x"03",	--9918
		x"07",	--9919
		x"27",	--9920
		x"2e",	--9921
		x"c1",	--9922
		x"2e",	--9923
		x"07",	--9924
		x"e1",	--9925
		x"01",	--9926
		x"1f",	--9927
		x"26",	--9928
		x"c1",	--9929
		x"03",	--9930
		x"06",	--9931
		x"c1",	--9932
		x"2a",	--9933
		x"03",	--9934
		x"91",	--9935
		x"26",	--9936
		x"30",	--9937
		x"0e",	--9938
		x"02",	--9939
		x"3e",	--9940
		x"ae",	--9941
		x"11",	--9942
		x"04",	--9943
		x"11",	--9944
		x"04",	--9945
		x"1d",	--9946
		x"34",	--9947
		x"1f",	--9948
		x"3e",	--9949
		x"b0",	--9950
		x"a2",	--9951
		x"21",	--9952
		x"81",	--9953
		x"2c",	--9954
		x"05",	--9955
		x"30",	--9956
		x"90",	--9957
		x"07",	--9958
		x"27",	--9959
		x"29",	--9960
		x"81",	--9961
		x"1e",	--9962
		x"5e",	--9963
		x"09",	--9964
		x"01",	--9965
		x"4e",	--9966
		x"4e",	--9967
		x"4e",	--9968
		x"4e",	--9969
		x"6a",	--9970
		x"7a",	--9971
		x"f7",	--9972
		x"4a",	--9973
		x"c1",	--9974
		x"00",	--9975
		x"05",	--9976
		x"b1",	--9977
		x"10",	--9978
		x"28",	--9979
		x"53",	--9980
		x"d1",	--9981
		x"01",	--9982
		x"06",	--9983
		x"e1",	--9984
		x"00",	--9985
		x"b1",	--9986
		x"0a",	--9987
		x"28",	--9988
		x"03",	--9989
		x"b1",	--9990
		x"10",	--9991
		x"28",	--9992
		x"6b",	--9993
		x"6b",	--9994
		x"24",	--9995
		x"0c",	--9996
		x"3c",	--9997
		x"28",	--9998
		x"17",	--9999
		x"02",	--10000
		x"16",	--10001
		x"04",	--10002
		x"1b",	--10003
		x"06",	--10004
		x"81",	--10005
		x"1e",	--10006
		x"81",	--10007
		x"20",	--10008
		x"81",	--10009
		x"22",	--10010
		x"81",	--10011
		x"24",	--10012
		x"d1",	--10013
		x"2b",	--10014
		x"08",	--10015
		x"06",	--10016
		x"07",	--10017
		x"04",	--10018
		x"06",	--10019
		x"02",	--10020
		x"0b",	--10021
		x"02",	--10022
		x"c1",	--10023
		x"2b",	--10024
		x"0b",	--10025
		x"0b",	--10026
		x"0b",	--10027
		x"c1",	--10028
		x"2f",	--10029
		x"05",	--10030
		x"20",	--10031
		x"5b",	--10032
		x"07",	--10033
		x"0d",	--10034
		x"27",	--10035
		x"28",	--10036
		x"1b",	--10037
		x"02",	--10038
		x"81",	--10039
		x"1e",	--10040
		x"81",	--10041
		x"20",	--10042
		x"d1",	--10043
		x"2b",	--10044
		x"08",	--10045
		x"09",	--10046
		x"06",	--10047
		x"27",	--10048
		x"2b",	--10049
		x"81",	--10050
		x"1e",	--10051
		x"d1",	--10052
		x"2b",	--10053
		x"0b",	--10054
		x"02",	--10055
		x"c1",	--10056
		x"2b",	--10057
		x"0b",	--10058
		x"0b",	--10059
		x"0b",	--10060
		x"c1",	--10061
		x"2f",	--10062
		x"05",	--10063
		x"f1",	--10064
		x"00",	--10065
		x"12",	--10066
		x"c1",	--10067
		x"2b",	--10068
		x"0f",	--10069
		x"68",	--10070
		x"b1",	--10071
		x"10",	--10072
		x"28",	--10073
		x"03",	--10074
		x"78",	--10075
		x"40",	--10076
		x"05",	--10077
		x"b1",	--10078
		x"28",	--10079
		x"04",	--10080
		x"78",	--10081
		x"20",	--10082
		x"c1",	--10083
		x"00",	--10084
		x"68",	--10085
		x"68",	--10086
		x"30",	--10087
		x"c1",	--10088
		x"2f",	--10089
		x"2d",	--10090
		x"f1",	--10091
		x"2d",	--10092
		x"02",	--10093
		x"68",	--10094
		x"11",	--10095
		x"b1",	--10096
		x"1e",	--10097
		x"b1",	--10098
		x"20",	--10099
		x"b1",	--10100
		x"22",	--10101
		x"b1",	--10102
		x"24",	--10103
		x"91",	--10104
		x"1e",	--10105
		x"81",	--10106
		x"20",	--10107
		x"81",	--10108
		x"22",	--10109
		x"81",	--10110
		x"24",	--10111
		x"17",	--10112
		x"58",	--10113
		x"0f",	--10114
		x"1a",	--10115
		x"1e",	--10116
		x"1b",	--10117
		x"20",	--10118
		x"3a",	--10119
		x"3b",	--10120
		x"0e",	--10121
		x"0f",	--10122
		x"1e",	--10123
		x"0f",	--10124
		x"81",	--10125
		x"1e",	--10126
		x"81",	--10127
		x"20",	--10128
		x"06",	--10129
		x"1a",	--10130
		x"1e",	--10131
		x"3a",	--10132
		x"1a",	--10133
		x"81",	--10134
		x"1e",	--10135
		x"c1",	--10136
		x"1b",	--10137
		x"68",	--10138
		x"6a",	--10139
		x"16",	--10140
		x"1e",	--10141
		x"91",	--10142
		x"20",	--10143
		x"3c",	--10144
		x"18",	--10145
		x"22",	--10146
		x"14",	--10147
		x"24",	--10148
		x"07",	--10149
		x"37",	--10150
		x"1a",	--10151
		x"09",	--10152
		x"91",	--10153
		x"28",	--10154
		x"32",	--10155
		x"1b",	--10156
		x"28",	--10157
		x"8b",	--10158
		x"8b",	--10159
		x"8b",	--10160
		x"8b",	--10161
		x"81",	--10162
		x"34",	--10163
		x"81",	--10164
		x"36",	--10165
		x"81",	--10166
		x"38",	--10167
		x"11",	--10168
		x"3a",	--10169
		x"11",	--10170
		x"3a",	--10171
		x"11",	--10172
		x"3a",	--10173
		x"11",	--10174
		x"3a",	--10175
		x"0c",	--10176
		x"1d",	--10177
		x"44",	--10178
		x"0e",	--10179
		x"0f",	--10180
		x"b0",	--10181
		x"44",	--10182
		x"31",	--10183
		x"0b",	--10184
		x"3c",	--10185
		x"0a",	--10186
		x"05",	--10187
		x"7b",	--10188
		x"30",	--10189
		x"c7",	--10190
		x"00",	--10191
		x"0c",	--10192
		x"4b",	--10193
		x"d1",	--10194
		x"01",	--10195
		x"03",	--10196
		x"7a",	--10197
		x"37",	--10198
		x"02",	--10199
		x"7a",	--10200
		x"57",	--10201
		x"4a",	--10202
		x"c7",	--10203
		x"00",	--10204
		x"06",	--10205
		x"36",	--10206
		x"11",	--10207
		x"3a",	--10208
		x"11",	--10209
		x"3a",	--10210
		x"11",	--10211
		x"3a",	--10212
		x"11",	--10213
		x"3a",	--10214
		x"0c",	--10215
		x"1d",	--10216
		x"44",	--10217
		x"0e",	--10218
		x"0f",	--10219
		x"b0",	--10220
		x"1e",	--10221
		x"31",	--10222
		x"09",	--10223
		x"81",	--10224
		x"3c",	--10225
		x"08",	--10226
		x"04",	--10227
		x"37",	--10228
		x"0c",	--10229
		x"b2",	--10230
		x"0d",	--10231
		x"b0",	--10232
		x"0e",	--10233
		x"ae",	--10234
		x"0f",	--10235
		x"ac",	--10236
		x"81",	--10237
		x"1e",	--10238
		x"81",	--10239
		x"20",	--10240
		x"81",	--10241
		x"22",	--10242
		x"81",	--10243
		x"24",	--10244
		x"6c",	--10245
		x"58",	--10246
		x"3e",	--10247
		x"14",	--10248
		x"1e",	--10249
		x"17",	--10250
		x"20",	--10251
		x"08",	--10252
		x"38",	--10253
		x"1a",	--10254
		x"19",	--10255
		x"28",	--10256
		x"89",	--10257
		x"89",	--10258
		x"89",	--10259
		x"89",	--10260
		x"1c",	--10261
		x"28",	--10262
		x"0d",	--10263
		x"0e",	--10264
		x"0f",	--10265
		x"b0",	--10266
		x"48",	--10267
		x"0b",	--10268
		x"3e",	--10269
		x"0a",	--10270
		x"05",	--10271
		x"7b",	--10272
		x"30",	--10273
		x"c8",	--10274
		x"00",	--10275
		x"0c",	--10276
		x"4b",	--10277
		x"d1",	--10278
		x"01",	--10279
		x"03",	--10280
		x"7a",	--10281
		x"37",	--10282
		x"02",	--10283
		x"7a",	--10284
		x"57",	--10285
		x"4a",	--10286
		x"c8",	--10287
		x"00",	--10288
		x"06",	--10289
		x"36",	--10290
		x"1c",	--10291
		x"28",	--10292
		x"0d",	--10293
		x"0e",	--10294
		x"0f",	--10295
		x"b0",	--10296
		x"12",	--10297
		x"04",	--10298
		x"07",	--10299
		x"38",	--10300
		x"0e",	--10301
		x"d0",	--10302
		x"0f",	--10303
		x"ce",	--10304
		x"81",	--10305
		x"1e",	--10306
		x"81",	--10307
		x"20",	--10308
		x"2c",	--10309
		x"17",	--10310
		x"1e",	--10311
		x"08",	--10312
		x"38",	--10313
		x"1a",	--10314
		x"1e",	--10315
		x"28",	--10316
		x"0f",	--10317
		x"b0",	--10318
		x"b8",	--10319
		x"0d",	--10320
		x"3f",	--10321
		x"0a",	--10322
		x"05",	--10323
		x"7d",	--10324
		x"30",	--10325
		x"c8",	--10326
		x"00",	--10327
		x"0c",	--10328
		x"4d",	--10329
		x"d1",	--10330
		x"01",	--10331
		x"03",	--10332
		x"7c",	--10333
		x"37",	--10334
		x"02",	--10335
		x"7c",	--10336
		x"57",	--10337
		x"4c",	--10338
		x"c8",	--10339
		x"00",	--10340
		x"06",	--10341
		x"36",	--10342
		x"1e",	--10343
		x"28",	--10344
		x"0f",	--10345
		x"b0",	--10346
		x"9e",	--10347
		x"07",	--10348
		x"38",	--10349
		x"0f",	--10350
		x"db",	--10351
		x"81",	--10352
		x"1e",	--10353
		x"b1",	--10354
		x"0a",	--10355
		x"28",	--10356
		x"02",	--10357
		x"c1",	--10358
		x"02",	--10359
		x"c1",	--10360
		x"2e",	--10361
		x"2a",	--10362
		x"0f",	--10363
		x"3f",	--10364
		x"1c",	--10365
		x"81",	--10366
		x"42",	--10367
		x"1a",	--10368
		x"1c",	--10369
		x"8a",	--10370
		x"8a",	--10371
		x"8a",	--10372
		x"8a",	--10373
		x"81",	--10374
		x"44",	--10375
		x"81",	--10376
		x"46",	--10377
		x"0a",	--10378
		x"8a",	--10379
		x"8a",	--10380
		x"8a",	--10381
		x"8a",	--10382
		x"81",	--10383
		x"48",	--10384
		x"1c",	--10385
		x"42",	--10386
		x"1d",	--10387
		x"44",	--10388
		x"1c",	--10389
		x"46",	--10390
		x"1d",	--10391
		x"48",	--10392
		x"2c",	--10393
		x"1c",	--10394
		x"26",	--10395
		x"0e",	--10396
		x"e1",	--10397
		x"01",	--10398
		x"5e",	--10399
		x"26",	--10400
		x"4e",	--10401
		x"c1",	--10402
		x"03",	--10403
		x"06",	--10404
		x"c1",	--10405
		x"2a",	--10406
		x"03",	--10407
		x"91",	--10408
		x"26",	--10409
		x"30",	--10410
		x"11",	--10411
		x"04",	--10412
		x"11",	--10413
		x"04",	--10414
		x"1d",	--10415
		x"34",	--10416
		x"0e",	--10417
		x"1e",	--10418
		x"1f",	--10419
		x"3e",	--10420
		x"b0",	--10421
		x"a2",	--10422
		x"21",	--10423
		x"81",	--10424
		x"2c",	--10425
		x"0d",	--10426
		x"7f",	--10427
		x"8f",	--10428
		x"91",	--10429
		x"3c",	--10430
		x"0e",	--10431
		x"0e",	--10432
		x"19",	--10433
		x"40",	--10434
		x"f7",	--10435
		x"81",	--10436
		x"3e",	--10437
		x"81",	--10438
		x"2c",	--10439
		x"07",	--10440
		x"0e",	--10441
		x"91",	--10442
		x"26",	--10443
		x"30",	--10444
		x"d1",	--10445
		x"2e",	--10446
		x"c1",	--10447
		x"2a",	--10448
		x"03",	--10449
		x"05",	--10450
		x"d1",	--10451
		x"2a",	--10452
		x"81",	--10453
		x"26",	--10454
		x"17",	--10455
		x"16",	--10456
		x"40",	--10457
		x"6e",	--10458
		x"4e",	--10459
		x"02",	--10460
		x"30",	--10461
		x"86",	--10462
		x"1f",	--10463
		x"2c",	--10464
		x"31",	--10465
		x"4a",	--10466
		x"34",	--10467
		x"35",	--10468
		x"36",	--10469
		x"37",	--10470
		x"38",	--10471
		x"39",	--10472
		x"3a",	--10473
		x"3b",	--10474
		x"30",	--10475
		x"0d",	--10476
		x"0f",	--10477
		x"04",	--10478
		x"3d",	--10479
		x"03",	--10480
		x"3f",	--10481
		x"1f",	--10482
		x"0e",	--10483
		x"03",	--10484
		x"5d",	--10485
		x"3e",	--10486
		x"1e",	--10487
		x"0d",	--10488
		x"b0",	--10489
		x"9e",	--10490
		x"3d",	--10491
		x"6d",	--10492
		x"02",	--10493
		x"3e",	--10494
		x"1e",	--10495
		x"5d",	--10496
		x"02",	--10497
		x"3f",	--10498
		x"1f",	--10499
		x"30",	--10500
		x"b0",	--10501
		x"d8",	--10502
		x"0f",	--10503
		x"30",	--10504
		x"0b",	--10505
		x"0a",	--10506
		x"09",	--10507
		x"79",	--10508
		x"20",	--10509
		x"0a",	--10510
		x"0b",	--10511
		x"0c",	--10512
		x"0d",	--10513
		x"0e",	--10514
		x"0f",	--10515
		x"0c",	--10516
		x"0d",	--10517
		x"0d",	--10518
		x"06",	--10519
		x"02",	--10520
		x"0c",	--10521
		x"03",	--10522
		x"0c",	--10523
		x"0d",	--10524
		x"1e",	--10525
		x"19",	--10526
		x"f2",	--10527
		x"39",	--10528
		x"3a",	--10529
		x"3b",	--10530
		x"30",	--10531
		x"b0",	--10532
		x"12",	--10533
		x"0e",	--10534
		x"0f",	--10535
		x"30",	--10536
		x"0b",	--10537
		x"0b",	--10538
		x"0f",	--10539
		x"06",	--10540
		x"3b",	--10541
		x"03",	--10542
		x"3e",	--10543
		x"3f",	--10544
		x"1e",	--10545
		x"0f",	--10546
		x"0d",	--10547
		x"05",	--10548
		x"5b",	--10549
		x"3c",	--10550
		x"3d",	--10551
		x"1c",	--10552
		x"0d",	--10553
		x"b0",	--10554
		x"12",	--10555
		x"6b",	--10556
		x"04",	--10557
		x"3c",	--10558
		x"3d",	--10559
		x"1c",	--10560
		x"0d",	--10561
		x"5b",	--10562
		x"04",	--10563
		x"3e",	--10564
		x"3f",	--10565
		x"1e",	--10566
		x"0f",	--10567
		x"3b",	--10568
		x"30",	--10569
		x"b0",	--10570
		x"52",	--10571
		x"0e",	--10572
		x"0f",	--10573
		x"30",	--10574
		x"7c",	--10575
		x"10",	--10576
		x"0d",	--10577
		x"0e",	--10578
		x"0f",	--10579
		x"0e",	--10580
		x"0e",	--10581
		x"02",	--10582
		x"0e",	--10583
		x"1f",	--10584
		x"1c",	--10585
		x"f8",	--10586
		x"30",	--10587
		x"b0",	--10588
		x"9e",	--10589
		x"0f",	--10590
		x"30",	--10591
		x"07",	--10592
		x"06",	--10593
		x"05",	--10594
		x"04",	--10595
		x"30",	--10596
		x"40",	--10597
		x"04",	--10598
		x"05",	--10599
		x"06",	--10600
		x"07",	--10601
		x"08",	--10602
		x"09",	--10603
		x"0a",	--10604
		x"0b",	--10605
		x"0c",	--10606
		x"0d",	--10607
		x"0e",	--10608
		x"0f",	--10609
		x"08",	--10610
		x"09",	--10611
		x"0a",	--10612
		x"0b",	--10613
		x"0b",	--10614
		x"0e",	--10615
		x"08",	--10616
		x"0a",	--10617
		x"0b",	--10618
		x"05",	--10619
		x"09",	--10620
		x"08",	--10621
		x"02",	--10622
		x"08",	--10623
		x"05",	--10624
		x"08",	--10625
		x"09",	--10626
		x"0a",	--10627
		x"0b",	--10628
		x"1c",	--10629
		x"91",	--10630
		x"00",	--10631
		x"e5",	--10632
		x"21",	--10633
		x"34",	--10634
		x"35",	--10635
		x"36",	--10636
		x"37",	--10637
		x"30",	--10638
		x"0b",	--10639
		x"0a",	--10640
		x"09",	--10641
		x"08",	--10642
		x"18",	--10643
		x"0a",	--10644
		x"19",	--10645
		x"0c",	--10646
		x"1a",	--10647
		x"0e",	--10648
		x"1b",	--10649
		x"10",	--10650
		x"b0",	--10651
		x"c0",	--10652
		x"38",	--10653
		x"39",	--10654
		x"3a",	--10655
		x"3b",	--10656
		x"30",	--10657
		x"0b",	--10658
		x"0a",	--10659
		x"09",	--10660
		x"08",	--10661
		x"18",	--10662
		x"0a",	--10663
		x"19",	--10664
		x"0c",	--10665
		x"1a",	--10666
		x"0e",	--10667
		x"1b",	--10668
		x"10",	--10669
		x"b0",	--10670
		x"c0",	--10671
		x"0c",	--10672
		x"0d",	--10673
		x"0e",	--10674
		x"0f",	--10675
		x"38",	--10676
		x"39",	--10677
		x"3a",	--10678
		x"3b",	--10679
		x"30",	--10680
		x"0b",	--10681
		x"0a",	--10682
		x"09",	--10683
		x"08",	--10684
		x"07",	--10685
		x"18",	--10686
		x"0c",	--10687
		x"19",	--10688
		x"0e",	--10689
		x"1a",	--10690
		x"10",	--10691
		x"1b",	--10692
		x"12",	--10693
		x"b0",	--10694
		x"c0",	--10695
		x"17",	--10696
		x"14",	--10697
		x"87",	--10698
		x"00",	--10699
		x"87",	--10700
		x"02",	--10701
		x"87",	--10702
		x"04",	--10703
		x"87",	--10704
		x"06",	--10705
		x"37",	--10706
		x"38",	--10707
		x"39",	--10708
		x"3a",	--10709
		x"3b",	--10710
		x"30",	--10711
		x"00",	--10712
		x"32",	--10713
		x"f0",	--10714
		x"fd",	--10715
		x"78",	--10716
		x"25",	--10717
		x"20",	--10718
		x"3d",	--10719
		x"64",	--10720
		x"74",	--10721
		x"25",	--10722
		x"00",	--10723
		x"73",	--10724
		x"0a",	--10725
		x"25",	--10726
		x"20",	--10727
		x"0d",	--10728
		x"00",	--10729
		x"ae",	--10730
		x"d6",	--10731
		x"dc",	--10732
		x"e4",	--10733
		x"ec",	--10734
		x"f4",	--10735
		x"c6",	--10736
		x"ce",	--10737
		x"0d",	--10738
		x"3d",	--10739
		x"3d",	--10740
		x"3d",	--10741
		x"20",	--10742
		x"61",	--10743
		x"63",	--10744
		x"6c",	--10745
		x"4d",	--10746
		x"55",	--10747
		x"3d",	--10748
		x"3d",	--10749
		x"3d",	--10750
		x"0d",	--10751
		x"00",	--10752
		x"6e",	--10753
		x"65",	--10754
		x"61",	--10755
		x"74",	--10756
		x"76",	--10757
		x"20",	--10758
		x"6f",	--10759
		x"65",	--10760
		x"77",	--10761
		x"69",	--10762
		x"65",	--10763
		x"72",	--10764
		x"61",	--10765
		x"00",	--10766
		x"75",	--10767
		x"7a",	--10768
		x"72",	--10769
		x"70",	--10770
		x"6d",	--10771
		x"65",	--10772
		x"63",	--10773
		x"64",	--10774
		x"72",	--10775
		x"73",	--10776
		x"65",	--10777
		x"64",	--10778
		x"63",	--10779
		x"6e",	--10780
		x"72",	--10781
		x"6c",	--10782
		x"65",	--10783
		x"00",	--10784
		x"64",	--10785
		x"6d",	--10786
		x"74",	--10787
		x"79",	--10788
		x"73",	--10789
		x"65",	--10790
		x"64",	--10791
		x"63",	--10792
		x"6e",	--10793
		x"69",	--10794
		x"75",	--10795
		x"61",	--10796
		x"69",	--10797
		x"6e",	--10798
		x"6f",	--10799
		x"73",	--10800
		x"61",	--10801
		x"6c",	--10802
		x"20",	--10803
		x"76",	--10804
		x"69",	--10805
		x"61",	--10806
		x"63",	--10807
		x"00",	--10808
		x"6f",	--10809
		x"6d",	--10810
		x"62",	--10811
		x"6f",	--10812
		x"6c",	--10813
		x"61",	--10814
		x"65",	--10815
		x"00",	--10816
		x"0a",	--10817
		x"08",	--10818
		x"08",	--10819
		x"25",	--10820
		x"00",	--10821
		x"50",	--10822
		x"0a",	--10823
		x"44",	--10824
		x"57",	--10825
		x"0d",	--10826
		x"00",	--10827
		x"49",	--10828
		x"48",	--10829
		x"0d",	--10830
		x"00",	--10831
		x"45",	--10832
		x"54",	--10833
		x"0a",	--10834
		x"53",	--10835
		x"6f",	--10836
		x"0d",	--10837
		x"00",	--10838
		x"6f",	--10839
		x"72",	--10840
		x"63",	--10841
		x"20",	--10842
		x"73",	--10843
		x"67",	--10844
		x"3a",	--10845
		x"0a",	--10846
		x"09",	--10847
		x"63",	--10848
		x"5b",	--10849
		x"5d",	--10850
		x"4c",	--10851
		x"46",	--10852
		x"20",	--10853
		x"49",	--10854
		x"48",	--10855
		x"20",	--10856
		x"54",	--10857
		x"4d",	--10858
		x"4f",	--10859
		x"54",	--10860
		x"0d",	--10861
		x"00",	--10862
		x"64",	--10863
		x"25",	--10864
		x"0d",	--10865
		x"00",	--10866
		x"6f",	--10867
		x"20",	--10868
		x"6d",	--10869
		x"6c",	--10870
		x"6d",	--10871
		x"6e",	--10872
		x"65",	--10873
		x"20",	--10874
		x"65",	--10875
		x"0d",	--10876
		x"00",	--10877
		x"61",	--10878
		x"74",	--10879
		x"6e",	--10880
		x"20",	--10881
		x"6f",	--10882
		x"20",	--10883
		x"20",	--10884
		x"65",	--10885
		x"20",	--10886
		x"62",	--10887
		x"6e",	--10888
		x"66",	--10889
		x"6c",	--10890
		x"0d",	--10891
		x"00",	--10892
		x"65",	--10893
		x"73",	--10894
		x"6f",	--10895
		x"6c",	--10896
		x"20",	--10897
		x"6f",	--10898
		x"20",	--10899
		x"65",	--10900
		x"20",	--10901
		x"68",	--10902
		x"74",	--10903
		x"0a",	--10904
		x"25",	--10905
		x"20",	--10906
		x"73",	--10907
		x"6e",	--10908
		x"74",	--10909
		x"61",	--10910
		x"6e",	--10911
		x"6d",	--10912
		x"65",	--10913
		x"0d",	--10914
		x"00",	--10915
		x"74",	--10916
		x"70",	--10917
		x"0a",	--10918
		x"65",	--10919
		x"72",	--10920
		x"72",	--10921
		x"20",	--10922
		x"69",	--10923
		x"73",	--10924
		x"6e",	--10925
		x"20",	--10926
		x"72",	--10927
		x"75",	--10928
		x"65",	--10929
		x"74",	--10930
		x"0a",	--10931
		x"63",	--10932
		x"72",	--10933
		x"65",	--10934
		x"74",	--10935
		x"75",	--10936
		x"61",	--10937
		x"65",	--10938
		x"0d",	--10939
		x"00",	--10940
		x"25",	--10941
		x"20",	--10942
		x"45",	--10943
		x"54",	--10944
		x"52",	--10945
		x"47",	--10946
		x"54",	--10947
		x"3c",	--10948
		x"49",	--10949
		x"45",	--10950
		x"55",	--10951
		x"3e",	--10952
		x"0a",	--10953
		x"25",	--10954
		x"20",	--10955
		x"64",	--10956
		x"0a",	--10957
		x"25",	--10958
		x"64",	--10959
		x"25",	--10960
		x"64",	--10961
		x"25",	--10962
		x"0d",	--10963
		x"00",	--10964
		x"64",	--10965
		x"25",	--10966
		x"0d",	--10967
		x"00",	--10968
		x"64",	--10969
		x"00",	--10970
		x"0a",	--10971
		x"59",	--10972
		x"20",	--10973
		x"65",	--10974
		x"69",	--10975
		x"64",	--10976
		x"6d",	--10977
		x"20",	--10978
		x"75",	--10979
		x"20",	--10980
		x"20",	--10981
		x"6f",	--10982
		x"27",	--10983
		x"20",	--10984
		x"69",	--10985
		x"65",	--10986
		x"61",	--10987
		x"73",	--10988
		x"69",	--10989
		x"21",	--10990
		x"0a",	--10991
		x"59",	--10992
		x"20",	--10993
		x"6e",	--10994
		x"66",	--10995
		x"6f",	--10996
		x"74",	--10997
		x"0a",	--10998
		x"59",	--10999
		x"20",	--11000
		x"6e",	--11001
		x"74",	--11002
		x"65",	--11003
		x"72",	--11004
		x"67",	--11005
		x"74",	--11006
		x"0a",	--11007
		x"59",	--11008
		x"20",	--11009
		x"6e",	--11010
		x"74",	--11011
		x"65",	--11012
		x"6c",	--11013
		x"66",	--11014
		x"0d",	--11015
		x"00",	--11016
		x"64",	--11017
		x"0a",	--11018
		x"73",	--11019
		x"6f",	--11020
		x"0d",	--11021
		x"00",	--11022
		x"72",	--11023
		x"6e",	--11024
		x"3a",	--11025
		x"6f",	--11026
		x"61",	--11027
		x"69",	--11028
		x"6e",	--11029
		x"0a",	--11030
		x"6c",	--11031
		x"66",	--11032
		x"3a",	--11033
		x"6f",	--11034
		x"61",	--11035
		x"69",	--11036
		x"6e",	--11037
		x"0a",	--11038
		x"72",	--11039
		x"67",	--11040
		x"74",	--11041
		x"72",	--11042
		x"74",	--11043
		x"74",	--11044
		x"6f",	--11045
		x"0d",	--11046
		x"00",	--11047
		x"6f",	--11048
		x"6d",	--11049
		x"6e",	--11050
		x"20",	--11051
		x"63",	--11052
		x"69",	--11053
		x"61",	--11054
		x"65",	--11055
		x"0d",	--11056
		x"00",	--11057
		x"6f",	--11058
		x"6d",	--11059
		x"6e",	--11060
		x"20",	--11061
		x"65",	--11062
		x"63",	--11063
		x"69",	--11064
		x"61",	--11065
		x"65",	--11066
		x"0d",	--11067
		x"00",	--11068
		x"72",	--11069
		x"74",	--11070
		x"0a",	--11071
		x"00",	--11072
		x"72",	--11073
		x"6f",	--11074
		x"3a",	--11075
		x"6d",	--11076
		x"73",	--11077
		x"69",	--11078
		x"67",	--11079
		x"61",	--11080
		x"67",	--11081
		x"6d",	--11082
		x"6e",	--11083
		x"0d",	--11084
		x"00",	--11085
		x"6f",	--11086
		x"72",	--11087
		x"63",	--11088
		x"20",	--11089
		x"73",	--11090
		x"67",	--11091
		x"3a",	--11092
		x"0a",	--11093
		x"09",	--11094
		x"73",	--11095
		x"52",	--11096
		x"47",	--11097
		x"53",	--11098
		x"45",	--11099
		x"20",	--11100
		x"41",	--11101
		x"55",	--11102
		x"0d",	--11103
		x"00",	--11104
		x"3d",	--11105
		x"64",	--11106
		x"76",	--11107
		x"25",	--11108
		x"0d",	--11109
		x"00",	--11110
		x"25",	--11111
		x"20",	--11112
		x"45",	--11113
		x"49",	--11114
		x"54",	--11115
		x"52",	--11116
		x"0a",	--11117
		x"72",	--11118
		x"61",	--11119
		x"0a",	--11120
		x"00",	--11121
		x"63",	--11122
		x"25",	--11123
		x"0d",	--11124
		x"00",	--11125
		x"63",	--11126
		x"20",	--11127
		x"6f",	--11128
		x"73",	--11129
		x"63",	--11130
		x"20",	--11131
		x"6f",	--11132
		x"6d",	--11133
		x"6e",	--11134
		x"0d",	--11135
		x"00",	--11136
		x"82",	--11137
		x"b0",	--11138
		x"b0",	--11139
		x"b0",	--11140
		x"b0",	--11141
		x"b0",	--11142
		x"b0",	--11143
		x"b0",	--11144
		x"b0",	--11145
		x"b0",	--11146
		x"b0",	--11147
		x"b0",	--11148
		x"b0",	--11149
		x"b0",	--11150
		x"b0",	--11151
		x"b0",	--11152
		x"b0",	--11153
		x"b0",	--11154
		x"b0",	--11155
		x"b0",	--11156
		x"b0",	--11157
		x"b0",	--11158
		x"b0",	--11159
		x"b0",	--11160
		x"b0",	--11161
		x"b0",	--11162
		x"b0",	--11163
		x"b0",	--11164
		x"b0",	--11165
		x"74",	--11166
		x"b0",	--11167
		x"b0",	--11168
		x"b0",	--11169
		x"b0",	--11170
		x"b0",	--11171
		x"b0",	--11172
		x"b0",	--11173
		x"b0",	--11174
		x"b0",	--11175
		x"b0",	--11176
		x"b0",	--11177
		x"b0",	--11178
		x"b0",	--11179
		x"b0",	--11180
		x"b0",	--11181
		x"b0",	--11182
		x"b0",	--11183
		x"b0",	--11184
		x"b0",	--11185
		x"b0",	--11186
		x"b0",	--11187
		x"b0",	--11188
		x"b0",	--11189
		x"b0",	--11190
		x"b0",	--11191
		x"b0",	--11192
		x"b0",	--11193
		x"b0",	--11194
		x"b0",	--11195
		x"b0",	--11196
		x"b0",	--11197
		x"66",	--11198
		x"58",	--11199
		x"4a",	--11200
		x"b0",	--11201
		x"b0",	--11202
		x"b0",	--11203
		x"b0",	--11204
		x"b0",	--11205
		x"b0",	--11206
		x"b0",	--11207
		x"32",	--11208
		x"b0",	--11209
		x"20",	--11210
		x"b0",	--11211
		x"b0",	--11212
		x"b0",	--11213
		x"b0",	--11214
		x"04",	--11215
		x"b0",	--11216
		x"b0",	--11217
		x"b0",	--11218
		x"f6",	--11219
		x"e4",	--11220
		x"30",	--11221
		x"32",	--11222
		x"34",	--11223
		x"36",	--11224
		x"38",	--11225
		x"61",	--11226
		x"63",	--11227
		x"65",	--11228
		x"00",	--11229
		x"38",	--11230
		x"ed",	--11231
		x"da",	--11232
		x"49",	--11233
		x"5e",	--11234
		x"7b",	--11235
		x"da",	--11236
		x"c9",	--11237
		x"69",	--11238
		x"ac",	--11239
		x"68",	--11240
		x"22",	--11241
		x"b4",	--11242
		x"14",	--11243
		x"68",	--11244
		x"a2",	--11245
		x"00",	--11246
		x"c9",	--11247
		x"00",	--11248
		x"49",	--11249
		x"00",	--11250
		x"96",	--11251
		x"00",	--11252
		x"c9",	--11253
		x"00",	--11254
		x"fb",	--11255
		x"00",	--11256
		x"16",	--11257
		x"00",	--11258
		x"2f",	--11259
		x"00",	--11260
		x"49",	--11261
		x"00",	--11262
		x"62",	--11263
		x"00",	--11264
		x"7b",	--11265
		x"00",	--11266
		x"8a",	--11267
		x"00",	--11268
		x"96",	--11269
		x"00",	--11270
		x"a3",	--11271
		x"00",	--11272
		x"af",	--11273
		x"00",	--11274
		x"bc",	--11275
		x"00",	--11276
		x"c9",	--11277
		x"00",	--11278
		x"d5",	--11279
		x"00",	--11280
		x"e2",	--11281
		x"00",	--11282
		x"ee",	--11283
		x"00",	--11284
		x"fb",	--11285
		x"00",	--11286
		x"03",	--11287
		x"00",	--11288
		x"0a",	--11289
		x"00",	--11290
		x"10",	--11291
		x"00",	--11292
		x"16",	--11293
		x"00",	--11294
		x"1d",	--11295
		x"00",	--11296
		x"23",	--11297
		x"00",	--11298
		x"29",	--11299
		x"00",	--11300
		x"2f",	--11301
		x"00",	--11302
		x"36",	--11303
		x"00",	--11304
		x"3c",	--11305
		x"00",	--11306
		x"42",	--11307
		x"00",	--11308
		x"49",	--11309
		x"a2",	--11310
		x"00",	--11311
		x"f9",	--11312
		x"00",	--11313
		x"83",	--11314
		x"00",	--11315
		x"6e",	--11316
		x"00",	--11317
		x"4e",	--11318
		x"00",	--11319
		x"44",	--11320
		x"00",	--11321
		x"15",	--11322
		x"00",	--11323
		x"29",	--11324
		x"00",	--11325
		x"fc",	--11326
		x"00",	--11327
		x"27",	--11328
		x"00",	--11329
		x"57",	--11330
		x"00",	--11331
		x"d1",	--11332
		x"00",	--11333
		x"f5",	--11334
		x"00",	--11335
		x"34",	--11336
		x"00",	--11337
		x"dd",	--11338
		x"00",	--11339
		x"c0",	--11340
		x"00",	--11341
		x"db",	--11342
		x"00",	--11343
		x"62",	--11344
		x"00",	--11345
		x"95",	--11346
		x"00",	--11347
		x"99",	--11348
		x"00",	--11349
		x"3c",	--11350
		x"00",	--11351
		x"43",	--11352
		x"00",	--11353
		x"90",	--11354
		x"00",	--11355
		x"41",	--11356
		x"00",	--11357
		x"fe",	--11358
		x"00",	--11359
		x"51",	--11360
		x"00",	--11361
		x"63",	--11362
		x"00",	--11363
		x"ab",	--11364
		x"00",	--11365
		x"de",	--11366
		x"00",	--11367
		x"bb",	--11368
		x"00",	--11369
		x"c5",	--11370
		x"00",	--11371
		x"61",	--11372
		x"00",	--11373
		x"b7",	--11374
		x"00",	--11375
		x"24",	--11376
		x"00",	--11377
		x"6e",	--11378
		x"00",	--11379
		x"3a",	--11380
		x"00",	--11381
		x"42",	--11382
		x"00",	--11383
		x"4d",	--11384
		x"00",	--11385
		x"d2",	--11386
		x"00",	--11387
		x"e0",	--11388
		x"00",	--11389
		x"06",	--11390
		x"00",	--11391
		x"49",	--11392
		x"00",	--11393
		x"2e",	--11394
		x"00",	--11395
		x"ea",	--11396
		x"00",	--11397
		x"09",	--11398
		x"00",	--11399
		x"d1",	--11400
		x"00",	--11401
		x"92",	--11402
		x"00",	--11403
		x"1c",	--11404
		x"00",	--11405
		x"fe",	--11406
		x"00",	--11407
		x"1d",	--11408
		x"00",	--11409
		x"eb",	--11410
		x"00",	--11411
		x"1c",	--11412
		x"00",	--11413
		x"b1",	--11414
		x"00",	--11415
		x"29",	--11416
		x"00",	--11417
		x"a7",	--11418
		x"00",	--11419
		x"3e",	--11420
		x"00",	--11421
		x"e8",	--11422
		x"00",	--11423
		x"82",	--11424
		x"00",	--11425
		x"35",	--11426
		x"00",	--11427
		x"f5",	--11428
		x"00",	--11429
		x"2e",	--11430
		x"00",	--11431
		x"bb",	--11432
		x"00",	--11433
		x"44",	--11434
		x"00",	--11435
		x"84",	--11436
		x"00",	--11437
		x"e9",	--11438
		x"00",	--11439
		x"9c",	--11440
		x"00",	--11441
		x"70",	--11442
		x"00",	--11443
		x"26",	--11444
		x"00",	--11445
		x"b4",	--11446
		x"00",	--11447
		x"5f",	--11448
		x"00",	--11449
		x"7e",	--11450
		x"00",	--11451
		x"41",	--11452
		x"00",	--11453
		x"39",	--11454
		x"00",	--11455
		x"91",	--11456
		x"00",	--11457
		x"d6",	--11458
		x"00",	--11459
		x"39",	--11460
		x"00",	--11461
		x"83",	--11462
		x"00",	--11463
		x"53",	--11464
		x"00",	--11465
		x"39",	--11466
		x"00",	--11467
		x"f4",	--11468
		x"00",	--11469
		x"9c",	--11470
		x"00",	--11471
		x"84",	--11472
		x"00",	--11473
		x"5f",	--11474
		x"00",	--11475
		x"8b",	--11476
		x"00",	--11477
		x"bd",	--11478
		x"00",	--11479
		x"f9",	--11480
		x"00",	--11481
		x"28",	--11482
		x"00",	--11483
		x"3b",	--11484
		x"00",	--11485
		x"1f",	--11486
		x"00",	--11487
		x"f8",	--11488
		x"00",	--11489
		x"97",	--11490
		x"00",	--11491
		x"ff",	--11492
		x"00",	--11493
		x"de",	--11494
		x"00",	--11495
		x"05",	--11496
		x"00",	--11497
		x"98",	--11498
		x"00",	--11499
		x"0f",	--11500
		x"00",	--11501
		x"ef",	--11502
		x"00",	--11503
		x"2f",	--11504
		x"00",	--11505
		x"11",	--11506
		x"00",	--11507
		x"8b",	--11508
		x"00",	--11509
		x"5a",	--11510
		x"00",	--11511
		x"0a",	--11512
		x"00",	--11513
		x"6d",	--11514
		x"00",	--11515
		x"1f",	--11516
		x"00",	--11517
		x"6d",	--11518
		x"00",	--11519
		x"36",	--11520
		x"00",	--11521
		x"7e",	--11522
		x"00",	--11523
		x"cf",	--11524
		x"00",	--11525
		x"27",	--11526
		x"00",	--11527
		x"cb",	--11528
		x"00",	--11529
		x"09",	--11530
		x"00",	--11531
		x"b7",	--11532
		x"00",	--11533
		x"4f",	--11534
		x"00",	--11535
		x"46",	--11536
		x"00",	--11537
		x"3f",	--11538
		x"00",	--11539
		x"66",	--11540
		x"00",	--11541
		x"9e",	--11542
		x"00",	--11543
		x"5f",	--11544
		x"00",	--11545
		x"ea",	--11546
		x"00",	--11547
		x"2d",	--11548
		x"00",	--11549
		x"75",	--11550
		x"00",	--11551
		x"27",	--11552
		x"00",	--11553
		x"ba",	--11554
		x"00",	--11555
		x"c7",	--11556
		x"00",	--11557
		x"eb",	--11558
		x"00",	--11559
		x"e5",	--11560
		x"00",	--11561
		x"f1",	--11562
		x"00",	--11563
		x"7b",	--11564
		x"00",	--11565
		x"3d",	--11566
		x"00",	--11567
		x"07",	--11568
		x"00",	--11569
		x"39",	--11570
		x"00",	--11571
		x"f7",	--11572
		x"00",	--11573
		x"8a",	--11574
		x"00",	--11575
		x"52",	--11576
		x"00",	--11577
		x"92",	--11578
		x"00",	--11579
		x"ea",	--11580
		x"00",	--11581
		x"6b",	--11582
		x"00",	--11583
		x"fb",	--11584
		x"00",	--11585
		x"5f",	--11586
		x"00",	--11587
		x"b1",	--11588
		x"00",	--11589
		x"1f",	--11590
		x"00",	--11591
		x"8d",	--11592
		x"00",	--11593
		x"5d",	--11594
		x"00",	--11595
		x"08",	--11596
		x"00",	--11597
		x"56",	--11598
		x"00",	--11599
		x"03",	--11600
		x"00",	--11601
		x"30",	--11602
		x"00",	--11603
		x"46",	--11604
		x"00",	--11605
		x"fc",	--11606
		x"00",	--11607
		x"7b",	--11608
		x"00",	--11609
		x"6b",	--11610
		x"00",	--11611
		x"ab",	--11612
		x"00",	--11613
		x"f0",	--11614
		x"00",	--11615
		x"cf",	--11616
		x"00",	--11617
		x"bc",	--11618
		x"00",	--11619
		x"20",	--11620
		x"00",	--11621
		x"9a",	--11622
		x"00",	--11623
		x"f4",	--11624
		x"00",	--11625
		x"36",	--11626
		x"00",	--11627
		x"1d",	--11628
		x"00",	--11629
		x"a9",	--11630
		x"00",	--11631
		x"e3",	--11632
		x"00",	--11633
		x"91",	--11634
		x"00",	--11635
		x"61",	--11636
		x"00",	--11637
		x"5e",	--11638
		x"00",	--11639
		x"e6",	--11640
		x"00",	--11641
		x"1b",	--11642
		x"00",	--11643
		x"08",	--11644
		x"00",	--11645
		x"65",	--11646
		x"00",	--11647
		x"99",	--11648
		x"00",	--11649
		x"85",	--11650
		x"00",	--11651
		x"5f",	--11652
		x"00",	--11653
		x"14",	--11654
		x"00",	--11655
		x"a0",	--11656
		x"00",	--11657
		x"68",	--11658
		x"00",	--11659
		x"40",	--11660
		x"00",	--11661
		x"8d",	--11662
		x"00",	--11663
		x"ff",	--11664
		x"00",	--11665
		x"d8",	--11666
		x"00",	--11667
		x"80",	--11668
		x"00",	--11669
		x"4d",	--11670
		x"00",	--11671
		x"73",	--11672
		x"00",	--11673
		x"27",	--11674
		x"00",	--11675
		x"31",	--11676
		x"00",	--11677
		x"06",	--11678
		x"00",	--11679
		x"06",	--11680
		x"00",	--11681
		x"15",	--11682
		x"00",	--11683
		x"56",	--11684
		x"00",	--11685
		x"ca",	--11686
		x"00",	--11687
		x"73",	--11688
		x"00",	--11689
		x"a8",	--11690
		x"00",	--11691
		x"c9",	--11692
		x"00",	--11693
		x"60",	--11694
		x"00",	--11695
		x"e2",	--11696
		x"00",	--11697
		x"7b",	--11698
		x"00",	--11699
		x"c0",	--11700
		x"00",	--11701
		x"8c",	--11702
		x"00",	--11703
		x"6b",	--11704
		x"00",	--11705
		x"04",	--11706
		x"07",	--11707
		x"09",	--11708
		x"00",	--11709
		x"c9",	--11710
		x"00",	--11711
		x"f0",	--11712
		x"00",	--11713
		x"da",	--11714
		x"00",	--11715
		x"a2",	--11716
		x"00",	--11717
		x"84",	--11718
		x"00",	--11719
		x"50",	--11720
		x"00",	--11721
		x"c2",	--11722
		x"00",	--11723
		x"d0",	--11724
		x"00",	--11725
		x"c4",	--11726
		x"00",	--11727
		x"c6",	--11728
		x"00",	--11729
		x"44",	--11730
		x"00",	--11731
		x"00",	--11732
		x"00",	--11733
		x"00",	--11734
		x"00",	--11735
		x"02",	--11736
		x"03",	--11737
		x"03",	--11738
		x"04",	--11739
		x"04",	--11740
		x"04",	--11741
		x"04",	--11742
		x"05",	--11743
		x"05",	--11744
		x"05",	--11745
		x"05",	--11746
		x"05",	--11747
		x"05",	--11748
		x"05",	--11749
		x"05",	--11750
		x"06",	--11751
		x"06",	--11752
		x"06",	--11753
		x"06",	--11754
		x"06",	--11755
		x"06",	--11756
		x"06",	--11757
		x"06",	--11758
		x"06",	--11759
		x"06",	--11760
		x"06",	--11761
		x"06",	--11762
		x"06",	--11763
		x"06",	--11764
		x"06",	--11765
		x"06",	--11766
		x"07",	--11767
		x"07",	--11768
		x"07",	--11769
		x"07",	--11770
		x"07",	--11771
		x"07",	--11772
		x"07",	--11773
		x"07",	--11774
		x"07",	--11775
		x"07",	--11776
		x"07",	--11777
		x"07",	--11778
		x"07",	--11779
		x"07",	--11780
		x"07",	--11781
		x"07",	--11782
		x"07",	--11783
		x"07",	--11784
		x"07",	--11785
		x"07",	--11786
		x"07",	--11787
		x"07",	--11788
		x"07",	--11789
		x"07",	--11790
		x"07",	--11791
		x"07",	--11792
		x"07",	--11793
		x"07",	--11794
		x"07",	--11795
		x"07",	--11796
		x"07",	--11797
		x"07",	--11798
		x"08",	--11799
		x"08",	--11800
		x"08",	--11801
		x"08",	--11802
		x"08",	--11803
		x"08",	--11804
		x"08",	--11805
		x"08",	--11806
		x"08",	--11807
		x"08",	--11808
		x"08",	--11809
		x"08",	--11810
		x"08",	--11811
		x"08",	--11812
		x"08",	--11813
		x"08",	--11814
		x"08",	--11815
		x"08",	--11816
		x"08",	--11817
		x"08",	--11818
		x"08",	--11819
		x"08",	--11820
		x"08",	--11821
		x"08",	--11822
		x"08",	--11823
		x"08",	--11824
		x"08",	--11825
		x"08",	--11826
		x"08",	--11827
		x"08",	--11828
		x"08",	--11829
		x"08",	--11830
		x"08",	--11831
		x"08",	--11832
		x"08",	--11833
		x"08",	--11834
		x"08",	--11835
		x"08",	--11836
		x"08",	--11837
		x"08",	--11838
		x"08",	--11839
		x"08",	--11840
		x"08",	--11841
		x"08",	--11842
		x"08",	--11843
		x"08",	--11844
		x"08",	--11845
		x"08",	--11846
		x"08",	--11847
		x"08",	--11848
		x"08",	--11849
		x"08",	--11850
		x"08",	--11851
		x"08",	--11852
		x"08",	--11853
		x"08",	--11854
		x"08",	--11855
		x"08",	--11856
		x"08",	--11857
		x"08",	--11858
		x"08",	--11859
		x"08",	--11860
		x"08",	--11861
		x"08",	--11862
		x"28",	--11863
		x"75",	--11864
		x"6c",	--11865
		x"00",	--11866
		x"ff",	--11867
		x"ff",	--11868
		x"ff",	--11869
		x"ff",	--11870
		x"2c",	--11871
		x"2c",	--11872
		x"2c",	--11873
		x"2c",	--11874
		x"2c",	--11875
		x"68",	--11876
		x"6c",	--11877
		x"00",	--11878
		x"ff",	--11879
		x"ff",	--11880
		x"ff",	--11881
		x"ff",	--11882
		x"ff",	--11883
		x"ff",	--11884
		x"ff",	--11885
		x"ff",	--11886
		x"ff",	--11887
		x"ff",	--11888
		x"ff",	--11889
		x"ff",	--11890
		x"ff",	--11891
		x"ff",	--11892
		x"ff",	--11893
		x"ff",	--11894
		x"ff",	--11895
		x"ff",	--11896
		x"ff",	--11897
		x"ff",	--11898
		x"ff",	--11899
		x"ff",	--11900
		x"ff",	--11901
		x"ff",	--11902
		x"ff",	--11903
		x"ff",	--11904
		x"ff",	--11905
		x"ff",	--11906
		x"ff",	--11907
		x"ff",	--11908
		x"ff",	--11909
		x"ff",	--11910
		x"ff",	--11911
		x"ff",	--11912
		x"ff",	--11913
		x"ff",	--11914
		x"ff",	--11915
		x"ff",	--11916
		x"ff",	--11917
		x"ff",	--11918
		x"ff",	--11919
		x"ff",	--11920
		x"ff",	--11921
		x"ff",	--11922
		x"ff",	--11923
		x"ff",	--11924
		x"ff",	--11925
		x"ff",	--11926
		x"ff",	--11927
		x"ff",	--11928
		x"ff",	--11929
		x"ff",	--11930
		x"ff",	--11931
		x"ff",	--11932
		x"ff",	--11933
		x"ff",	--11934
		x"ff",	--11935
		x"ff",	--11936
		x"ff",	--11937
		x"ff",	--11938
		x"ff",	--11939
		x"ff",	--11940
		x"ff",	--11941
		x"ff",	--11942
		x"ff",	--11943
		x"ff",	--11944
		x"ff",	--11945
		x"ff",	--11946
		x"ff",	--11947
		x"ff",	--11948
		x"ff",	--11949
		x"ff",	--11950
		x"ff",	--11951
		x"ff",	--11952
		x"ff",	--11953
		x"ff",	--11954
		x"ff",	--11955
		x"ff",	--11956
		x"ff",	--11957
		x"ff",	--11958
		x"ff",	--11959
		x"ff",	--11960
		x"ff",	--11961
		x"ff",	--11962
		x"ff",	--11963
		x"ff",	--11964
		x"ff",	--11965
		x"ff",	--11966
		x"ff",	--11967
		x"ff",	--11968
		x"ff",	--11969
		x"ff",	--11970
		x"ff",	--11971
		x"ff",	--11972
		x"ff",	--11973
		x"ff",	--11974
		x"ff",	--11975
		x"ff",	--11976
		x"ff",	--11977
		x"ff",	--11978
		x"ff",	--11979
		x"ff",	--11980
		x"ff",	--11981
		x"ff",	--11982
		x"ff",	--11983
		x"ff",	--11984
		x"ff",	--11985
		x"ff",	--11986
		x"ff",	--11987
		x"ff",	--11988
		x"ff",	--11989
		x"ff",	--11990
		x"ff",	--11991
		x"ff",	--11992
		x"ff",	--11993
		x"ff",	--11994
		x"ff",	--11995
		x"ff",	--11996
		x"ff",	--11997
		x"ff",	--11998
		x"ff",	--11999
		x"ff",	--12000
		x"ff",	--12001
		x"ff",	--12002
		x"ff",	--12003
		x"ff",	--12004
		x"ff",	--12005
		x"ff",	--12006
		x"ff",	--12007
		x"ff",	--12008
		x"ff",	--12009
		x"ff",	--12010
		x"ff",	--12011
		x"ff",	--12012
		x"ff",	--12013
		x"ff",	--12014
		x"ff",	--12015
		x"ff",	--12016
		x"ff",	--12017
		x"ff",	--12018
		x"ff",	--12019
		x"ff",	--12020
		x"ff",	--12021
		x"ff",	--12022
		x"ff",	--12023
		x"ff",	--12024
		x"ff",	--12025
		x"ff",	--12026
		x"ff",	--12027
		x"ff",	--12028
		x"ff",	--12029
		x"ff",	--12030
		x"ff",	--12031
		x"ff",	--12032
		x"ff",	--12033
		x"ff",	--12034
		x"ff",	--12035
		x"ff",	--12036
		x"ff",	--12037
		x"ff",	--12038
		x"ff",	--12039
		x"ff",	--12040
		x"ff",	--12041
		x"ff",	--12042
		x"ff",	--12043
		x"ff",	--12044
		x"ff",	--12045
		x"ff",	--12046
		x"ff",	--12047
		x"ff",	--12048
		x"ff",	--12049
		x"ff",	--12050
		x"ff",	--12051
		x"ff",	--12052
		x"ff",	--12053
		x"ff",	--12054
		x"ff",	--12055
		x"ff",	--12056
		x"ff",	--12057
		x"ff",	--12058
		x"ff",	--12059
		x"ff",	--12060
		x"ff",	--12061
		x"ff",	--12062
		x"ff",	--12063
		x"ff",	--12064
		x"ff",	--12065
		x"ff",	--12066
		x"ff",	--12067
		x"ff",	--12068
		x"ff",	--12069
		x"ff",	--12070
		x"ff",	--12071
		x"ff",	--12072
		x"ff",	--12073
		x"ff",	--12074
		x"ff",	--12075
		x"ff",	--12076
		x"ff",	--12077
		x"ff",	--12078
		x"ff",	--12079
		x"ff",	--12080
		x"ff",	--12081
		x"ff",	--12082
		x"ff",	--12083
		x"ff",	--12084
		x"ff",	--12085
		x"ff",	--12086
		x"ff",	--12087
		x"ff",	--12088
		x"ff",	--12089
		x"ff",	--12090
		x"ff",	--12091
		x"ff",	--12092
		x"ff",	--12093
		x"ff",	--12094
		x"ff",	--12095
		x"ff",	--12096
		x"ff",	--12097
		x"ff",	--12098
		x"ff",	--12099
		x"ff",	--12100
		x"ff",	--12101
		x"ff",	--12102
		x"ff",	--12103
		x"ff",	--12104
		x"ff",	--12105
		x"ff",	--12106
		x"ff",	--12107
		x"ff",	--12108
		x"ff",	--12109
		x"ff",	--12110
		x"ff",	--12111
		x"ff",	--12112
		x"ff",	--12113
		x"ff",	--12114
		x"ff",	--12115
		x"ff",	--12116
		x"ff",	--12117
		x"ff",	--12118
		x"ff",	--12119
		x"ff",	--12120
		x"ff",	--12121
		x"ff",	--12122
		x"ff",	--12123
		x"ff",	--12124
		x"ff",	--12125
		x"ff",	--12126
		x"ff",	--12127
		x"ff",	--12128
		x"ff",	--12129
		x"ff",	--12130
		x"ff",	--12131
		x"ff",	--12132
		x"ff",	--12133
		x"ff",	--12134
		x"ff",	--12135
		x"ff",	--12136
		x"ff",	--12137
		x"ff",	--12138
		x"ff",	--12139
		x"ff",	--12140
		x"ff",	--12141
		x"ff",	--12142
		x"ff",	--12143
		x"ff",	--12144
		x"ff",	--12145
		x"ff",	--12146
		x"ff",	--12147
		x"ff",	--12148
		x"ff",	--12149
		x"ff",	--12150
		x"ff",	--12151
		x"ff",	--12152
		x"ff",	--12153
		x"ff",	--12154
		x"ff",	--12155
		x"ff",	--12156
		x"ff",	--12157
		x"ff",	--12158
		x"ff",	--12159
		x"ff",	--12160
		x"ff",	--12161
		x"ff",	--12162
		x"ff",	--12163
		x"ff",	--12164
		x"ff",	--12165
		x"ff",	--12166
		x"ff",	--12167
		x"ff",	--12168
		x"ff",	--12169
		x"ff",	--12170
		x"ff",	--12171
		x"ff",	--12172
		x"ff",	--12173
		x"ff",	--12174
		x"ff",	--12175
		x"ff",	--12176
		x"ff",	--12177
		x"ff",	--12178
		x"ff",	--12179
		x"ff",	--12180
		x"ff",	--12181
		x"ff",	--12182
		x"ff",	--12183
		x"ff",	--12184
		x"ff",	--12185
		x"ff",	--12186
		x"ff",	--12187
		x"ff",	--12188
		x"ff",	--12189
		x"ff",	--12190
		x"ff",	--12191
		x"ff",	--12192
		x"ff",	--12193
		x"ff",	--12194
		x"ff",	--12195
		x"ff",	--12196
		x"ff",	--12197
		x"ff",	--12198
		x"ff",	--12199
		x"ff",	--12200
		x"ff",	--12201
		x"ff",	--12202
		x"ff",	--12203
		x"ff",	--12204
		x"ff",	--12205
		x"ff",	--12206
		x"ff",	--12207
		x"ff",	--12208
		x"ff",	--12209
		x"ff",	--12210
		x"ff",	--12211
		x"ff",	--12212
		x"ff",	--12213
		x"ff",	--12214
		x"ff",	--12215
		x"ff",	--12216
		x"ff",	--12217
		x"ff",	--12218
		x"ff",	--12219
		x"ff",	--12220
		x"ff",	--12221
		x"ff",	--12222
		x"ff",	--12223
		x"ff",	--12224
		x"ff",	--12225
		x"ff",	--12226
		x"ff",	--12227
		x"ff",	--12228
		x"ff",	--12229
		x"ff",	--12230
		x"ff",	--12231
		x"ff",	--12232
		x"ff",	--12233
		x"ff",	--12234
		x"ff",	--12235
		x"ff",	--12236
		x"ff",	--12237
		x"ff",	--12238
		x"ff",	--12239
		x"ff",	--12240
		x"ff",	--12241
		x"ff",	--12242
		x"ff",	--12243
		x"ff",	--12244
		x"ff",	--12245
		x"ff",	--12246
		x"ff",	--12247
		x"ff",	--12248
		x"ff",	--12249
		x"ff",	--12250
		x"ff",	--12251
		x"ff",	--12252
		x"ff",	--12253
		x"ff",	--12254
		x"ff",	--12255
		x"ff",	--12256
		x"ff",	--12257
		x"ff",	--12258
		x"ff",	--12259
		x"ff",	--12260
		x"ff",	--12261
		x"ff",	--12262
		x"ff",	--12263
		x"ff",	--12264
		x"ff",	--12265
		x"ff",	--12266
		x"ff",	--12267
		x"ff",	--12268
		x"ff",	--12269
		x"ff",	--12270
		x"ff",	--12271
		x"ff",	--12272
		x"ff",	--12273
		x"ff",	--12274
		x"ff",	--12275
		x"ff",	--12276
		x"ff",	--12277
		x"ff",	--12278
		x"ff",	--12279
		x"ff",	--12280
		x"ff",	--12281
		x"ff",	--12282
		x"ff",	--12283
		x"ff",	--12284
		x"ff",	--12285
		x"ff",	--12286
		x"ff",	--12287
		x"ff",	--12288
		x"ff",	--12289
		x"ff",	--12290
		x"ff",	--12291
		x"ff",	--12292
		x"ff",	--12293
		x"ff",	--12294
		x"ff",	--12295
		x"ff",	--12296
		x"ff",	--12297
		x"ff",	--12298
		x"ff",	--12299
		x"ff",	--12300
		x"ff",	--12301
		x"ff",	--12302
		x"ff",	--12303
		x"ff",	--12304
		x"ff",	--12305
		x"ff",	--12306
		x"ff",	--12307
		x"ff",	--12308
		x"ff",	--12309
		x"ff",	--12310
		x"ff",	--12311
		x"ff",	--12312
		x"ff",	--12313
		x"ff",	--12314
		x"ff",	--12315
		x"ff",	--12316
		x"ff",	--12317
		x"ff",	--12318
		x"ff",	--12319
		x"ff",	--12320
		x"ff",	--12321
		x"ff",	--12322
		x"ff",	--12323
		x"ff",	--12324
		x"ff",	--12325
		x"ff",	--12326
		x"ff",	--12327
		x"ff",	--12328
		x"ff",	--12329
		x"ff",	--12330
		x"ff",	--12331
		x"ff",	--12332
		x"ff",	--12333
		x"ff",	--12334
		x"ff",	--12335
		x"ff",	--12336
		x"ff",	--12337
		x"ff",	--12338
		x"ff",	--12339
		x"ff",	--12340
		x"ff",	--12341
		x"ff",	--12342
		x"ff",	--12343
		x"ff",	--12344
		x"ff",	--12345
		x"ff",	--12346
		x"ff",	--12347
		x"ff",	--12348
		x"ff",	--12349
		x"ff",	--12350
		x"ff",	--12351
		x"ff",	--12352
		x"ff",	--12353
		x"ff",	--12354
		x"ff",	--12355
		x"ff",	--12356
		x"ff",	--12357
		x"ff",	--12358
		x"ff",	--12359
		x"ff",	--12360
		x"ff",	--12361
		x"ff",	--12362
		x"ff",	--12363
		x"ff",	--12364
		x"ff",	--12365
		x"ff",	--12366
		x"ff",	--12367
		x"ff",	--12368
		x"ff",	--12369
		x"ff",	--12370
		x"ff",	--12371
		x"ff",	--12372
		x"ff",	--12373
		x"ff",	--12374
		x"ff",	--12375
		x"ff",	--12376
		x"ff",	--12377
		x"ff",	--12378
		x"ff",	--12379
		x"ff",	--12380
		x"ff",	--12381
		x"ff",	--12382
		x"ff",	--12383
		x"ff",	--12384
		x"ff",	--12385
		x"ff",	--12386
		x"ff",	--12387
		x"ff",	--12388
		x"ff",	--12389
		x"ff",	--12390
		x"ff",	--12391
		x"ff",	--12392
		x"ff",	--12393
		x"ff",	--12394
		x"ff",	--12395
		x"ff",	--12396
		x"ff",	--12397
		x"ff",	--12398
		x"ff",	--12399
		x"ff",	--12400
		x"ff",	--12401
		x"ff",	--12402
		x"ff",	--12403
		x"ff",	--12404
		x"ff",	--12405
		x"ff",	--12406
		x"ff",	--12407
		x"ff",	--12408
		x"ff",	--12409
		x"ff",	--12410
		x"ff",	--12411
		x"ff",	--12412
		x"ff",	--12413
		x"ff",	--12414
		x"ff",	--12415
		x"ff",	--12416
		x"ff",	--12417
		x"ff",	--12418
		x"ff",	--12419
		x"ff",	--12420
		x"ff",	--12421
		x"ff",	--12422
		x"ff",	--12423
		x"ff",	--12424
		x"ff",	--12425
		x"ff",	--12426
		x"ff",	--12427
		x"ff",	--12428
		x"ff",	--12429
		x"ff",	--12430
		x"ff",	--12431
		x"ff",	--12432
		x"ff",	--12433
		x"ff",	--12434
		x"ff",	--12435
		x"ff",	--12436
		x"ff",	--12437
		x"ff",	--12438
		x"ff",	--12439
		x"ff",	--12440
		x"ff",	--12441
		x"ff",	--12442
		x"ff",	--12443
		x"ff",	--12444
		x"ff",	--12445
		x"ff",	--12446
		x"ff",	--12447
		x"ff",	--12448
		x"ff",	--12449
		x"ff",	--12450
		x"ff",	--12451
		x"ff",	--12452
		x"ff",	--12453
		x"ff",	--12454
		x"ff",	--12455
		x"ff",	--12456
		x"ff",	--12457
		x"ff",	--12458
		x"ff",	--12459
		x"ff",	--12460
		x"ff",	--12461
		x"ff",	--12462
		x"ff",	--12463
		x"ff",	--12464
		x"ff",	--12465
		x"ff",	--12466
		x"ff",	--12467
		x"ff",	--12468
		x"ff",	--12469
		x"ff",	--12470
		x"ff",	--12471
		x"ff",	--12472
		x"ff",	--12473
		x"ff",	--12474
		x"ff",	--12475
		x"ff",	--12476
		x"ff",	--12477
		x"ff",	--12478
		x"ff",	--12479
		x"ff",	--12480
		x"ff",	--12481
		x"ff",	--12482
		x"ff",	--12483
		x"ff",	--12484
		x"ff",	--12485
		x"ff",	--12486
		x"ff",	--12487
		x"ff",	--12488
		x"ff",	--12489
		x"ff",	--12490
		x"ff",	--12491
		x"ff",	--12492
		x"ff",	--12493
		x"ff",	--12494
		x"ff",	--12495
		x"ff",	--12496
		x"ff",	--12497
		x"ff",	--12498
		x"ff",	--12499
		x"ff",	--12500
		x"ff",	--12501
		x"ff",	--12502
		x"ff",	--12503
		x"ff",	--12504
		x"ff",	--12505
		x"ff",	--12506
		x"ff",	--12507
		x"ff",	--12508
		x"ff",	--12509
		x"ff",	--12510
		x"ff",	--12511
		x"ff",	--12512
		x"ff",	--12513
		x"ff",	--12514
		x"ff",	--12515
		x"ff",	--12516
		x"ff",	--12517
		x"ff",	--12518
		x"ff",	--12519
		x"ff",	--12520
		x"ff",	--12521
		x"ff",	--12522
		x"ff",	--12523
		x"ff",	--12524
		x"ff",	--12525
		x"ff",	--12526
		x"ff",	--12527
		x"ff",	--12528
		x"ff",	--12529
		x"ff",	--12530
		x"ff",	--12531
		x"ff",	--12532
		x"ff",	--12533
		x"ff",	--12534
		x"ff",	--12535
		x"ff",	--12536
		x"ff",	--12537
		x"ff",	--12538
		x"ff",	--12539
		x"ff",	--12540
		x"ff",	--12541
		x"ff",	--12542
		x"ff",	--12543
		x"ff",	--12544
		x"ff",	--12545
		x"ff",	--12546
		x"ff",	--12547
		x"ff",	--12548
		x"ff",	--12549
		x"ff",	--12550
		x"ff",	--12551
		x"ff",	--12552
		x"ff",	--12553
		x"ff",	--12554
		x"ff",	--12555
		x"ff",	--12556
		x"ff",	--12557
		x"ff",	--12558
		x"ff",	--12559
		x"ff",	--12560
		x"ff",	--12561
		x"ff",	--12562
		x"ff",	--12563
		x"ff",	--12564
		x"ff",	--12565
		x"ff",	--12566
		x"ff",	--12567
		x"ff",	--12568
		x"ff",	--12569
		x"ff",	--12570
		x"ff",	--12571
		x"ff",	--12572
		x"ff",	--12573
		x"ff",	--12574
		x"ff",	--12575
		x"ff",	--12576
		x"ff",	--12577
		x"ff",	--12578
		x"ff",	--12579
		x"ff",	--12580
		x"ff",	--12581
		x"ff",	--12582
		x"ff",	--12583
		x"ff",	--12584
		x"ff",	--12585
		x"ff",	--12586
		x"ff",	--12587
		x"ff",	--12588
		x"ff",	--12589
		x"ff",	--12590
		x"ff",	--12591
		x"ff",	--12592
		x"ff",	--12593
		x"ff",	--12594
		x"ff",	--12595
		x"ff",	--12596
		x"ff",	--12597
		x"ff",	--12598
		x"ff",	--12599
		x"ff",	--12600
		x"ff",	--12601
		x"ff",	--12602
		x"ff",	--12603
		x"ff",	--12604
		x"ff",	--12605
		x"ff",	--12606
		x"ff",	--12607
		x"ff",	--12608
		x"ff",	--12609
		x"ff",	--12610
		x"ff",	--12611
		x"ff",	--12612
		x"ff",	--12613
		x"ff",	--12614
		x"ff",	--12615
		x"ff",	--12616
		x"ff",	--12617
		x"ff",	--12618
		x"ff",	--12619
		x"ff",	--12620
		x"ff",	--12621
		x"ff",	--12622
		x"ff",	--12623
		x"ff",	--12624
		x"ff",	--12625
		x"ff",	--12626
		x"ff",	--12627
		x"ff",	--12628
		x"ff",	--12629
		x"ff",	--12630
		x"ff",	--12631
		x"ff",	--12632
		x"ff",	--12633
		x"ff",	--12634
		x"ff",	--12635
		x"ff",	--12636
		x"ff",	--12637
		x"ff",	--12638
		x"ff",	--12639
		x"ff",	--12640
		x"ff",	--12641
		x"ff",	--12642
		x"ff",	--12643
		x"ff",	--12644
		x"ff",	--12645
		x"ff",	--12646
		x"ff",	--12647
		x"ff",	--12648
		x"ff",	--12649
		x"ff",	--12650
		x"ff",	--12651
		x"ff",	--12652
		x"ff",	--12653
		x"ff",	--12654
		x"ff",	--12655
		x"ff",	--12656
		x"ff",	--12657
		x"ff",	--12658
		x"ff",	--12659
		x"ff",	--12660
		x"ff",	--12661
		x"ff",	--12662
		x"ff",	--12663
		x"ff",	--12664
		x"ff",	--12665
		x"ff",	--12666
		x"ff",	--12667
		x"ff",	--12668
		x"ff",	--12669
		x"ff",	--12670
		x"ff",	--12671
		x"ff",	--12672
		x"ff",	--12673
		x"ff",	--12674
		x"ff",	--12675
		x"ff",	--12676
		x"ff",	--12677
		x"ff",	--12678
		x"ff",	--12679
		x"ff",	--12680
		x"ff",	--12681
		x"ff",	--12682
		x"ff",	--12683
		x"ff",	--12684
		x"ff",	--12685
		x"ff",	--12686
		x"ff",	--12687
		x"ff",	--12688
		x"ff",	--12689
		x"ff",	--12690
		x"ff",	--12691
		x"ff",	--12692
		x"ff",	--12693
		x"ff",	--12694
		x"ff",	--12695
		x"ff",	--12696
		x"ff",	--12697
		x"ff",	--12698
		x"ff",	--12699
		x"ff",	--12700
		x"ff",	--12701
		x"ff",	--12702
		x"ff",	--12703
		x"ff",	--12704
		x"ff",	--12705
		x"ff",	--12706
		x"ff",	--12707
		x"ff",	--12708
		x"ff",	--12709
		x"ff",	--12710
		x"ff",	--12711
		x"ff",	--12712
		x"ff",	--12713
		x"ff",	--12714
		x"ff",	--12715
		x"ff",	--12716
		x"ff",	--12717
		x"ff",	--12718
		x"ff",	--12719
		x"ff",	--12720
		x"ff",	--12721
		x"ff",	--12722
		x"ff",	--12723
		x"ff",	--12724
		x"ff",	--12725
		x"ff",	--12726
		x"ff",	--12727
		x"ff",	--12728
		x"ff",	--12729
		x"ff",	--12730
		x"ff",	--12731
		x"ff",	--12732
		x"ff",	--12733
		x"ff",	--12734
		x"ff",	--12735
		x"ff",	--12736
		x"ff",	--12737
		x"ff",	--12738
		x"ff",	--12739
		x"ff",	--12740
		x"ff",	--12741
		x"ff",	--12742
		x"ff",	--12743
		x"ff",	--12744
		x"ff",	--12745
		x"ff",	--12746
		x"ff",	--12747
		x"ff",	--12748
		x"ff",	--12749
		x"ff",	--12750
		x"ff",	--12751
		x"ff",	--12752
		x"ff",	--12753
		x"ff",	--12754
		x"ff",	--12755
		x"ff",	--12756
		x"ff",	--12757
		x"ff",	--12758
		x"ff",	--12759
		x"ff",	--12760
		x"ff",	--12761
		x"ff",	--12762
		x"ff",	--12763
		x"ff",	--12764
		x"ff",	--12765
		x"ff",	--12766
		x"ff",	--12767
		x"ff",	--12768
		x"ff",	--12769
		x"ff",	--12770
		x"ff",	--12771
		x"ff",	--12772
		x"ff",	--12773
		x"ff",	--12774
		x"ff",	--12775
		x"ff",	--12776
		x"ff",	--12777
		x"ff",	--12778
		x"ff",	--12779
		x"ff",	--12780
		x"ff",	--12781
		x"ff",	--12782
		x"ff",	--12783
		x"ff",	--12784
		x"ff",	--12785
		x"ff",	--12786
		x"ff",	--12787
		x"ff",	--12788
		x"ff",	--12789
		x"ff",	--12790
		x"ff",	--12791
		x"ff",	--12792
		x"ff",	--12793
		x"ff",	--12794
		x"ff",	--12795
		x"ff",	--12796
		x"ff",	--12797
		x"ff",	--12798
		x"ff",	--12799
		x"ff",	--12800
		x"ff",	--12801
		x"ff",	--12802
		x"ff",	--12803
		x"ff",	--12804
		x"ff",	--12805
		x"ff",	--12806
		x"ff",	--12807
		x"ff",	--12808
		x"ff",	--12809
		x"ff",	--12810
		x"ff",	--12811
		x"ff",	--12812
		x"ff",	--12813
		x"ff",	--12814
		x"ff",	--12815
		x"ff",	--12816
		x"ff",	--12817
		x"ff",	--12818
		x"ff",	--12819
		x"ff",	--12820
		x"ff",	--12821
		x"ff",	--12822
		x"ff",	--12823
		x"ff",	--12824
		x"ff",	--12825
		x"ff",	--12826
		x"ff",	--12827
		x"ff",	--12828
		x"ff",	--12829
		x"ff",	--12830
		x"ff",	--12831
		x"ff",	--12832
		x"ff",	--12833
		x"ff",	--12834
		x"ff",	--12835
		x"ff",	--12836
		x"ff",	--12837
		x"ff",	--12838
		x"ff",	--12839
		x"ff",	--12840
		x"ff",	--12841
		x"ff",	--12842
		x"ff",	--12843
		x"ff",	--12844
		x"ff",	--12845
		x"ff",	--12846
		x"ff",	--12847
		x"ff",	--12848
		x"ff",	--12849
		x"ff",	--12850
		x"ff",	--12851
		x"ff",	--12852
		x"ff",	--12853
		x"ff",	--12854
		x"ff",	--12855
		x"ff",	--12856
		x"ff",	--12857
		x"ff",	--12858
		x"ff",	--12859
		x"ff",	--12860
		x"ff",	--12861
		x"ff",	--12862
		x"ff",	--12863
		x"ff",	--12864
		x"ff",	--12865
		x"ff",	--12866
		x"ff",	--12867
		x"ff",	--12868
		x"ff",	--12869
		x"ff",	--12870
		x"ff",	--12871
		x"ff",	--12872
		x"ff",	--12873
		x"ff",	--12874
		x"ff",	--12875
		x"ff",	--12876
		x"ff",	--12877
		x"ff",	--12878
		x"ff",	--12879
		x"ff",	--12880
		x"ff",	--12881
		x"ff",	--12882
		x"ff",	--12883
		x"ff",	--12884
		x"ff",	--12885
		x"ff",	--12886
		x"ff",	--12887
		x"ff",	--12888
		x"ff",	--12889
		x"ff",	--12890
		x"ff",	--12891
		x"ff",	--12892
		x"ff",	--12893
		x"ff",	--12894
		x"ff",	--12895
		x"ff",	--12896
		x"ff",	--12897
		x"ff",	--12898
		x"ff",	--12899
		x"ff",	--12900
		x"ff",	--12901
		x"ff",	--12902
		x"ff",	--12903
		x"ff",	--12904
		x"ff",	--12905
		x"ff",	--12906
		x"ff",	--12907
		x"ff",	--12908
		x"ff",	--12909
		x"ff",	--12910
		x"ff",	--12911
		x"ff",	--12912
		x"ff",	--12913
		x"ff",	--12914
		x"ff",	--12915
		x"ff",	--12916
		x"ff",	--12917
		x"ff",	--12918
		x"ff",	--12919
		x"ff",	--12920
		x"ff",	--12921
		x"ff",	--12922
		x"ff",	--12923
		x"ff",	--12924
		x"ff",	--12925
		x"ff",	--12926
		x"ff",	--12927
		x"ff",	--12928
		x"ff",	--12929
		x"ff",	--12930
		x"ff",	--12931
		x"ff",	--12932
		x"ff",	--12933
		x"ff",	--12934
		x"ff",	--12935
		x"ff",	--12936
		x"ff",	--12937
		x"ff",	--12938
		x"ff",	--12939
		x"ff",	--12940
		x"ff",	--12941
		x"ff",	--12942
		x"ff",	--12943
		x"ff",	--12944
		x"ff",	--12945
		x"ff",	--12946
		x"ff",	--12947
		x"ff",	--12948
		x"ff",	--12949
		x"ff",	--12950
		x"ff",	--12951
		x"ff",	--12952
		x"ff",	--12953
		x"ff",	--12954
		x"ff",	--12955
		x"ff",	--12956
		x"ff",	--12957
		x"ff",	--12958
		x"ff",	--12959
		x"ff",	--12960
		x"ff",	--12961
		x"ff",	--12962
		x"ff",	--12963
		x"ff",	--12964
		x"ff",	--12965
		x"ff",	--12966
		x"ff",	--12967
		x"ff",	--12968
		x"ff",	--12969
		x"ff",	--12970
		x"ff",	--12971
		x"ff",	--12972
		x"ff",	--12973
		x"ff",	--12974
		x"ff",	--12975
		x"ff",	--12976
		x"ff",	--12977
		x"ff",	--12978
		x"ff",	--12979
		x"ff",	--12980
		x"ff",	--12981
		x"ff",	--12982
		x"ff",	--12983
		x"ff",	--12984
		x"ff",	--12985
		x"ff",	--12986
		x"ff",	--12987
		x"ff",	--12988
		x"ff",	--12989
		x"ff",	--12990
		x"ff",	--12991
		x"ff",	--12992
		x"ff",	--12993
		x"ff",	--12994
		x"ff",	--12995
		x"ff",	--12996
		x"ff",	--12997
		x"ff",	--12998
		x"ff",	--12999
		x"ff",	--13000
		x"ff",	--13001
		x"ff",	--13002
		x"ff",	--13003
		x"ff",	--13004
		x"ff",	--13005
		x"ff",	--13006
		x"ff",	--13007
		x"ff",	--13008
		x"ff",	--13009
		x"ff",	--13010
		x"ff",	--13011
		x"ff",	--13012
		x"ff",	--13013
		x"ff",	--13014
		x"ff",	--13015
		x"ff",	--13016
		x"ff",	--13017
		x"ff",	--13018
		x"ff",	--13019
		x"ff",	--13020
		x"ff",	--13021
		x"ff",	--13022
		x"ff",	--13023
		x"ff",	--13024
		x"ff",	--13025
		x"ff",	--13026
		x"ff",	--13027
		x"ff",	--13028
		x"ff",	--13029
		x"ff",	--13030
		x"ff",	--13031
		x"ff",	--13032
		x"ff",	--13033
		x"ff",	--13034
		x"ff",	--13035
		x"ff",	--13036
		x"ff",	--13037
		x"ff",	--13038
		x"ff",	--13039
		x"ff",	--13040
		x"ff",	--13041
		x"ff",	--13042
		x"ff",	--13043
		x"ff",	--13044
		x"ff",	--13045
		x"ff",	--13046
		x"ff",	--13047
		x"ff",	--13048
		x"ff",	--13049
		x"ff",	--13050
		x"ff",	--13051
		x"ff",	--13052
		x"ff",	--13053
		x"ff",	--13054
		x"ff",	--13055
		x"ff",	--13056
		x"ff",	--13057
		x"ff",	--13058
		x"ff",	--13059
		x"ff",	--13060
		x"ff",	--13061
		x"ff",	--13062
		x"ff",	--13063
		x"ff",	--13064
		x"ff",	--13065
		x"ff",	--13066
		x"ff",	--13067
		x"ff",	--13068
		x"ff",	--13069
		x"ff",	--13070
		x"ff",	--13071
		x"ff",	--13072
		x"ff",	--13073
		x"ff",	--13074
		x"ff",	--13075
		x"ff",	--13076
		x"ff",	--13077
		x"ff",	--13078
		x"ff",	--13079
		x"ff",	--13080
		x"ff",	--13081
		x"ff",	--13082
		x"ff",	--13083
		x"ff",	--13084
		x"ff",	--13085
		x"ff",	--13086
		x"ff",	--13087
		x"ff",	--13088
		x"ff",	--13089
		x"ff",	--13090
		x"ff",	--13091
		x"ff",	--13092
		x"ff",	--13093
		x"ff",	--13094
		x"ff",	--13095
		x"ff",	--13096
		x"ff",	--13097
		x"ff",	--13098
		x"ff",	--13099
		x"ff",	--13100
		x"ff",	--13101
		x"ff",	--13102
		x"ff",	--13103
		x"ff",	--13104
		x"ff",	--13105
		x"ff",	--13106
		x"ff",	--13107
		x"ff",	--13108
		x"ff",	--13109
		x"ff",	--13110
		x"ff",	--13111
		x"ff",	--13112
		x"ff",	--13113
		x"ff",	--13114
		x"ff",	--13115
		x"ff",	--13116
		x"ff",	--13117
		x"ff",	--13118
		x"ff",	--13119
		x"ff",	--13120
		x"ff",	--13121
		x"ff",	--13122
		x"ff",	--13123
		x"ff",	--13124
		x"ff",	--13125
		x"ff",	--13126
		x"ff",	--13127
		x"ff",	--13128
		x"ff",	--13129
		x"ff",	--13130
		x"ff",	--13131
		x"ff",	--13132
		x"ff",	--13133
		x"ff",	--13134
		x"ff",	--13135
		x"ff",	--13136
		x"ff",	--13137
		x"ff",	--13138
		x"ff",	--13139
		x"ff",	--13140
		x"ff",	--13141
		x"ff",	--13142
		x"ff",	--13143
		x"ff",	--13144
		x"ff",	--13145
		x"ff",	--13146
		x"ff",	--13147
		x"ff",	--13148
		x"ff",	--13149
		x"ff",	--13150
		x"ff",	--13151
		x"ff",	--13152
		x"ff",	--13153
		x"ff",	--13154
		x"ff",	--13155
		x"ff",	--13156
		x"ff",	--13157
		x"ff",	--13158
		x"ff",	--13159
		x"ff",	--13160
		x"ff",	--13161
		x"ff",	--13162
		x"ff",	--13163
		x"ff",	--13164
		x"ff",	--13165
		x"ff",	--13166
		x"ff",	--13167
		x"ff",	--13168
		x"ff",	--13169
		x"ff",	--13170
		x"ff",	--13171
		x"ff",	--13172
		x"ff",	--13173
		x"ff",	--13174
		x"ff",	--13175
		x"ff",	--13176
		x"ff",	--13177
		x"ff",	--13178
		x"ff",	--13179
		x"ff",	--13180
		x"ff",	--13181
		x"ff",	--13182
		x"ff",	--13183
		x"ff",	--13184
		x"ff",	--13185
		x"ff",	--13186
		x"ff",	--13187
		x"ff",	--13188
		x"ff",	--13189
		x"ff",	--13190
		x"ff",	--13191
		x"ff",	--13192
		x"ff",	--13193
		x"ff",	--13194
		x"ff",	--13195
		x"ff",	--13196
		x"ff",	--13197
		x"ff",	--13198
		x"ff",	--13199
		x"ff",	--13200
		x"ff",	--13201
		x"ff",	--13202
		x"ff",	--13203
		x"ff",	--13204
		x"ff",	--13205
		x"ff",	--13206
		x"ff",	--13207
		x"ff",	--13208
		x"ff",	--13209
		x"ff",	--13210
		x"ff",	--13211
		x"ff",	--13212
		x"ff",	--13213
		x"ff",	--13214
		x"ff",	--13215
		x"ff",	--13216
		x"ff",	--13217
		x"ff",	--13218
		x"ff",	--13219
		x"ff",	--13220
		x"ff",	--13221
		x"ff",	--13222
		x"ff",	--13223
		x"ff",	--13224
		x"ff",	--13225
		x"ff",	--13226
		x"ff",	--13227
		x"ff",	--13228
		x"ff",	--13229
		x"ff",	--13230
		x"ff",	--13231
		x"ff",	--13232
		x"ff",	--13233
		x"ff",	--13234
		x"ff",	--13235
		x"ff",	--13236
		x"ff",	--13237
		x"ff",	--13238
		x"ff",	--13239
		x"ff",	--13240
		x"ff",	--13241
		x"ff",	--13242
		x"ff",	--13243
		x"ff",	--13244
		x"ff",	--13245
		x"ff",	--13246
		x"ff",	--13247
		x"ff",	--13248
		x"ff",	--13249
		x"ff",	--13250
		x"ff",	--13251
		x"ff",	--13252
		x"ff",	--13253
		x"ff",	--13254
		x"ff",	--13255
		x"ff",	--13256
		x"ff",	--13257
		x"ff",	--13258
		x"ff",	--13259
		x"ff",	--13260
		x"ff",	--13261
		x"ff",	--13262
		x"ff",	--13263
		x"ff",	--13264
		x"ff",	--13265
		x"ff",	--13266
		x"ff",	--13267
		x"ff",	--13268
		x"ff",	--13269
		x"ff",	--13270
		x"ff",	--13271
		x"ff",	--13272
		x"ff",	--13273
		x"ff",	--13274
		x"ff",	--13275
		x"ff",	--13276
		x"ff",	--13277
		x"ff",	--13278
		x"ff",	--13279
		x"ff",	--13280
		x"ff",	--13281
		x"ff",	--13282
		x"ff",	--13283
		x"ff",	--13284
		x"ff",	--13285
		x"ff",	--13286
		x"ff",	--13287
		x"ff",	--13288
		x"ff",	--13289
		x"ff",	--13290
		x"ff",	--13291
		x"ff",	--13292
		x"ff",	--13293
		x"ff",	--13294
		x"ff",	--13295
		x"ff",	--13296
		x"ff",	--13297
		x"ff",	--13298
		x"ff",	--13299
		x"ff",	--13300
		x"ff",	--13301
		x"ff",	--13302
		x"ff",	--13303
		x"ff",	--13304
		x"ff",	--13305
		x"ff",	--13306
		x"ff",	--13307
		x"ff",	--13308
		x"ff",	--13309
		x"ff",	--13310
		x"ff",	--13311
		x"ff",	--13312
		x"ff",	--13313
		x"ff",	--13314
		x"ff",	--13315
		x"ff",	--13316
		x"ff",	--13317
		x"ff",	--13318
		x"ff",	--13319
		x"ff",	--13320
		x"ff",	--13321
		x"ff",	--13322
		x"ff",	--13323
		x"ff",	--13324
		x"ff",	--13325
		x"ff",	--13326
		x"ff",	--13327
		x"ff",	--13328
		x"ff",	--13329
		x"ff",	--13330
		x"ff",	--13331
		x"ff",	--13332
		x"ff",	--13333
		x"ff",	--13334
		x"ff",	--13335
		x"ff",	--13336
		x"ff",	--13337
		x"ff",	--13338
		x"ff",	--13339
		x"ff",	--13340
		x"ff",	--13341
		x"ff",	--13342
		x"ff",	--13343
		x"ff",	--13344
		x"ff",	--13345
		x"ff",	--13346
		x"ff",	--13347
		x"ff",	--13348
		x"ff",	--13349
		x"ff",	--13350
		x"ff",	--13351
		x"ff",	--13352
		x"ff",	--13353
		x"ff",	--13354
		x"ff",	--13355
		x"ff",	--13356
		x"ff",	--13357
		x"ff",	--13358
		x"ff",	--13359
		x"ff",	--13360
		x"ff",	--13361
		x"ff",	--13362
		x"ff",	--13363
		x"ff",	--13364
		x"ff",	--13365
		x"ff",	--13366
		x"ff",	--13367
		x"ff",	--13368
		x"ff",	--13369
		x"ff",	--13370
		x"ff",	--13371
		x"ff",	--13372
		x"ff",	--13373
		x"ff",	--13374
		x"ff",	--13375
		x"ff",	--13376
		x"ff",	--13377
		x"ff",	--13378
		x"ff",	--13379
		x"ff",	--13380
		x"ff",	--13381
		x"ff",	--13382
		x"ff",	--13383
		x"ff",	--13384
		x"ff",	--13385
		x"ff",	--13386
		x"ff",	--13387
		x"ff",	--13388
		x"ff",	--13389
		x"ff",	--13390
		x"ff",	--13391
		x"ff",	--13392
		x"ff",	--13393
		x"ff",	--13394
		x"ff",	--13395
		x"ff",	--13396
		x"ff",	--13397
		x"ff",	--13398
		x"ff",	--13399
		x"ff",	--13400
		x"ff",	--13401
		x"ff",	--13402
		x"ff",	--13403
		x"ff",	--13404
		x"ff",	--13405
		x"ff",	--13406
		x"ff",	--13407
		x"ff",	--13408
		x"ff",	--13409
		x"ff",	--13410
		x"ff",	--13411
		x"ff",	--13412
		x"ff",	--13413
		x"ff",	--13414
		x"ff",	--13415
		x"ff",	--13416
		x"ff",	--13417
		x"ff",	--13418
		x"ff",	--13419
		x"ff",	--13420
		x"ff",	--13421
		x"ff",	--13422
		x"ff",	--13423
		x"ff",	--13424
		x"ff",	--13425
		x"ff",	--13426
		x"ff",	--13427
		x"ff",	--13428
		x"ff",	--13429
		x"ff",	--13430
		x"ff",	--13431
		x"ff",	--13432
		x"ff",	--13433
		x"ff",	--13434
		x"ff",	--13435
		x"ff",	--13436
		x"ff",	--13437
		x"ff",	--13438
		x"ff",	--13439
		x"ff",	--13440
		x"ff",	--13441
		x"ff",	--13442
		x"ff",	--13443
		x"ff",	--13444
		x"ff",	--13445
		x"ff",	--13446
		x"ff",	--13447
		x"ff",	--13448
		x"ff",	--13449
		x"ff",	--13450
		x"ff",	--13451
		x"ff",	--13452
		x"ff",	--13453
		x"ff",	--13454
		x"ff",	--13455
		x"ff",	--13456
		x"ff",	--13457
		x"ff",	--13458
		x"ff",	--13459
		x"ff",	--13460
		x"ff",	--13461
		x"ff",	--13462
		x"ff",	--13463
		x"ff",	--13464
		x"ff",	--13465
		x"ff",	--13466
		x"ff",	--13467
		x"ff",	--13468
		x"ff",	--13469
		x"ff",	--13470
		x"ff",	--13471
		x"ff",	--13472
		x"ff",	--13473
		x"ff",	--13474
		x"ff",	--13475
		x"ff",	--13476
		x"ff",	--13477
		x"ff",	--13478
		x"ff",	--13479
		x"ff",	--13480
		x"ff",	--13481
		x"ff",	--13482
		x"ff",	--13483
		x"ff",	--13484
		x"ff",	--13485
		x"ff",	--13486
		x"ff",	--13487
		x"ff",	--13488
		x"ff",	--13489
		x"ff",	--13490
		x"ff",	--13491
		x"ff",	--13492
		x"ff",	--13493
		x"ff",	--13494
		x"ff",	--13495
		x"ff",	--13496
		x"ff",	--13497
		x"ff",	--13498
		x"ff",	--13499
		x"ff",	--13500
		x"ff",	--13501
		x"ff",	--13502
		x"ff",	--13503
		x"ff",	--13504
		x"ff",	--13505
		x"ff",	--13506
		x"ff",	--13507
		x"ff",	--13508
		x"ff",	--13509
		x"ff",	--13510
		x"ff",	--13511
		x"ff",	--13512
		x"ff",	--13513
		x"ff",	--13514
		x"ff",	--13515
		x"ff",	--13516
		x"ff",	--13517
		x"ff",	--13518
		x"ff",	--13519
		x"ff",	--13520
		x"ff",	--13521
		x"ff",	--13522
		x"ff",	--13523
		x"ff",	--13524
		x"ff",	--13525
		x"ff",	--13526
		x"ff",	--13527
		x"ff",	--13528
		x"ff",	--13529
		x"ff",	--13530
		x"ff",	--13531
		x"ff",	--13532
		x"ff",	--13533
		x"ff",	--13534
		x"ff",	--13535
		x"ff",	--13536
		x"ff",	--13537
		x"ff",	--13538
		x"ff",	--13539
		x"ff",	--13540
		x"ff",	--13541
		x"ff",	--13542
		x"ff",	--13543
		x"ff",	--13544
		x"ff",	--13545
		x"ff",	--13546
		x"ff",	--13547
		x"ff",	--13548
		x"ff",	--13549
		x"ff",	--13550
		x"ff",	--13551
		x"ff",	--13552
		x"ff",	--13553
		x"ff",	--13554
		x"ff",	--13555
		x"ff",	--13556
		x"ff",	--13557
		x"ff",	--13558
		x"ff",	--13559
		x"ff",	--13560
		x"ff",	--13561
		x"ff",	--13562
		x"ff",	--13563
		x"ff",	--13564
		x"ff",	--13565
		x"ff",	--13566
		x"ff",	--13567
		x"ff",	--13568
		x"ff",	--13569
		x"ff",	--13570
		x"ff",	--13571
		x"ff",	--13572
		x"ff",	--13573
		x"ff",	--13574
		x"ff",	--13575
		x"ff",	--13576
		x"ff",	--13577
		x"ff",	--13578
		x"ff",	--13579
		x"ff",	--13580
		x"ff",	--13581
		x"ff",	--13582
		x"ff",	--13583
		x"ff",	--13584
		x"ff",	--13585
		x"ff",	--13586
		x"ff",	--13587
		x"ff",	--13588
		x"ff",	--13589
		x"ff",	--13590
		x"ff",	--13591
		x"ff",	--13592
		x"ff",	--13593
		x"ff",	--13594
		x"ff",	--13595
		x"ff",	--13596
		x"ff",	--13597
		x"ff",	--13598
		x"ff",	--13599
		x"ff",	--13600
		x"ff",	--13601
		x"ff",	--13602
		x"ff",	--13603
		x"ff",	--13604
		x"ff",	--13605
		x"ff",	--13606
		x"ff",	--13607
		x"ff",	--13608
		x"ff",	--13609
		x"ff",	--13610
		x"ff",	--13611
		x"ff",	--13612
		x"ff",	--13613
		x"ff",	--13614
		x"ff",	--13615
		x"ff",	--13616
		x"ff",	--13617
		x"ff",	--13618
		x"ff",	--13619
		x"ff",	--13620
		x"ff",	--13621
		x"ff",	--13622
		x"ff",	--13623
		x"ff",	--13624
		x"ff",	--13625
		x"ff",	--13626
		x"ff",	--13627
		x"ff",	--13628
		x"ff",	--13629
		x"ff",	--13630
		x"ff",	--13631
		x"ff",	--13632
		x"ff",	--13633
		x"ff",	--13634
		x"ff",	--13635
		x"ff",	--13636
		x"ff",	--13637
		x"ff",	--13638
		x"ff",	--13639
		x"ff",	--13640
		x"ff",	--13641
		x"ff",	--13642
		x"ff",	--13643
		x"ff",	--13644
		x"ff",	--13645
		x"ff",	--13646
		x"ff",	--13647
		x"ff",	--13648
		x"ff",	--13649
		x"ff",	--13650
		x"ff",	--13651
		x"ff",	--13652
		x"ff",	--13653
		x"ff",	--13654
		x"ff",	--13655
		x"ff",	--13656
		x"ff",	--13657
		x"ff",	--13658
		x"ff",	--13659
		x"ff",	--13660
		x"ff",	--13661
		x"ff",	--13662
		x"ff",	--13663
		x"ff",	--13664
		x"ff",	--13665
		x"ff",	--13666
		x"ff",	--13667
		x"ff",	--13668
		x"ff",	--13669
		x"ff",	--13670
		x"ff",	--13671
		x"ff",	--13672
		x"ff",	--13673
		x"ff",	--13674
		x"ff",	--13675
		x"ff",	--13676
		x"ff",	--13677
		x"ff",	--13678
		x"ff",	--13679
		x"ff",	--13680
		x"ff",	--13681
		x"ff",	--13682
		x"ff",	--13683
		x"ff",	--13684
		x"ff",	--13685
		x"ff",	--13686
		x"ff",	--13687
		x"ff",	--13688
		x"ff",	--13689
		x"ff",	--13690
		x"ff",	--13691
		x"ff",	--13692
		x"ff",	--13693
		x"ff",	--13694
		x"ff",	--13695
		x"ff",	--13696
		x"ff",	--13697
		x"ff",	--13698
		x"ff",	--13699
		x"ff",	--13700
		x"ff",	--13701
		x"ff",	--13702
		x"ff",	--13703
		x"ff",	--13704
		x"ff",	--13705
		x"ff",	--13706
		x"ff",	--13707
		x"ff",	--13708
		x"ff",	--13709
		x"ff",	--13710
		x"ff",	--13711
		x"ff",	--13712
		x"ff",	--13713
		x"ff",	--13714
		x"ff",	--13715
		x"ff",	--13716
		x"ff",	--13717
		x"ff",	--13718
		x"ff",	--13719
		x"ff",	--13720
		x"ff",	--13721
		x"ff",	--13722
		x"ff",	--13723
		x"ff",	--13724
		x"ff",	--13725
		x"ff",	--13726
		x"ff",	--13727
		x"ff",	--13728
		x"ff",	--13729
		x"ff",	--13730
		x"ff",	--13731
		x"ff",	--13732
		x"ff",	--13733
		x"ff",	--13734
		x"ff",	--13735
		x"ff",	--13736
		x"ff",	--13737
		x"ff",	--13738
		x"ff",	--13739
		x"ff",	--13740
		x"ff",	--13741
		x"ff",	--13742
		x"ff",	--13743
		x"ff",	--13744
		x"ff",	--13745
		x"ff",	--13746
		x"ff",	--13747
		x"ff",	--13748
		x"ff",	--13749
		x"ff",	--13750
		x"ff",	--13751
		x"ff",	--13752
		x"ff",	--13753
		x"ff",	--13754
		x"ff",	--13755
		x"ff",	--13756
		x"ff",	--13757
		x"ff",	--13758
		x"ff",	--13759
		x"ff",	--13760
		x"ff",	--13761
		x"ff",	--13762
		x"ff",	--13763
		x"ff",	--13764
		x"ff",	--13765
		x"ff",	--13766
		x"ff",	--13767
		x"ff",	--13768
		x"ff",	--13769
		x"ff",	--13770
		x"ff",	--13771
		x"ff",	--13772
		x"ff",	--13773
		x"ff",	--13774
		x"ff",	--13775
		x"ff",	--13776
		x"ff",	--13777
		x"ff",	--13778
		x"ff",	--13779
		x"ff",	--13780
		x"ff",	--13781
		x"ff",	--13782
		x"ff",	--13783
		x"ff",	--13784
		x"ff",	--13785
		x"ff",	--13786
		x"ff",	--13787
		x"ff",	--13788
		x"ff",	--13789
		x"ff",	--13790
		x"ff",	--13791
		x"ff",	--13792
		x"ff",	--13793
		x"ff",	--13794
		x"ff",	--13795
		x"ff",	--13796
		x"ff",	--13797
		x"ff",	--13798
		x"ff",	--13799
		x"ff",	--13800
		x"ff",	--13801
		x"ff",	--13802
		x"ff",	--13803
		x"ff",	--13804
		x"ff",	--13805
		x"ff",	--13806
		x"ff",	--13807
		x"ff",	--13808
		x"ff",	--13809
		x"ff",	--13810
		x"ff",	--13811
		x"ff",	--13812
		x"ff",	--13813
		x"ff",	--13814
		x"ff",	--13815
		x"ff",	--13816
		x"ff",	--13817
		x"ff",	--13818
		x"ff",	--13819
		x"ff",	--13820
		x"ff",	--13821
		x"ff",	--13822
		x"ff",	--13823
		x"ff",	--13824
		x"ff",	--13825
		x"ff",	--13826
		x"ff",	--13827
		x"ff",	--13828
		x"ff",	--13829
		x"ff",	--13830
		x"ff",	--13831
		x"ff",	--13832
		x"ff",	--13833
		x"ff",	--13834
		x"ff",	--13835
		x"ff",	--13836
		x"ff",	--13837
		x"ff",	--13838
		x"ff",	--13839
		x"ff",	--13840
		x"ff",	--13841
		x"ff",	--13842
		x"ff",	--13843
		x"ff",	--13844
		x"ff",	--13845
		x"ff",	--13846
		x"ff",	--13847
		x"ff",	--13848
		x"ff",	--13849
		x"ff",	--13850
		x"ff",	--13851
		x"ff",	--13852
		x"ff",	--13853
		x"ff",	--13854
		x"ff",	--13855
		x"ff",	--13856
		x"ff",	--13857
		x"ff",	--13858
		x"ff",	--13859
		x"ff",	--13860
		x"ff",	--13861
		x"ff",	--13862
		x"ff",	--13863
		x"ff",	--13864
		x"ff",	--13865
		x"ff",	--13866
		x"ff",	--13867
		x"ff",	--13868
		x"ff",	--13869
		x"ff",	--13870
		x"ff",	--13871
		x"ff",	--13872
		x"ff",	--13873
		x"ff",	--13874
		x"ff",	--13875
		x"ff",	--13876
		x"ff",	--13877
		x"ff",	--13878
		x"ff",	--13879
		x"ff",	--13880
		x"ff",	--13881
		x"ff",	--13882
		x"ff",	--13883
		x"ff",	--13884
		x"ff",	--13885
		x"ff",	--13886
		x"ff",	--13887
		x"ff",	--13888
		x"ff",	--13889
		x"ff",	--13890
		x"ff",	--13891
		x"ff",	--13892
		x"ff",	--13893
		x"ff",	--13894
		x"ff",	--13895
		x"ff",	--13896
		x"ff",	--13897
		x"ff",	--13898
		x"ff",	--13899
		x"ff",	--13900
		x"ff",	--13901
		x"ff",	--13902
		x"ff",	--13903
		x"ff",	--13904
		x"ff",	--13905
		x"ff",	--13906
		x"ff",	--13907
		x"ff",	--13908
		x"ff",	--13909
		x"ff",	--13910
		x"ff",	--13911
		x"ff",	--13912
		x"ff",	--13913
		x"ff",	--13914
		x"ff",	--13915
		x"ff",	--13916
		x"ff",	--13917
		x"ff",	--13918
		x"ff",	--13919
		x"ff",	--13920
		x"ff",	--13921
		x"ff",	--13922
		x"ff",	--13923
		x"ff",	--13924
		x"ff",	--13925
		x"ff",	--13926
		x"ff",	--13927
		x"ff",	--13928
		x"ff",	--13929
		x"ff",	--13930
		x"ff",	--13931
		x"ff",	--13932
		x"ff",	--13933
		x"ff",	--13934
		x"ff",	--13935
		x"ff",	--13936
		x"ff",	--13937
		x"ff",	--13938
		x"ff",	--13939
		x"ff",	--13940
		x"ff",	--13941
		x"ff",	--13942
		x"ff",	--13943
		x"ff",	--13944
		x"ff",	--13945
		x"ff",	--13946
		x"ff",	--13947
		x"ff",	--13948
		x"ff",	--13949
		x"ff",	--13950
		x"ff",	--13951
		x"ff",	--13952
		x"ff",	--13953
		x"ff",	--13954
		x"ff",	--13955
		x"ff",	--13956
		x"ff",	--13957
		x"ff",	--13958
		x"ff",	--13959
		x"ff",	--13960
		x"ff",	--13961
		x"ff",	--13962
		x"ff",	--13963
		x"ff",	--13964
		x"ff",	--13965
		x"ff",	--13966
		x"ff",	--13967
		x"ff",	--13968
		x"ff",	--13969
		x"ff",	--13970
		x"ff",	--13971
		x"ff",	--13972
		x"ff",	--13973
		x"ff",	--13974
		x"ff",	--13975
		x"ff",	--13976
		x"ff",	--13977
		x"ff",	--13978
		x"ff",	--13979
		x"ff",	--13980
		x"ff",	--13981
		x"ff",	--13982
		x"ff",	--13983
		x"ff",	--13984
		x"ff",	--13985
		x"ff",	--13986
		x"ff",	--13987
		x"ff",	--13988
		x"ff",	--13989
		x"ff",	--13990
		x"ff",	--13991
		x"ff",	--13992
		x"ff",	--13993
		x"ff",	--13994
		x"ff",	--13995
		x"ff",	--13996
		x"ff",	--13997
		x"ff",	--13998
		x"ff",	--13999
		x"ff",	--14000
		x"ff",	--14001
		x"ff",	--14002
		x"ff",	--14003
		x"ff",	--14004
		x"ff",	--14005
		x"ff",	--14006
		x"ff",	--14007
		x"ff",	--14008
		x"ff",	--14009
		x"ff",	--14010
		x"ff",	--14011
		x"ff",	--14012
		x"ff",	--14013
		x"ff",	--14014
		x"ff",	--14015
		x"ff",	--14016
		x"ff",	--14017
		x"ff",	--14018
		x"ff",	--14019
		x"ff",	--14020
		x"ff",	--14021
		x"ff",	--14022
		x"ff",	--14023
		x"ff",	--14024
		x"ff",	--14025
		x"ff",	--14026
		x"ff",	--14027
		x"ff",	--14028
		x"ff",	--14029
		x"ff",	--14030
		x"ff",	--14031
		x"ff",	--14032
		x"ff",	--14033
		x"ff",	--14034
		x"ff",	--14035
		x"ff",	--14036
		x"ff",	--14037
		x"ff",	--14038
		x"ff",	--14039
		x"ff",	--14040
		x"ff",	--14041
		x"ff",	--14042
		x"ff",	--14043
		x"ff",	--14044
		x"ff",	--14045
		x"ff",	--14046
		x"ff",	--14047
		x"ff",	--14048
		x"ff",	--14049
		x"ff",	--14050
		x"ff",	--14051
		x"ff",	--14052
		x"ff",	--14053
		x"ff",	--14054
		x"ff",	--14055
		x"ff",	--14056
		x"ff",	--14057
		x"ff",	--14058
		x"ff",	--14059
		x"ff",	--14060
		x"ff",	--14061
		x"ff",	--14062
		x"ff",	--14063
		x"ff",	--14064
		x"ff",	--14065
		x"ff",	--14066
		x"ff",	--14067
		x"ff",	--14068
		x"ff",	--14069
		x"ff",	--14070
		x"ff",	--14071
		x"ff",	--14072
		x"ff",	--14073
		x"ff",	--14074
		x"ff",	--14075
		x"ff",	--14076
		x"ff",	--14077
		x"ff",	--14078
		x"ff",	--14079
		x"ff",	--14080
		x"ff",	--14081
		x"ff",	--14082
		x"ff",	--14083
		x"ff",	--14084
		x"ff",	--14085
		x"ff",	--14086
		x"ff",	--14087
		x"ff",	--14088
		x"ff",	--14089
		x"ff",	--14090
		x"ff",	--14091
		x"ff",	--14092
		x"ff",	--14093
		x"ff",	--14094
		x"ff",	--14095
		x"ff",	--14096
		x"ff",	--14097
		x"ff",	--14098
		x"ff",	--14099
		x"ff",	--14100
		x"ff",	--14101
		x"ff",	--14102
		x"ff",	--14103
		x"ff",	--14104
		x"ff",	--14105
		x"ff",	--14106
		x"ff",	--14107
		x"ff",	--14108
		x"ff",	--14109
		x"ff",	--14110
		x"ff",	--14111
		x"ff",	--14112
		x"ff",	--14113
		x"ff",	--14114
		x"ff",	--14115
		x"ff",	--14116
		x"ff",	--14117
		x"ff",	--14118
		x"ff",	--14119
		x"ff",	--14120
		x"ff",	--14121
		x"ff",	--14122
		x"ff",	--14123
		x"ff",	--14124
		x"ff",	--14125
		x"ff",	--14126
		x"ff",	--14127
		x"ff",	--14128
		x"ff",	--14129
		x"ff",	--14130
		x"ff",	--14131
		x"ff",	--14132
		x"ff",	--14133
		x"ff",	--14134
		x"ff",	--14135
		x"ff",	--14136
		x"ff",	--14137
		x"ff",	--14138
		x"ff",	--14139
		x"ff",	--14140
		x"ff",	--14141
		x"ff",	--14142
		x"ff",	--14143
		x"ff",	--14144
		x"ff",	--14145
		x"ff",	--14146
		x"ff",	--14147
		x"ff",	--14148
		x"ff",	--14149
		x"ff",	--14150
		x"ff",	--14151
		x"ff",	--14152
		x"ff",	--14153
		x"ff",	--14154
		x"ff",	--14155
		x"ff",	--14156
		x"ff",	--14157
		x"ff",	--14158
		x"ff",	--14159
		x"ff",	--14160
		x"ff",	--14161
		x"ff",	--14162
		x"ff",	--14163
		x"ff",	--14164
		x"ff",	--14165
		x"ff",	--14166
		x"ff",	--14167
		x"ff",	--14168
		x"ff",	--14169
		x"ff",	--14170
		x"ff",	--14171
		x"ff",	--14172
		x"ff",	--14173
		x"ff",	--14174
		x"ff",	--14175
		x"ff",	--14176
		x"ff",	--14177
		x"ff",	--14178
		x"ff",	--14179
		x"ff",	--14180
		x"ff",	--14181
		x"ff",	--14182
		x"ff",	--14183
		x"ff",	--14184
		x"ff",	--14185
		x"ff",	--14186
		x"ff",	--14187
		x"ff",	--14188
		x"ff",	--14189
		x"ff",	--14190
		x"ff",	--14191
		x"ff",	--14192
		x"ff",	--14193
		x"ff",	--14194
		x"ff",	--14195
		x"ff",	--14196
		x"ff",	--14197
		x"ff",	--14198
		x"ff",	--14199
		x"ff",	--14200
		x"ff",	--14201
		x"ff",	--14202
		x"ff",	--14203
		x"ff",	--14204
		x"ff",	--14205
		x"ff",	--14206
		x"ff",	--14207
		x"ff",	--14208
		x"ff",	--14209
		x"ff",	--14210
		x"ff",	--14211
		x"ff",	--14212
		x"ff",	--14213
		x"ff",	--14214
		x"ff",	--14215
		x"ff",	--14216
		x"ff",	--14217
		x"ff",	--14218
		x"ff",	--14219
		x"ff",	--14220
		x"ff",	--14221
		x"ff",	--14222
		x"ff",	--14223
		x"ff",	--14224
		x"ff",	--14225
		x"ff",	--14226
		x"ff",	--14227
		x"ff",	--14228
		x"ff",	--14229
		x"ff",	--14230
		x"ff",	--14231
		x"ff",	--14232
		x"ff",	--14233
		x"ff",	--14234
		x"ff",	--14235
		x"ff",	--14236
		x"ff",	--14237
		x"ff",	--14238
		x"ff",	--14239
		x"ff",	--14240
		x"ff",	--14241
		x"ff",	--14242
		x"ff",	--14243
		x"ff",	--14244
		x"ff",	--14245
		x"ff",	--14246
		x"ff",	--14247
		x"ff",	--14248
		x"ff",	--14249
		x"ff",	--14250
		x"ff",	--14251
		x"ff",	--14252
		x"ff",	--14253
		x"ff",	--14254
		x"ff",	--14255
		x"ff",	--14256
		x"ff",	--14257
		x"ff",	--14258
		x"ff",	--14259
		x"ff",	--14260
		x"ff",	--14261
		x"ff",	--14262
		x"ff",	--14263
		x"ff",	--14264
		x"ff",	--14265
		x"ff",	--14266
		x"ff",	--14267
		x"ff",	--14268
		x"ff",	--14269
		x"ff",	--14270
		x"ff",	--14271
		x"ff",	--14272
		x"ff",	--14273
		x"ff",	--14274
		x"ff",	--14275
		x"ff",	--14276
		x"ff",	--14277
		x"ff",	--14278
		x"ff",	--14279
		x"ff",	--14280
		x"ff",	--14281
		x"ff",	--14282
		x"ff",	--14283
		x"ff",	--14284
		x"ff",	--14285
		x"ff",	--14286
		x"ff",	--14287
		x"ff",	--14288
		x"ff",	--14289
		x"ff",	--14290
		x"ff",	--14291
		x"ff",	--14292
		x"ff",	--14293
		x"ff",	--14294
		x"ff",	--14295
		x"ff",	--14296
		x"ff",	--14297
		x"ff",	--14298
		x"ff",	--14299
		x"ff",	--14300
		x"ff",	--14301
		x"ff",	--14302
		x"ff",	--14303
		x"ff",	--14304
		x"ff",	--14305
		x"ff",	--14306
		x"ff",	--14307
		x"ff",	--14308
		x"ff",	--14309
		x"ff",	--14310
		x"ff",	--14311
		x"ff",	--14312
		x"ff",	--14313
		x"ff",	--14314
		x"ff",	--14315
		x"ff",	--14316
		x"ff",	--14317
		x"ff",	--14318
		x"ff",	--14319
		x"ff",	--14320
		x"ff",	--14321
		x"ff",	--14322
		x"ff",	--14323
		x"ff",	--14324
		x"ff",	--14325
		x"ff",	--14326
		x"ff",	--14327
		x"ff",	--14328
		x"ff",	--14329
		x"ff",	--14330
		x"ff",	--14331
		x"ff",	--14332
		x"ff",	--14333
		x"ff",	--14334
		x"ff",	--14335
		x"ff",	--14336
		x"ff",	--14337
		x"ff",	--14338
		x"ff",	--14339
		x"ff",	--14340
		x"ff",	--14341
		x"ff",	--14342
		x"ff",	--14343
		x"ff",	--14344
		x"ff",	--14345
		x"ff",	--14346
		x"ff",	--14347
		x"ff",	--14348
		x"ff",	--14349
		x"ff",	--14350
		x"ff",	--14351
		x"ff",	--14352
		x"ff",	--14353
		x"ff",	--14354
		x"ff",	--14355
		x"ff",	--14356
		x"ff",	--14357
		x"ff",	--14358
		x"ff",	--14359
		x"ff",	--14360
		x"ff",	--14361
		x"ff",	--14362
		x"ff",	--14363
		x"ff",	--14364
		x"ff",	--14365
		x"ff",	--14366
		x"ff",	--14367
		x"ff",	--14368
		x"ff",	--14369
		x"ff",	--14370
		x"ff",	--14371
		x"ff",	--14372
		x"ff",	--14373
		x"ff",	--14374
		x"ff",	--14375
		x"ff",	--14376
		x"ff",	--14377
		x"ff",	--14378
		x"ff",	--14379
		x"ff",	--14380
		x"ff",	--14381
		x"ff",	--14382
		x"ff",	--14383
		x"ff",	--14384
		x"ff",	--14385
		x"ff",	--14386
		x"ff",	--14387
		x"ff",	--14388
		x"ff",	--14389
		x"ff",	--14390
		x"ff",	--14391
		x"ff",	--14392
		x"ff",	--14393
		x"ff",	--14394
		x"ff",	--14395
		x"ff",	--14396
		x"ff",	--14397
		x"ff",	--14398
		x"ff",	--14399
		x"ff",	--14400
		x"ff",	--14401
		x"ff",	--14402
		x"ff",	--14403
		x"ff",	--14404
		x"ff",	--14405
		x"ff",	--14406
		x"ff",	--14407
		x"ff",	--14408
		x"ff",	--14409
		x"ff",	--14410
		x"ff",	--14411
		x"ff",	--14412
		x"ff",	--14413
		x"ff",	--14414
		x"ff",	--14415
		x"ff",	--14416
		x"ff",	--14417
		x"ff",	--14418
		x"ff",	--14419
		x"ff",	--14420
		x"ff",	--14421
		x"ff",	--14422
		x"ff",	--14423
		x"ff",	--14424
		x"ff",	--14425
		x"ff",	--14426
		x"ff",	--14427
		x"ff",	--14428
		x"ff",	--14429
		x"ff",	--14430
		x"ff",	--14431
		x"ff",	--14432
		x"ff",	--14433
		x"ff",	--14434
		x"ff",	--14435
		x"ff",	--14436
		x"ff",	--14437
		x"ff",	--14438
		x"ff",	--14439
		x"ff",	--14440
		x"ff",	--14441
		x"ff",	--14442
		x"ff",	--14443
		x"ff",	--14444
		x"ff",	--14445
		x"ff",	--14446
		x"ff",	--14447
		x"ff",	--14448
		x"ff",	--14449
		x"ff",	--14450
		x"ff",	--14451
		x"ff",	--14452
		x"ff",	--14453
		x"ff",	--14454
		x"ff",	--14455
		x"ff",	--14456
		x"ff",	--14457
		x"ff",	--14458
		x"ff",	--14459
		x"ff",	--14460
		x"ff",	--14461
		x"ff",	--14462
		x"ff",	--14463
		x"ff",	--14464
		x"ff",	--14465
		x"ff",	--14466
		x"ff",	--14467
		x"ff",	--14468
		x"ff",	--14469
		x"ff",	--14470
		x"ff",	--14471
		x"ff",	--14472
		x"ff",	--14473
		x"ff",	--14474
		x"ff",	--14475
		x"ff",	--14476
		x"ff",	--14477
		x"ff",	--14478
		x"ff",	--14479
		x"ff",	--14480
		x"ff",	--14481
		x"ff",	--14482
		x"ff",	--14483
		x"ff",	--14484
		x"ff",	--14485
		x"ff",	--14486
		x"ff",	--14487
		x"ff",	--14488
		x"ff",	--14489
		x"ff",	--14490
		x"ff",	--14491
		x"ff",	--14492
		x"ff",	--14493
		x"ff",	--14494
		x"ff",	--14495
		x"ff",	--14496
		x"ff",	--14497
		x"ff",	--14498
		x"ff",	--14499
		x"ff",	--14500
		x"ff",	--14501
		x"ff",	--14502
		x"ff",	--14503
		x"ff",	--14504
		x"ff",	--14505
		x"ff",	--14506
		x"ff",	--14507
		x"ff",	--14508
		x"ff",	--14509
		x"ff",	--14510
		x"ff",	--14511
		x"ff",	--14512
		x"ff",	--14513
		x"ff",	--14514
		x"ff",	--14515
		x"ff",	--14516
		x"ff",	--14517
		x"ff",	--14518
		x"ff",	--14519
		x"ff",	--14520
		x"ff",	--14521
		x"ff",	--14522
		x"ff",	--14523
		x"ff",	--14524
		x"ff",	--14525
		x"ff",	--14526
		x"ff",	--14527
		x"ff",	--14528
		x"ff",	--14529
		x"ff",	--14530
		x"ff",	--14531
		x"ff",	--14532
		x"ff",	--14533
		x"ff",	--14534
		x"ff",	--14535
		x"ff",	--14536
		x"ff",	--14537
		x"ff",	--14538
		x"ff",	--14539
		x"ff",	--14540
		x"ff",	--14541
		x"ff",	--14542
		x"ff",	--14543
		x"ff",	--14544
		x"ff",	--14545
		x"ff",	--14546
		x"ff",	--14547
		x"ff",	--14548
		x"ff",	--14549
		x"ff",	--14550
		x"ff",	--14551
		x"ff",	--14552
		x"ff",	--14553
		x"ff",	--14554
		x"ff",	--14555
		x"ff",	--14556
		x"ff",	--14557
		x"ff",	--14558
		x"ff",	--14559
		x"ff",	--14560
		x"ff",	--14561
		x"ff",	--14562
		x"ff",	--14563
		x"ff",	--14564
		x"ff",	--14565
		x"ff",	--14566
		x"ff",	--14567
		x"ff",	--14568
		x"ff",	--14569
		x"ff",	--14570
		x"ff",	--14571
		x"ff",	--14572
		x"ff",	--14573
		x"ff",	--14574
		x"ff",	--14575
		x"ff",	--14576
		x"ff",	--14577
		x"ff",	--14578
		x"ff",	--14579
		x"ff",	--14580
		x"ff",	--14581
		x"ff",	--14582
		x"ff",	--14583
		x"ff",	--14584
		x"ff",	--14585
		x"ff",	--14586
		x"ff",	--14587
		x"ff",	--14588
		x"ff",	--14589
		x"ff",	--14590
		x"ff",	--14591
		x"ff",	--14592
		x"ff",	--14593
		x"ff",	--14594
		x"ff",	--14595
		x"ff",	--14596
		x"ff",	--14597
		x"ff",	--14598
		x"ff",	--14599
		x"ff",	--14600
		x"ff",	--14601
		x"ff",	--14602
		x"ff",	--14603
		x"ff",	--14604
		x"ff",	--14605
		x"ff",	--14606
		x"ff",	--14607
		x"ff",	--14608
		x"ff",	--14609
		x"ff",	--14610
		x"ff",	--14611
		x"ff",	--14612
		x"ff",	--14613
		x"ff",	--14614
		x"ff",	--14615
		x"ff",	--14616
		x"ff",	--14617
		x"ff",	--14618
		x"ff",	--14619
		x"ff",	--14620
		x"ff",	--14621
		x"ff",	--14622
		x"ff",	--14623
		x"ff",	--14624
		x"ff",	--14625
		x"ff",	--14626
		x"ff",	--14627
		x"ff",	--14628
		x"ff",	--14629
		x"ff",	--14630
		x"ff",	--14631
		x"ff",	--14632
		x"ff",	--14633
		x"ff",	--14634
		x"ff",	--14635
		x"ff",	--14636
		x"ff",	--14637
		x"ff",	--14638
		x"ff",	--14639
		x"ff",	--14640
		x"ff",	--14641
		x"ff",	--14642
		x"ff",	--14643
		x"ff",	--14644
		x"ff",	--14645
		x"ff",	--14646
		x"ff",	--14647
		x"ff",	--14648
		x"ff",	--14649
		x"ff",	--14650
		x"ff",	--14651
		x"ff",	--14652
		x"ff",	--14653
		x"ff",	--14654
		x"ff",	--14655
		x"ff",	--14656
		x"ff",	--14657
		x"ff",	--14658
		x"ff",	--14659
		x"ff",	--14660
		x"ff",	--14661
		x"ff",	--14662
		x"ff",	--14663
		x"ff",	--14664
		x"ff",	--14665
		x"ff",	--14666
		x"ff",	--14667
		x"ff",	--14668
		x"ff",	--14669
		x"ff",	--14670
		x"ff",	--14671
		x"ff",	--14672
		x"ff",	--14673
		x"ff",	--14674
		x"ff",	--14675
		x"ff",	--14676
		x"ff",	--14677
		x"ff",	--14678
		x"ff",	--14679
		x"ff",	--14680
		x"ff",	--14681
		x"ff",	--14682
		x"ff",	--14683
		x"ff",	--14684
		x"ff",	--14685
		x"ff",	--14686
		x"ff",	--14687
		x"ff",	--14688
		x"ff",	--14689
		x"ff",	--14690
		x"ff",	--14691
		x"ff",	--14692
		x"ff",	--14693
		x"ff",	--14694
		x"ff",	--14695
		x"ff",	--14696
		x"ff",	--14697
		x"ff",	--14698
		x"ff",	--14699
		x"ff",	--14700
		x"ff",	--14701
		x"ff",	--14702
		x"ff",	--14703
		x"ff",	--14704
		x"ff",	--14705
		x"ff",	--14706
		x"ff",	--14707
		x"ff",	--14708
		x"ff",	--14709
		x"ff",	--14710
		x"ff",	--14711
		x"ff",	--14712
		x"ff",	--14713
		x"ff",	--14714
		x"ff",	--14715
		x"ff",	--14716
		x"ff",	--14717
		x"ff",	--14718
		x"ff",	--14719
		x"ff",	--14720
		x"ff",	--14721
		x"ff",	--14722
		x"ff",	--14723
		x"ff",	--14724
		x"ff",	--14725
		x"ff",	--14726
		x"ff",	--14727
		x"ff",	--14728
		x"ff",	--14729
		x"ff",	--14730
		x"ff",	--14731
		x"ff",	--14732
		x"ff",	--14733
		x"ff",	--14734
		x"ff",	--14735
		x"ff",	--14736
		x"ff",	--14737
		x"ff",	--14738
		x"ff",	--14739
		x"ff",	--14740
		x"ff",	--14741
		x"ff",	--14742
		x"ff",	--14743
		x"ff",	--14744
		x"ff",	--14745
		x"ff",	--14746
		x"ff",	--14747
		x"ff",	--14748
		x"ff",	--14749
		x"ff",	--14750
		x"ff",	--14751
		x"ff",	--14752
		x"ff",	--14753
		x"ff",	--14754
		x"ff",	--14755
		x"ff",	--14756
		x"ff",	--14757
		x"ff",	--14758
		x"ff",	--14759
		x"ff",	--14760
		x"ff",	--14761
		x"ff",	--14762
		x"ff",	--14763
		x"ff",	--14764
		x"ff",	--14765
		x"ff",	--14766
		x"ff",	--14767
		x"ff",	--14768
		x"ff",	--14769
		x"ff",	--14770
		x"ff",	--14771
		x"ff",	--14772
		x"ff",	--14773
		x"ff",	--14774
		x"ff",	--14775
		x"ff",	--14776
		x"ff",	--14777
		x"ff",	--14778
		x"ff",	--14779
		x"ff",	--14780
		x"ff",	--14781
		x"ff",	--14782
		x"ff",	--14783
		x"ff",	--14784
		x"ff",	--14785
		x"ff",	--14786
		x"ff",	--14787
		x"ff",	--14788
		x"ff",	--14789
		x"ff",	--14790
		x"ff",	--14791
		x"ff",	--14792
		x"ff",	--14793
		x"ff",	--14794
		x"ff",	--14795
		x"ff",	--14796
		x"ff",	--14797
		x"ff",	--14798
		x"ff",	--14799
		x"ff",	--14800
		x"ff",	--14801
		x"ff",	--14802
		x"ff",	--14803
		x"ff",	--14804
		x"ff",	--14805
		x"ff",	--14806
		x"ff",	--14807
		x"ff",	--14808
		x"ff",	--14809
		x"ff",	--14810
		x"ff",	--14811
		x"ff",	--14812
		x"ff",	--14813
		x"ff",	--14814
		x"ff",	--14815
		x"ff",	--14816
		x"ff",	--14817
		x"ff",	--14818
		x"ff",	--14819
		x"ff",	--14820
		x"ff",	--14821
		x"ff",	--14822
		x"ff",	--14823
		x"ff",	--14824
		x"ff",	--14825
		x"ff",	--14826
		x"ff",	--14827
		x"ff",	--14828
		x"ff",	--14829
		x"ff",	--14830
		x"ff",	--14831
		x"ff",	--14832
		x"ff",	--14833
		x"ff",	--14834
		x"ff",	--14835
		x"ff",	--14836
		x"ff",	--14837
		x"ff",	--14838
		x"ff",	--14839
		x"ff",	--14840
		x"ff",	--14841
		x"ff",	--14842
		x"ff",	--14843
		x"ff",	--14844
		x"ff",	--14845
		x"ff",	--14846
		x"ff",	--14847
		x"ff",	--14848
		x"ff",	--14849
		x"ff",	--14850
		x"ff",	--14851
		x"ff",	--14852
		x"ff",	--14853
		x"ff",	--14854
		x"ff",	--14855
		x"ff",	--14856
		x"ff",	--14857
		x"ff",	--14858
		x"ff",	--14859
		x"ff",	--14860
		x"ff",	--14861
		x"ff",	--14862
		x"ff",	--14863
		x"ff",	--14864
		x"ff",	--14865
		x"ff",	--14866
		x"ff",	--14867
		x"ff",	--14868
		x"ff",	--14869
		x"ff",	--14870
		x"ff",	--14871
		x"ff",	--14872
		x"ff",	--14873
		x"ff",	--14874
		x"ff",	--14875
		x"ff",	--14876
		x"ff",	--14877
		x"ff",	--14878
		x"ff",	--14879
		x"ff",	--14880
		x"ff",	--14881
		x"ff",	--14882
		x"ff",	--14883
		x"ff",	--14884
		x"ff",	--14885
		x"ff",	--14886
		x"ff",	--14887
		x"ff",	--14888
		x"ff",	--14889
		x"ff",	--14890
		x"ff",	--14891
		x"ff",	--14892
		x"ff",	--14893
		x"ff",	--14894
		x"ff",	--14895
		x"ff",	--14896
		x"ff",	--14897
		x"ff",	--14898
		x"ff",	--14899
		x"ff",	--14900
		x"ff",	--14901
		x"ff",	--14902
		x"ff",	--14903
		x"ff",	--14904
		x"ff",	--14905
		x"ff",	--14906
		x"ff",	--14907
		x"ff",	--14908
		x"ff",	--14909
		x"ff",	--14910
		x"ff",	--14911
		x"ff",	--14912
		x"ff",	--14913
		x"ff",	--14914
		x"ff",	--14915
		x"ff",	--14916
		x"ff",	--14917
		x"ff",	--14918
		x"ff",	--14919
		x"ff",	--14920
		x"ff",	--14921
		x"ff",	--14922
		x"ff",	--14923
		x"ff",	--14924
		x"ff",	--14925
		x"ff",	--14926
		x"ff",	--14927
		x"ff",	--14928
		x"ff",	--14929
		x"ff",	--14930
		x"ff",	--14931
		x"ff",	--14932
		x"ff",	--14933
		x"ff",	--14934
		x"ff",	--14935
		x"ff",	--14936
		x"ff",	--14937
		x"ff",	--14938
		x"ff",	--14939
		x"ff",	--14940
		x"ff",	--14941
		x"ff",	--14942
		x"ff",	--14943
		x"ff",	--14944
		x"ff",	--14945
		x"ff",	--14946
		x"ff",	--14947
		x"ff",	--14948
		x"ff",	--14949
		x"ff",	--14950
		x"ff",	--14951
		x"ff",	--14952
		x"ff",	--14953
		x"ff",	--14954
		x"ff",	--14955
		x"ff",	--14956
		x"ff",	--14957
		x"ff",	--14958
		x"ff",	--14959
		x"ff",	--14960
		x"ff",	--14961
		x"ff",	--14962
		x"ff",	--14963
		x"ff",	--14964
		x"ff",	--14965
		x"ff",	--14966
		x"ff",	--14967
		x"ff",	--14968
		x"ff",	--14969
		x"ff",	--14970
		x"ff",	--14971
		x"ff",	--14972
		x"ff",	--14973
		x"ff",	--14974
		x"ff",	--14975
		x"ff",	--14976
		x"ff",	--14977
		x"ff",	--14978
		x"ff",	--14979
		x"ff",	--14980
		x"ff",	--14981
		x"ff",	--14982
		x"ff",	--14983
		x"ff",	--14984
		x"ff",	--14985
		x"ff",	--14986
		x"ff",	--14987
		x"ff",	--14988
		x"ff",	--14989
		x"ff",	--14990
		x"ff",	--14991
		x"ff",	--14992
		x"ff",	--14993
		x"ff",	--14994
		x"ff",	--14995
		x"ff",	--14996
		x"ff",	--14997
		x"ff",	--14998
		x"ff",	--14999
		x"ff",	--15000
		x"ff",	--15001
		x"ff",	--15002
		x"ff",	--15003
		x"ff",	--15004
		x"ff",	--15005
		x"ff",	--15006
		x"ff",	--15007
		x"ff",	--15008
		x"ff",	--15009
		x"ff",	--15010
		x"ff",	--15011
		x"ff",	--15012
		x"ff",	--15013
		x"ff",	--15014
		x"ff",	--15015
		x"ff",	--15016
		x"ff",	--15017
		x"ff",	--15018
		x"ff",	--15019
		x"ff",	--15020
		x"ff",	--15021
		x"ff",	--15022
		x"ff",	--15023
		x"ff",	--15024
		x"ff",	--15025
		x"ff",	--15026
		x"ff",	--15027
		x"ff",	--15028
		x"ff",	--15029
		x"ff",	--15030
		x"ff",	--15031
		x"ff",	--15032
		x"ff",	--15033
		x"ff",	--15034
		x"ff",	--15035
		x"ff",	--15036
		x"ff",	--15037
		x"ff",	--15038
		x"ff",	--15039
		x"ff",	--15040
		x"ff",	--15041
		x"ff",	--15042
		x"ff",	--15043
		x"ff",	--15044
		x"ff",	--15045
		x"ff",	--15046
		x"ff",	--15047
		x"ff",	--15048
		x"ff",	--15049
		x"ff",	--15050
		x"ff",	--15051
		x"ff",	--15052
		x"ff",	--15053
		x"ff",	--15054
		x"ff",	--15055
		x"ff",	--15056
		x"ff",	--15057
		x"ff",	--15058
		x"ff",	--15059
		x"ff",	--15060
		x"ff",	--15061
		x"ff",	--15062
		x"ff",	--15063
		x"ff",	--15064
		x"ff",	--15065
		x"ff",	--15066
		x"ff",	--15067
		x"ff",	--15068
		x"ff",	--15069
		x"ff",	--15070
		x"ff",	--15071
		x"ff",	--15072
		x"ff",	--15073
		x"ff",	--15074
		x"ff",	--15075
		x"ff",	--15076
		x"ff",	--15077
		x"ff",	--15078
		x"ff",	--15079
		x"ff",	--15080
		x"ff",	--15081
		x"ff",	--15082
		x"ff",	--15083
		x"ff",	--15084
		x"ff",	--15085
		x"ff",	--15086
		x"ff",	--15087
		x"ff",	--15088
		x"ff",	--15089
		x"ff",	--15090
		x"ff",	--15091
		x"ff",	--15092
		x"ff",	--15093
		x"ff",	--15094
		x"ff",	--15095
		x"ff",	--15096
		x"ff",	--15097
		x"ff",	--15098
		x"ff",	--15099
		x"ff",	--15100
		x"ff",	--15101
		x"ff",	--15102
		x"ff",	--15103
		x"ff",	--15104
		x"ff",	--15105
		x"ff",	--15106
		x"ff",	--15107
		x"ff",	--15108
		x"ff",	--15109
		x"ff",	--15110
		x"ff",	--15111
		x"ff",	--15112
		x"ff",	--15113
		x"ff",	--15114
		x"ff",	--15115
		x"ff",	--15116
		x"ff",	--15117
		x"ff",	--15118
		x"ff",	--15119
		x"ff",	--15120
		x"ff",	--15121
		x"ff",	--15122
		x"ff",	--15123
		x"ff",	--15124
		x"ff",	--15125
		x"ff",	--15126
		x"ff",	--15127
		x"ff",	--15128
		x"ff",	--15129
		x"ff",	--15130
		x"ff",	--15131
		x"ff",	--15132
		x"ff",	--15133
		x"ff",	--15134
		x"ff",	--15135
		x"ff",	--15136
		x"ff",	--15137
		x"ff",	--15138
		x"ff",	--15139
		x"ff",	--15140
		x"ff",	--15141
		x"ff",	--15142
		x"ff",	--15143
		x"ff",	--15144
		x"ff",	--15145
		x"ff",	--15146
		x"ff",	--15147
		x"ff",	--15148
		x"ff",	--15149
		x"ff",	--15150
		x"ff",	--15151
		x"ff",	--15152
		x"ff",	--15153
		x"ff",	--15154
		x"ff",	--15155
		x"ff",	--15156
		x"ff",	--15157
		x"ff",	--15158
		x"ff",	--15159
		x"ff",	--15160
		x"ff",	--15161
		x"ff",	--15162
		x"ff",	--15163
		x"ff",	--15164
		x"ff",	--15165
		x"ff",	--15166
		x"ff",	--15167
		x"ff",	--15168
		x"ff",	--15169
		x"ff",	--15170
		x"ff",	--15171
		x"ff",	--15172
		x"ff",	--15173
		x"ff",	--15174
		x"ff",	--15175
		x"ff",	--15176
		x"ff",	--15177
		x"ff",	--15178
		x"ff",	--15179
		x"ff",	--15180
		x"ff",	--15181
		x"ff",	--15182
		x"ff",	--15183
		x"ff",	--15184
		x"ff",	--15185
		x"ff",	--15186
		x"ff",	--15187
		x"ff",	--15188
		x"ff",	--15189
		x"ff",	--15190
		x"ff",	--15191
		x"ff",	--15192
		x"ff",	--15193
		x"ff",	--15194
		x"ff",	--15195
		x"ff",	--15196
		x"ff",	--15197
		x"ff",	--15198
		x"ff",	--15199
		x"ff",	--15200
		x"ff",	--15201
		x"ff",	--15202
		x"ff",	--15203
		x"ff",	--15204
		x"ff",	--15205
		x"ff",	--15206
		x"ff",	--15207
		x"ff",	--15208
		x"ff",	--15209
		x"ff",	--15210
		x"ff",	--15211
		x"ff",	--15212
		x"ff",	--15213
		x"ff",	--15214
		x"ff",	--15215
		x"ff",	--15216
		x"ff",	--15217
		x"ff",	--15218
		x"ff",	--15219
		x"ff",	--15220
		x"ff",	--15221
		x"ff",	--15222
		x"ff",	--15223
		x"ff",	--15224
		x"ff",	--15225
		x"ff",	--15226
		x"ff",	--15227
		x"ff",	--15228
		x"ff",	--15229
		x"ff",	--15230
		x"ff",	--15231
		x"ff",	--15232
		x"ff",	--15233
		x"ff",	--15234
		x"ff",	--15235
		x"ff",	--15236
		x"ff",	--15237
		x"ff",	--15238
		x"ff",	--15239
		x"ff",	--15240
		x"ff",	--15241
		x"ff",	--15242
		x"ff",	--15243
		x"ff",	--15244
		x"ff",	--15245
		x"ff",	--15246
		x"ff",	--15247
		x"ff",	--15248
		x"ff",	--15249
		x"ff",	--15250
		x"ff",	--15251
		x"ff",	--15252
		x"ff",	--15253
		x"ff",	--15254
		x"ff",	--15255
		x"ff",	--15256
		x"ff",	--15257
		x"ff",	--15258
		x"ff",	--15259
		x"ff",	--15260
		x"ff",	--15261
		x"ff",	--15262
		x"ff",	--15263
		x"ff",	--15264
		x"ff",	--15265
		x"ff",	--15266
		x"ff",	--15267
		x"ff",	--15268
		x"ff",	--15269
		x"ff",	--15270
		x"ff",	--15271
		x"ff",	--15272
		x"ff",	--15273
		x"ff",	--15274
		x"ff",	--15275
		x"ff",	--15276
		x"ff",	--15277
		x"ff",	--15278
		x"ff",	--15279
		x"ff",	--15280
		x"ff",	--15281
		x"ff",	--15282
		x"ff",	--15283
		x"ff",	--15284
		x"ff",	--15285
		x"ff",	--15286
		x"ff",	--15287
		x"ff",	--15288
		x"ff",	--15289
		x"ff",	--15290
		x"ff",	--15291
		x"ff",	--15292
		x"ff",	--15293
		x"ff",	--15294
		x"ff",	--15295
		x"ff",	--15296
		x"ff",	--15297
		x"ff",	--15298
		x"ff",	--15299
		x"ff",	--15300
		x"ff",	--15301
		x"ff",	--15302
		x"ff",	--15303
		x"ff",	--15304
		x"ff",	--15305
		x"ff",	--15306
		x"ff",	--15307
		x"ff",	--15308
		x"ff",	--15309
		x"ff",	--15310
		x"ff",	--15311
		x"ff",	--15312
		x"ff",	--15313
		x"ff",	--15314
		x"ff",	--15315
		x"ff",	--15316
		x"ff",	--15317
		x"ff",	--15318
		x"ff",	--15319
		x"ff",	--15320
		x"ff",	--15321
		x"ff",	--15322
		x"ff",	--15323
		x"ff",	--15324
		x"ff",	--15325
		x"ff",	--15326
		x"ff",	--15327
		x"ff",	--15328
		x"ff",	--15329
		x"ff",	--15330
		x"ff",	--15331
		x"ff",	--15332
		x"ff",	--15333
		x"ff",	--15334
		x"ff",	--15335
		x"ff",	--15336
		x"ff",	--15337
		x"ff",	--15338
		x"ff",	--15339
		x"ff",	--15340
		x"ff",	--15341
		x"ff",	--15342
		x"ff",	--15343
		x"ff",	--15344
		x"ff",	--15345
		x"ff",	--15346
		x"ff",	--15347
		x"ff",	--15348
		x"ff",	--15349
		x"ff",	--15350
		x"ff",	--15351
		x"ff",	--15352
		x"ff",	--15353
		x"ff",	--15354
		x"ff",	--15355
		x"ff",	--15356
		x"ff",	--15357
		x"ff",	--15358
		x"ff",	--15359
		x"ff",	--15360
		x"ff",	--15361
		x"ff",	--15362
		x"ff",	--15363
		x"ff",	--15364
		x"ff",	--15365
		x"ff",	--15366
		x"ff",	--15367
		x"ff",	--15368
		x"ff",	--15369
		x"ff",	--15370
		x"ff",	--15371
		x"ff",	--15372
		x"ff",	--15373
		x"ff",	--15374
		x"ff",	--15375
		x"ff",	--15376
		x"ff",	--15377
		x"ff",	--15378
		x"ff",	--15379
		x"ff",	--15380
		x"ff",	--15381
		x"ff",	--15382
		x"ff",	--15383
		x"ff",	--15384
		x"ff",	--15385
		x"ff",	--15386
		x"ff",	--15387
		x"ff",	--15388
		x"ff",	--15389
		x"ff",	--15390
		x"ff",	--15391
		x"ff",	--15392
		x"ff",	--15393
		x"ff",	--15394
		x"ff",	--15395
		x"ff",	--15396
		x"ff",	--15397
		x"ff",	--15398
		x"ff",	--15399
		x"ff",	--15400
		x"ff",	--15401
		x"ff",	--15402
		x"ff",	--15403
		x"ff",	--15404
		x"ff",	--15405
		x"ff",	--15406
		x"ff",	--15407
		x"ff",	--15408
		x"ff",	--15409
		x"ff",	--15410
		x"ff",	--15411
		x"ff",	--15412
		x"ff",	--15413
		x"ff",	--15414
		x"ff",	--15415
		x"ff",	--15416
		x"ff",	--15417
		x"ff",	--15418
		x"ff",	--15419
		x"ff",	--15420
		x"ff",	--15421
		x"ff",	--15422
		x"ff",	--15423
		x"ff",	--15424
		x"ff",	--15425
		x"ff",	--15426
		x"ff",	--15427
		x"ff",	--15428
		x"ff",	--15429
		x"ff",	--15430
		x"ff",	--15431
		x"ff",	--15432
		x"ff",	--15433
		x"ff",	--15434
		x"ff",	--15435
		x"ff",	--15436
		x"ff",	--15437
		x"ff",	--15438
		x"ff",	--15439
		x"ff",	--15440
		x"ff",	--15441
		x"ff",	--15442
		x"ff",	--15443
		x"ff",	--15444
		x"ff",	--15445
		x"ff",	--15446
		x"ff",	--15447
		x"ff",	--15448
		x"ff",	--15449
		x"ff",	--15450
		x"ff",	--15451
		x"ff",	--15452
		x"ff",	--15453
		x"ff",	--15454
		x"ff",	--15455
		x"ff",	--15456
		x"ff",	--15457
		x"ff",	--15458
		x"ff",	--15459
		x"ff",	--15460
		x"ff",	--15461
		x"ff",	--15462
		x"ff",	--15463
		x"ff",	--15464
		x"ff",	--15465
		x"ff",	--15466
		x"ff",	--15467
		x"ff",	--15468
		x"ff",	--15469
		x"ff",	--15470
		x"ff",	--15471
		x"ff",	--15472
		x"ff",	--15473
		x"ff",	--15474
		x"ff",	--15475
		x"ff",	--15476
		x"ff",	--15477
		x"ff",	--15478
		x"ff",	--15479
		x"ff",	--15480
		x"ff",	--15481
		x"ff",	--15482
		x"ff",	--15483
		x"ff",	--15484
		x"ff",	--15485
		x"ff",	--15486
		x"ff",	--15487
		x"ff",	--15488
		x"ff",	--15489
		x"ff",	--15490
		x"ff",	--15491
		x"ff",	--15492
		x"ff",	--15493
		x"ff",	--15494
		x"ff",	--15495
		x"ff",	--15496
		x"ff",	--15497
		x"ff",	--15498
		x"ff",	--15499
		x"ff",	--15500
		x"ff",	--15501
		x"ff",	--15502
		x"ff",	--15503
		x"ff",	--15504
		x"ff",	--15505
		x"ff",	--15506
		x"ff",	--15507
		x"ff",	--15508
		x"ff",	--15509
		x"ff",	--15510
		x"ff",	--15511
		x"ff",	--15512
		x"ff",	--15513
		x"ff",	--15514
		x"ff",	--15515
		x"ff",	--15516
		x"ff",	--15517
		x"ff",	--15518
		x"ff",	--15519
		x"ff",	--15520
		x"ff",	--15521
		x"ff",	--15522
		x"ff",	--15523
		x"ff",	--15524
		x"ff",	--15525
		x"ff",	--15526
		x"ff",	--15527
		x"ff",	--15528
		x"ff",	--15529
		x"ff",	--15530
		x"ff",	--15531
		x"ff",	--15532
		x"ff",	--15533
		x"ff",	--15534
		x"ff",	--15535
		x"ff",	--15536
		x"ff",	--15537
		x"ff",	--15538
		x"ff",	--15539
		x"ff",	--15540
		x"ff",	--15541
		x"ff",	--15542
		x"ff",	--15543
		x"ff",	--15544
		x"ff",	--15545
		x"ff",	--15546
		x"ff",	--15547
		x"ff",	--15548
		x"ff",	--15549
		x"ff",	--15550
		x"ff",	--15551
		x"ff",	--15552
		x"ff",	--15553
		x"ff",	--15554
		x"ff",	--15555
		x"ff",	--15556
		x"ff",	--15557
		x"ff",	--15558
		x"ff",	--15559
		x"ff",	--15560
		x"ff",	--15561
		x"ff",	--15562
		x"ff",	--15563
		x"ff",	--15564
		x"ff",	--15565
		x"ff",	--15566
		x"ff",	--15567
		x"ff",	--15568
		x"ff",	--15569
		x"ff",	--15570
		x"ff",	--15571
		x"ff",	--15572
		x"ff",	--15573
		x"ff",	--15574
		x"ff",	--15575
		x"ff",	--15576
		x"ff",	--15577
		x"ff",	--15578
		x"ff",	--15579
		x"ff",	--15580
		x"ff",	--15581
		x"ff",	--15582
		x"ff",	--15583
		x"ff",	--15584
		x"ff",	--15585
		x"ff",	--15586
		x"ff",	--15587
		x"ff",	--15588
		x"ff",	--15589
		x"ff",	--15590
		x"ff",	--15591
		x"ff",	--15592
		x"ff",	--15593
		x"ff",	--15594
		x"ff",	--15595
		x"ff",	--15596
		x"ff",	--15597
		x"ff",	--15598
		x"ff",	--15599
		x"ff",	--15600
		x"ff",	--15601
		x"ff",	--15602
		x"ff",	--15603
		x"ff",	--15604
		x"ff",	--15605
		x"ff",	--15606
		x"ff",	--15607
		x"ff",	--15608
		x"ff",	--15609
		x"ff",	--15610
		x"ff",	--15611
		x"ff",	--15612
		x"ff",	--15613
		x"ff",	--15614
		x"ff",	--15615
		x"ff",	--15616
		x"ff",	--15617
		x"ff",	--15618
		x"ff",	--15619
		x"ff",	--15620
		x"ff",	--15621
		x"ff",	--15622
		x"ff",	--15623
		x"ff",	--15624
		x"ff",	--15625
		x"ff",	--15626
		x"ff",	--15627
		x"ff",	--15628
		x"ff",	--15629
		x"ff",	--15630
		x"ff",	--15631
		x"ff",	--15632
		x"ff",	--15633
		x"ff",	--15634
		x"ff",	--15635
		x"ff",	--15636
		x"ff",	--15637
		x"ff",	--15638
		x"ff",	--15639
		x"ff",	--15640
		x"ff",	--15641
		x"ff",	--15642
		x"ff",	--15643
		x"ff",	--15644
		x"ff",	--15645
		x"ff",	--15646
		x"ff",	--15647
		x"ff",	--15648
		x"ff",	--15649
		x"ff",	--15650
		x"ff",	--15651
		x"ff",	--15652
		x"ff",	--15653
		x"ff",	--15654
		x"ff",	--15655
		x"ff",	--15656
		x"ff",	--15657
		x"ff",	--15658
		x"ff",	--15659
		x"ff",	--15660
		x"ff",	--15661
		x"ff",	--15662
		x"ff",	--15663
		x"ff",	--15664
		x"ff",	--15665
		x"ff",	--15666
		x"ff",	--15667
		x"ff",	--15668
		x"ff",	--15669
		x"ff",	--15670
		x"ff",	--15671
		x"ff",	--15672
		x"ff",	--15673
		x"ff",	--15674
		x"ff",	--15675
		x"ff",	--15676
		x"ff",	--15677
		x"ff",	--15678
		x"ff",	--15679
		x"ff",	--15680
		x"ff",	--15681
		x"ff",	--15682
		x"ff",	--15683
		x"ff",	--15684
		x"ff",	--15685
		x"ff",	--15686
		x"ff",	--15687
		x"ff",	--15688
		x"ff",	--15689
		x"ff",	--15690
		x"ff",	--15691
		x"ff",	--15692
		x"ff",	--15693
		x"ff",	--15694
		x"ff",	--15695
		x"ff",	--15696
		x"ff",	--15697
		x"ff",	--15698
		x"ff",	--15699
		x"ff",	--15700
		x"ff",	--15701
		x"ff",	--15702
		x"ff",	--15703
		x"ff",	--15704
		x"ff",	--15705
		x"ff",	--15706
		x"ff",	--15707
		x"ff",	--15708
		x"ff",	--15709
		x"ff",	--15710
		x"ff",	--15711
		x"ff",	--15712
		x"ff",	--15713
		x"ff",	--15714
		x"ff",	--15715
		x"ff",	--15716
		x"ff",	--15717
		x"ff",	--15718
		x"ff",	--15719
		x"ff",	--15720
		x"ff",	--15721
		x"ff",	--15722
		x"ff",	--15723
		x"ff",	--15724
		x"ff",	--15725
		x"ff",	--15726
		x"ff",	--15727
		x"ff",	--15728
		x"ff",	--15729
		x"ff",	--15730
		x"ff",	--15731
		x"ff",	--15732
		x"ff",	--15733
		x"ff",	--15734
		x"ff",	--15735
		x"ff",	--15736
		x"ff",	--15737
		x"ff",	--15738
		x"ff",	--15739
		x"ff",	--15740
		x"ff",	--15741
		x"ff",	--15742
		x"ff",	--15743
		x"ff",	--15744
		x"ff",	--15745
		x"ff",	--15746
		x"ff",	--15747
		x"ff",	--15748
		x"ff",	--15749
		x"ff",	--15750
		x"ff",	--15751
		x"ff",	--15752
		x"ff",	--15753
		x"ff",	--15754
		x"ff",	--15755
		x"ff",	--15756
		x"ff",	--15757
		x"ff",	--15758
		x"ff",	--15759
		x"ff",	--15760
		x"ff",	--15761
		x"ff",	--15762
		x"ff",	--15763
		x"ff",	--15764
		x"ff",	--15765
		x"ff",	--15766
		x"ff",	--15767
		x"ff",	--15768
		x"ff",	--15769
		x"ff",	--15770
		x"ff",	--15771
		x"ff",	--15772
		x"ff",	--15773
		x"ff",	--15774
		x"ff",	--15775
		x"ff",	--15776
		x"ff",	--15777
		x"ff",	--15778
		x"ff",	--15779
		x"ff",	--15780
		x"ff",	--15781
		x"ff",	--15782
		x"ff",	--15783
		x"ff",	--15784
		x"ff",	--15785
		x"ff",	--15786
		x"ff",	--15787
		x"ff",	--15788
		x"ff",	--15789
		x"ff",	--15790
		x"ff",	--15791
		x"ff",	--15792
		x"ff",	--15793
		x"ff",	--15794
		x"ff",	--15795
		x"ff",	--15796
		x"ff",	--15797
		x"ff",	--15798
		x"ff",	--15799
		x"ff",	--15800
		x"ff",	--15801
		x"ff",	--15802
		x"ff",	--15803
		x"ff",	--15804
		x"ff",	--15805
		x"ff",	--15806
		x"ff",	--15807
		x"ff",	--15808
		x"ff",	--15809
		x"ff",	--15810
		x"ff",	--15811
		x"ff",	--15812
		x"ff",	--15813
		x"ff",	--15814
		x"ff",	--15815
		x"ff",	--15816
		x"ff",	--15817
		x"ff",	--15818
		x"ff",	--15819
		x"ff",	--15820
		x"ff",	--15821
		x"ff",	--15822
		x"ff",	--15823
		x"ff",	--15824
		x"ff",	--15825
		x"ff",	--15826
		x"ff",	--15827
		x"ff",	--15828
		x"ff",	--15829
		x"ff",	--15830
		x"ff",	--15831
		x"ff",	--15832
		x"ff",	--15833
		x"ff",	--15834
		x"ff",	--15835
		x"ff",	--15836
		x"ff",	--15837
		x"ff",	--15838
		x"ff",	--15839
		x"ff",	--15840
		x"ff",	--15841
		x"ff",	--15842
		x"ff",	--15843
		x"ff",	--15844
		x"ff",	--15845
		x"ff",	--15846
		x"ff",	--15847
		x"ff",	--15848
		x"ff",	--15849
		x"ff",	--15850
		x"ff",	--15851
		x"ff",	--15852
		x"ff",	--15853
		x"ff",	--15854
		x"ff",	--15855
		x"ff",	--15856
		x"ff",	--15857
		x"ff",	--15858
		x"ff",	--15859
		x"ff",	--15860
		x"ff",	--15861
		x"ff",	--15862
		x"ff",	--15863
		x"ff",	--15864
		x"ff",	--15865
		x"ff",	--15866
		x"ff",	--15867
		x"ff",	--15868
		x"ff",	--15869
		x"ff",	--15870
		x"ff",	--15871
		x"ff",	--15872
		x"ff",	--15873
		x"ff",	--15874
		x"ff",	--15875
		x"ff",	--15876
		x"ff",	--15877
		x"ff",	--15878
		x"ff",	--15879
		x"ff",	--15880
		x"ff",	--15881
		x"ff",	--15882
		x"ff",	--15883
		x"ff",	--15884
		x"ff",	--15885
		x"ff",	--15886
		x"ff",	--15887
		x"ff",	--15888
		x"ff",	--15889
		x"ff",	--15890
		x"ff",	--15891
		x"ff",	--15892
		x"ff",	--15893
		x"ff",	--15894
		x"ff",	--15895
		x"ff",	--15896
		x"ff",	--15897
		x"ff",	--15898
		x"ff",	--15899
		x"ff",	--15900
		x"ff",	--15901
		x"ff",	--15902
		x"ff",	--15903
		x"ff",	--15904
		x"ff",	--15905
		x"ff",	--15906
		x"ff",	--15907
		x"ff",	--15908
		x"ff",	--15909
		x"ff",	--15910
		x"ff",	--15911
		x"ff",	--15912
		x"ff",	--15913
		x"ff",	--15914
		x"ff",	--15915
		x"ff",	--15916
		x"ff",	--15917
		x"ff",	--15918
		x"ff",	--15919
		x"ff",	--15920
		x"ff",	--15921
		x"ff",	--15922
		x"ff",	--15923
		x"ff",	--15924
		x"ff",	--15925
		x"ff",	--15926
		x"ff",	--15927
		x"ff",	--15928
		x"ff",	--15929
		x"ff",	--15930
		x"ff",	--15931
		x"ff",	--15932
		x"ff",	--15933
		x"ff",	--15934
		x"ff",	--15935
		x"ff",	--15936
		x"ff",	--15937
		x"ff",	--15938
		x"ff",	--15939
		x"ff",	--15940
		x"ff",	--15941
		x"ff",	--15942
		x"ff",	--15943
		x"ff",	--15944
		x"ff",	--15945
		x"ff",	--15946
		x"ff",	--15947
		x"ff",	--15948
		x"ff",	--15949
		x"ff",	--15950
		x"ff",	--15951
		x"ff",	--15952
		x"ff",	--15953
		x"ff",	--15954
		x"ff",	--15955
		x"ff",	--15956
		x"ff",	--15957
		x"ff",	--15958
		x"ff",	--15959
		x"ff",	--15960
		x"ff",	--15961
		x"ff",	--15962
		x"ff",	--15963
		x"ff",	--15964
		x"ff",	--15965
		x"ff",	--15966
		x"ff",	--15967
		x"ff",	--15968
		x"ff",	--15969
		x"ff",	--15970
		x"ff",	--15971
		x"ff",	--15972
		x"ff",	--15973
		x"ff",	--15974
		x"ff",	--15975
		x"ff",	--15976
		x"ff",	--15977
		x"ff",	--15978
		x"ff",	--15979
		x"ff",	--15980
		x"ff",	--15981
		x"ff",	--15982
		x"ff",	--15983
		x"ff",	--15984
		x"ff",	--15985
		x"ff",	--15986
		x"ff",	--15987
		x"ff",	--15988
		x"ff",	--15989
		x"ff",	--15990
		x"ff",	--15991
		x"ff",	--15992
		x"ff",	--15993
		x"ff",	--15994
		x"ff",	--15995
		x"ff",	--15996
		x"ff",	--15997
		x"ff",	--15998
		x"ff",	--15999
		x"ff",	--16000
		x"ff",	--16001
		x"ff",	--16002
		x"ff",	--16003
		x"ff",	--16004
		x"ff",	--16005
		x"ff",	--16006
		x"ff",	--16007
		x"ff",	--16008
		x"ff",	--16009
		x"ff",	--16010
		x"ff",	--16011
		x"ff",	--16012
		x"ff",	--16013
		x"ff",	--16014
		x"ff",	--16015
		x"ff",	--16016
		x"ff",	--16017
		x"ff",	--16018
		x"ff",	--16019
		x"ff",	--16020
		x"ff",	--16021
		x"ff",	--16022
		x"ff",	--16023
		x"ff",	--16024
		x"ff",	--16025
		x"ff",	--16026
		x"ff",	--16027
		x"ff",	--16028
		x"ff",	--16029
		x"ff",	--16030
		x"ff",	--16031
		x"ff",	--16032
		x"ff",	--16033
		x"ff",	--16034
		x"ff",	--16035
		x"ff",	--16036
		x"ff",	--16037
		x"ff",	--16038
		x"ff",	--16039
		x"ff",	--16040
		x"ff",	--16041
		x"ff",	--16042
		x"ff",	--16043
		x"ff",	--16044
		x"ff",	--16045
		x"ff",	--16046
		x"ff",	--16047
		x"ff",	--16048
		x"ff",	--16049
		x"ff",	--16050
		x"ff",	--16051
		x"ff",	--16052
		x"ff",	--16053
		x"ff",	--16054
		x"ff",	--16055
		x"ff",	--16056
		x"ff",	--16057
		x"ff",	--16058
		x"ff",	--16059
		x"ff",	--16060
		x"ff",	--16061
		x"ff",	--16062
		x"ff",	--16063
		x"ff",	--16064
		x"ff",	--16065
		x"ff",	--16066
		x"ff",	--16067
		x"ff",	--16068
		x"ff",	--16069
		x"ff",	--16070
		x"ff",	--16071
		x"ff",	--16072
		x"ff",	--16073
		x"ff",	--16074
		x"ff",	--16075
		x"ff",	--16076
		x"ff",	--16077
		x"ff",	--16078
		x"ff",	--16079
		x"ff",	--16080
		x"ff",	--16081
		x"ff",	--16082
		x"ff",	--16083
		x"ff",	--16084
		x"ff",	--16085
		x"ff",	--16086
		x"ff",	--16087
		x"ff",	--16088
		x"ff",	--16089
		x"ff",	--16090
		x"ff",	--16091
		x"ff",	--16092
		x"ff",	--16093
		x"ff",	--16094
		x"ff",	--16095
		x"ff",	--16096
		x"ff",	--16097
		x"ff",	--16098
		x"ff",	--16099
		x"ff",	--16100
		x"ff",	--16101
		x"ff",	--16102
		x"ff",	--16103
		x"ff",	--16104
		x"ff",	--16105
		x"ff",	--16106
		x"ff",	--16107
		x"ff",	--16108
		x"ff",	--16109
		x"ff",	--16110
		x"ff",	--16111
		x"ff",	--16112
		x"ff",	--16113
		x"ff",	--16114
		x"ff",	--16115
		x"ff",	--16116
		x"ff",	--16117
		x"ff",	--16118
		x"ff",	--16119
		x"ff",	--16120
		x"ff",	--16121
		x"ff",	--16122
		x"ff",	--16123
		x"ff",	--16124
		x"ff",	--16125
		x"ff",	--16126
		x"ff",	--16127
		x"ff",	--16128
		x"ff",	--16129
		x"ff",	--16130
		x"ff",	--16131
		x"ff",	--16132
		x"ff",	--16133
		x"ff",	--16134
		x"ff",	--16135
		x"ff",	--16136
		x"ff",	--16137
		x"ff",	--16138
		x"ff",	--16139
		x"ff",	--16140
		x"ff",	--16141
		x"ff",	--16142
		x"ff",	--16143
		x"ff",	--16144
		x"ff",	--16145
		x"ff",	--16146
		x"ff",	--16147
		x"ff",	--16148
		x"ff",	--16149
		x"ff",	--16150
		x"ff",	--16151
		x"ff",	--16152
		x"ff",	--16153
		x"ff",	--16154
		x"ff",	--16155
		x"ff",	--16156
		x"ff",	--16157
		x"ff",	--16158
		x"ff",	--16159
		x"ff",	--16160
		x"ff",	--16161
		x"ff",	--16162
		x"ff",	--16163
		x"ff",	--16164
		x"ff",	--16165
		x"ff",	--16166
		x"ff",	--16167
		x"ff",	--16168
		x"ff",	--16169
		x"ff",	--16170
		x"ff",	--16171
		x"ff",	--16172
		x"ff",	--16173
		x"ff",	--16174
		x"ff",	--16175
		x"ff",	--16176
		x"ff",	--16177
		x"ff",	--16178
		x"ff",	--16179
		x"ff",	--16180
		x"ff",	--16181
		x"ff",	--16182
		x"ff",	--16183
		x"ff",	--16184
		x"ff",	--16185
		x"ff",	--16186
		x"ff",	--16187
		x"ff",	--16188
		x"ff",	--16189
		x"ff",	--16190
		x"ff",	--16191
		x"ff",	--16192
		x"ff",	--16193
		x"ff",	--16194
		x"ff",	--16195
		x"ff",	--16196
		x"ff",	--16197
		x"ff",	--16198
		x"ff",	--16199
		x"ff",	--16200
		x"ff",	--16201
		x"ff",	--16202
		x"ff",	--16203
		x"ff",	--16204
		x"ff",	--16205
		x"ff",	--16206
		x"ff",	--16207
		x"ff",	--16208
		x"ff",	--16209
		x"ff",	--16210
		x"ff",	--16211
		x"ff",	--16212
		x"ff",	--16213
		x"ff",	--16214
		x"ff",	--16215
		x"ff",	--16216
		x"ff",	--16217
		x"ff",	--16218
		x"ff",	--16219
		x"ff",	--16220
		x"ff",	--16221
		x"ff",	--16222
		x"ff",	--16223
		x"ff",	--16224
		x"ff",	--16225
		x"ff",	--16226
		x"ff",	--16227
		x"ff",	--16228
		x"ff",	--16229
		x"ff",	--16230
		x"ff",	--16231
		x"ff",	--16232
		x"ff",	--16233
		x"ff",	--16234
		x"ff",	--16235
		x"ff",	--16236
		x"ff",	--16237
		x"ff",	--16238
		x"ff",	--16239
		x"ff",	--16240
		x"ff",	--16241
		x"ff",	--16242
		x"ff",	--16243
		x"ff",	--16244
		x"ff",	--16245
		x"ff",	--16246
		x"ff",	--16247
		x"ff",	--16248
		x"ff",	--16249
		x"ff",	--16250
		x"ff",	--16251
		x"ff",	--16252
		x"ff",	--16253
		x"ff",	--16254
		x"ff",	--16255
		x"ff",	--16256
		x"ff",	--16257
		x"ff",	--16258
		x"ff",	--16259
		x"ff",	--16260
		x"ff",	--16261
		x"ff",	--16262
		x"ff",	--16263
		x"ff",	--16264
		x"ff",	--16265
		x"ff",	--16266
		x"ff",	--16267
		x"ff",	--16268
		x"ff",	--16269
		x"ff",	--16270
		x"ff",	--16271
		x"ff",	--16272
		x"ff",	--16273
		x"ff",	--16274
		x"ff",	--16275
		x"ff",	--16276
		x"ff",	--16277
		x"ff",	--16278
		x"ff",	--16279
		x"ff",	--16280
		x"ff",	--16281
		x"ff",	--16282
		x"ff",	--16283
		x"ff",	--16284
		x"ff",	--16285
		x"ff",	--16286
		x"ff",	--16287
		x"ff",	--16288
		x"ff",	--16289
		x"ff",	--16290
		x"ff",	--16291
		x"ff",	--16292
		x"ff",	--16293
		x"ff",	--16294
		x"ff",	--16295
		x"ff",	--16296
		x"ff",	--16297
		x"ff",	--16298
		x"ff",	--16299
		x"ff",	--16300
		x"ff",	--16301
		x"ff",	--16302
		x"ff",	--16303
		x"ff",	--16304
		x"ff",	--16305
		x"ff",	--16306
		x"ff",	--16307
		x"ff",	--16308
		x"ff",	--16309
		x"ff",	--16310
		x"ff",	--16311
		x"ff",	--16312
		x"ff",	--16313
		x"ff",	--16314
		x"ff",	--16315
		x"ff",	--16316
		x"ff",	--16317
		x"ff",	--16318
		x"ff",	--16319
		x"ff",	--16320
		x"ff",	--16321
		x"ff",	--16322
		x"ff",	--16323
		x"ff",	--16324
		x"ff",	--16325
		x"ff",	--16326
		x"ff",	--16327
		x"ff",	--16328
		x"ff",	--16329
		x"ff",	--16330
		x"ff",	--16331
		x"ff",	--16332
		x"ff",	--16333
		x"ff",	--16334
		x"ff",	--16335
		x"ff",	--16336
		x"ff",	--16337
		x"ff",	--16338
		x"ff",	--16339
		x"ff",	--16340
		x"ff",	--16341
		x"ff",	--16342
		x"ff",	--16343
		x"ff",	--16344
		x"ff",	--16345
		x"ff",	--16346
		x"ff",	--16347
		x"ff",	--16348
		x"ff",	--16349
		x"ff",	--16350
		x"ff",	--16351
		x"ff",	--16352
		x"ff",	--16353
		x"ff",	--16354
		x"ff",	--16355
		x"ff",	--16356
		x"ff",	--16357
		x"ff",	--16358
		x"ff",	--16359
		x"ff",	--16360
		x"ff",	--16361
		x"ff",	--16362
		x"ff",	--16363
		x"ff",	--16364
		x"ff",	--16365
		x"ff",	--16366
		x"ff",	--16367
		x"fc",	--16368
		x"fc",	--16369
		x"fc",	--16370
		x"fc",	--16371
		x"fc",	--16372
		x"fc",	--16373
		x"fc",	--16374
		x"8c",	--16375
		x"de",	--16376
		x"fc",	--16377
		x"fc",	--16378
		x"fc",	--16379
		x"fc",	--16380
		x"fc",	--16381
		x"fc",	--16382
		x"00");	--16383
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"dc",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"9c",	--44
		x"12",	--45
		x"97",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"d3",	--50
		x"12",	--51
		x"9b",	--52
		x"53",	--53
		x"40",	--54
		x"d4",	--55
		x"40",	--56
		x"85",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"97",	--61
		x"40",	--62
		x"d4",	--63
		x"40",	--64
		x"91",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"97",	--69
		x"40",	--70
		x"d4",	--71
		x"40",	--72
		x"91",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"97",	--77
		x"40",	--78
		x"d4",	--79
		x"40",	--80
		x"85",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"97",	--85
		x"40",	--86
		x"d4",	--87
		x"40",	--88
		x"8a",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"97",	--93
		x"40",	--94
		x"d4",	--95
		x"40",	--96
		x"8b",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"97",	--101
		x"40",	--102
		x"d4",	--103
		x"40",	--104
		x"86",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"97",	--109
		x"40",	--110
		x"d4",	--111
		x"40",	--112
		x"84",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"97",	--117
		x"40",	--118
		x"d4",	--119
		x"40",	--120
		x"87",	--121
		x"40",	--122
		x"00",	--123
		x"12",	--124
		x"97",	--125
		x"40",	--126
		x"d4",	--127
		x"40",	--128
		x"84",	--129
		x"40",	--130
		x"00",	--131
		x"12",	--132
		x"97",	--133
		x"40",	--134
		x"d4",	--135
		x"40",	--136
		x"8f",	--137
		x"40",	--138
		x"00",	--139
		x"12",	--140
		x"97",	--141
		x"40",	--142
		x"d4",	--143
		x"40",	--144
		x"87",	--145
		x"40",	--146
		x"00",	--147
		x"12",	--148
		x"97",	--149
		x"43",	--150
		x"43",	--151
		x"12",	--152
		x"96",	--153
		x"43",	--154
		x"40",	--155
		x"4e",	--156
		x"40",	--157
		x"01",	--158
		x"41",	--159
		x"50",	--160
		x"00",	--161
		x"12",	--162
		x"95",	--163
		x"41",	--164
		x"50",	--165
		x"00",	--166
		x"12",	--167
		x"96",	--168
		x"43",	--169
		x"40",	--170
		x"4e",	--171
		x"40",	--172
		x"01",	--173
		x"41",	--174
		x"52",	--175
		x"12",	--176
		x"95",	--177
		x"41",	--178
		x"52",	--179
		x"12",	--180
		x"96",	--181
		x"41",	--182
		x"52",	--183
		x"41",	--184
		x"50",	--185
		x"00",	--186
		x"12",	--187
		x"8a",	--188
		x"40",	--189
		x"01",	--190
		x"41",	--191
		x"50",	--192
		x"00",	--193
		x"12",	--194
		x"99",	--195
		x"40",	--196
		x"01",	--197
		x"41",	--198
		x"52",	--199
		x"12",	--200
		x"99",	--201
		x"41",	--202
		x"52",	--203
		x"41",	--204
		x"50",	--205
		x"00",	--206
		x"12",	--207
		x"8b",	--208
		x"41",	--209
		x"52",	--210
		x"41",	--211
		x"50",	--212
		x"00",	--213
		x"12",	--214
		x"8b",	--215
		x"12",	--216
		x"98",	--217
		x"40",	--218
		x"01",	--219
		x"41",	--220
		x"53",	--221
		x"12",	--222
		x"99",	--223
		x"41",	--224
		x"53",	--225
		x"12",	--226
		x"85",	--227
		x"40",	--228
		x"00",	--229
		x"40",	--230
		x"11",	--231
		x"41",	--232
		x"53",	--233
		x"12",	--234
		x"99",	--235
		x"40",	--236
		x"01",	--237
		x"41",	--238
		x"12",	--239
		x"98",	--240
		x"41",	--241
		x"12",	--242
		x"84",	--243
		x"12",	--244
		x"41",	--245
		x"12",	--246
		x"12",	--247
		x"12",	--248
		x"12",	--249
		x"39",	--250
		x"12",	--251
		x"b7",	--252
		x"12",	--253
		x"3a",	--254
		x"12",	--255
		x"49",	--256
		x"40",	--257
		x"00",	--258
		x"41",	--259
		x"50",	--260
		x"00",	--261
		x"41",	--262
		x"50",	--263
		x"00",	--264
		x"41",	--265
		x"50",	--266
		x"00",	--267
		x"12",	--268
		x"89",	--269
		x"50",	--270
		x"00",	--271
		x"12",	--272
		x"41",	--273
		x"12",	--274
		x"12",	--275
		x"12",	--276
		x"12",	--277
		x"39",	--278
		x"12",	--279
		x"b7",	--280
		x"12",	--281
		x"3a",	--282
		x"12",	--283
		x"49",	--284
		x"40",	--285
		x"00",	--286
		x"41",	--287
		x"50",	--288
		x"00",	--289
		x"41",	--290
		x"50",	--291
		x"00",	--292
		x"41",	--293
		x"50",	--294
		x"00",	--295
		x"12",	--296
		x"89",	--297
		x"50",	--298
		x"00",	--299
		x"41",	--300
		x"50",	--301
		x"00",	--302
		x"41",	--303
		x"50",	--304
		x"00",	--305
		x"12",	--306
		x"86",	--307
		x"41",	--308
		x"12",	--309
		x"86",	--310
		x"12",	--311
		x"86",	--312
		x"12",	--313
		x"04",	--314
		x"12",	--315
		x"3e",	--316
		x"12",	--317
		x"99",	--318
		x"40",	--319
		x"c2",	--320
		x"40",	--321
		x"3d",	--322
		x"41",	--323
		x"50",	--324
		x"00",	--325
		x"12",	--326
		x"92",	--327
		x"50",	--328
		x"00",	--329
		x"41",	--330
		x"50",	--331
		x"00",	--332
		x"41",	--333
		x"52",	--334
		x"41",	--335
		x"50",	--336
		x"00",	--337
		x"12",	--338
		x"93",	--339
		x"40",	--340
		x"00",	--341
		x"41",	--342
		x"50",	--343
		x"00",	--344
		x"12",	--345
		x"95",	--346
		x"41",	--347
		x"50",	--348
		x"00",	--349
		x"12",	--350
		x"84",	--351
		x"41",	--352
		x"50",	--353
		x"00",	--354
		x"41",	--355
		x"50",	--356
		x"00",	--357
		x"12",	--358
		x"8f",	--359
		x"41",	--360
		x"12",	--361
		x"8f",	--362
		x"40",	--363
		x"00",	--364
		x"12",	--365
		x"8f",	--366
		x"40",	--367
		x"ff",	--368
		x"00",	--369
		x"d2",	--370
		x"43",	--371
		x"43",	--372
		x"3c",	--373
		x"43",	--374
		x"3c",	--375
		x"43",	--376
		x"3c",	--377
		x"43",	--378
		x"12",	--379
		x"9c",	--380
		x"93",	--381
		x"27",	--382
		x"12",	--383
		x"9d",	--384
		x"93",	--385
		x"20",	--386
		x"90",	--387
		x"00",	--388
		x"24",	--389
		x"90",	--390
		x"00",	--391
		x"27",	--392
		x"92",	--393
		x"20",	--394
		x"3c",	--395
		x"12",	--396
		x"d4",	--397
		x"12",	--398
		x"9b",	--399
		x"53",	--400
		x"40",	--401
		x"00",	--402
		x"51",	--403
		x"5f",	--404
		x"43",	--405
		x"00",	--406
		x"4f",	--407
		x"41",	--408
		x"00",	--409
		x"12",	--410
		x"97",	--411
		x"43",	--412
		x"3f",	--413
		x"93",	--414
		x"27",	--415
		x"53",	--416
		x"12",	--417
		x"d4",	--418
		x"12",	--419
		x"9b",	--420
		x"53",	--421
		x"3f",	--422
		x"90",	--423
		x"00",	--424
		x"2f",	--425
		x"93",	--426
		x"02",	--427
		x"24",	--428
		x"4f",	--429
		x"11",	--430
		x"12",	--431
		x"12",	--432
		x"d4",	--433
		x"4f",	--434
		x"00",	--435
		x"12",	--436
		x"9b",	--437
		x"52",	--438
		x"41",	--439
		x"00",	--440
		x"40",	--441
		x"00",	--442
		x"51",	--443
		x"5a",	--444
		x"4f",	--445
		x"00",	--446
		x"53",	--447
		x"3f",	--448
		x"93",	--449
		x"20",	--450
		x"90",	--451
		x"00",	--452
		x"23",	--453
		x"3f",	--454
		x"93",	--455
		x"23",	--456
		x"90",	--457
		x"00",	--458
		x"24",	--459
		x"90",	--460
		x"00",	--461
		x"34",	--462
		x"90",	--463
		x"00",	--464
		x"23",	--465
		x"3c",	--466
		x"90",	--467
		x"00",	--468
		x"24",	--469
		x"90",	--470
		x"00",	--471
		x"23",	--472
		x"3c",	--473
		x"12",	--474
		x"d4",	--475
		x"12",	--476
		x"9b",	--477
		x"53",	--478
		x"12",	--479
		x"86",	--480
		x"43",	--481
		x"3f",	--482
		x"12",	--483
		x"d4",	--484
		x"12",	--485
		x"9b",	--486
		x"53",	--487
		x"12",	--488
		x"87",	--489
		x"43",	--490
		x"3f",	--491
		x"12",	--492
		x"d4",	--493
		x"12",	--494
		x"9b",	--495
		x"53",	--496
		x"12",	--497
		x"87",	--498
		x"43",	--499
		x"3f",	--500
		x"12",	--501
		x"d4",	--502
		x"12",	--503
		x"9b",	--504
		x"53",	--505
		x"12",	--506
		x"87",	--507
		x"43",	--508
		x"3f",	--509
		x"40",	--510
		x"d3",	--511
		x"4f",	--512
		x"02",	--513
		x"41",	--514
		x"12",	--515
		x"42",	--516
		x"02",	--517
		x"43",	--518
		x"40",	--519
		x"44",	--520
		x"4b",	--521
		x"00",	--522
		x"4b",	--523
		x"00",	--524
		x"12",	--525
		x"bd",	--526
		x"12",	--527
		x"c3",	--528
		x"12",	--529
		x"43",	--530
		x"40",	--531
		x"44",	--532
		x"4b",	--533
		x"00",	--534
		x"4b",	--535
		x"00",	--536
		x"12",	--537
		x"bd",	--538
		x"12",	--539
		x"c3",	--540
		x"12",	--541
		x"43",	--542
		x"40",	--543
		x"44",	--544
		x"4b",	--545
		x"00",	--546
		x"4b",	--547
		x"00",	--548
		x"12",	--549
		x"bd",	--550
		x"12",	--551
		x"c3",	--552
		x"12",	--553
		x"12",	--554
		x"d3",	--555
		x"12",	--556
		x"02",	--557
		x"12",	--558
		x"c9",	--559
		x"50",	--560
		x"00",	--561
		x"12",	--562
		x"02",	--563
		x"12",	--564
		x"d3",	--565
		x"12",	--566
		x"9b",	--567
		x"52",	--568
		x"43",	--569
		x"41",	--570
		x"41",	--571
		x"12",	--572
		x"43",	--573
		x"4b",	--574
		x"42",	--575
		x"02",	--576
		x"12",	--577
		x"98",	--578
		x"12",	--579
		x"12",	--580
		x"d3",	--581
		x"12",	--582
		x"9b",	--583
		x"52",	--584
		x"53",	--585
		x"90",	--586
		x"00",	--587
		x"23",	--588
		x"12",	--589
		x"d3",	--590
		x"12",	--591
		x"9b",	--592
		x"53",	--593
		x"41",	--594
		x"41",	--595
		x"4f",	--596
		x"02",	--597
		x"41",	--598
		x"12",	--599
		x"83",	--600
		x"4e",	--601
		x"43",	--602
		x"00",	--603
		x"93",	--604
		x"24",	--605
		x"93",	--606
		x"02",	--607
		x"24",	--608
		x"43",	--609
		x"02",	--610
		x"41",	--611
		x"4b",	--612
		x"00",	--613
		x"12",	--614
		x"87",	--615
		x"43",	--616
		x"4f",	--617
		x"42",	--618
		x"02",	--619
		x"12",	--620
		x"98",	--621
		x"43",	--622
		x"53",	--623
		x"41",	--624
		x"41",	--625
		x"93",	--626
		x"02",	--627
		x"24",	--628
		x"43",	--629
		x"02",	--630
		x"42",	--631
		x"02",	--632
		x"12",	--633
		x"98",	--634
		x"43",	--635
		x"53",	--636
		x"41",	--637
		x"41",	--638
		x"43",	--639
		x"12",	--640
		x"84",	--641
		x"43",	--642
		x"53",	--643
		x"41",	--644
		x"41",	--645
		x"43",	--646
		x"40",	--647
		x"84",	--648
		x"12",	--649
		x"98",	--650
		x"4f",	--651
		x"02",	--652
		x"3f",	--653
		x"4f",	--654
		x"02",	--655
		x"41",	--656
		x"12",	--657
		x"12",	--658
		x"82",	--659
		x"4f",	--660
		x"4e",	--661
		x"93",	--662
		x"38",	--663
		x"41",	--664
		x"4b",	--665
		x"00",	--666
		x"12",	--667
		x"87",	--668
		x"4f",	--669
		x"93",	--670
		x"24",	--671
		x"41",	--672
		x"4b",	--673
		x"00",	--674
		x"4d",	--675
		x"00",	--676
		x"12",	--677
		x"87",	--678
		x"4f",	--679
		x"41",	--680
		x"00",	--681
		x"42",	--682
		x"02",	--683
		x"12",	--684
		x"99",	--685
		x"43",	--686
		x"52",	--687
		x"41",	--688
		x"41",	--689
		x"41",	--690
		x"40",	--691
		x"00",	--692
		x"40",	--693
		x"11",	--694
		x"3f",	--695
		x"40",	--696
		x"11",	--697
		x"3f",	--698
		x"43",	--699
		x"93",	--700
		x"02",	--701
		x"24",	--702
		x"43",	--703
		x"4f",	--704
		x"02",	--705
		x"43",	--706
		x"41",	--707
		x"42",	--708
		x"00",	--709
		x"4e",	--710
		x"be",	--711
		x"20",	--712
		x"df",	--713
		x"00",	--714
		x"41",	--715
		x"cf",	--716
		x"00",	--717
		x"41",	--718
		x"42",	--719
		x"02",	--720
		x"92",	--721
		x"2c",	--722
		x"4e",	--723
		x"5f",	--724
		x"4f",	--725
		x"d3",	--726
		x"43",	--727
		x"00",	--728
		x"90",	--729
		x"00",	--730
		x"38",	--731
		x"43",	--732
		x"02",	--733
		x"41",	--734
		x"53",	--735
		x"4e",	--736
		x"02",	--737
		x"41",	--738
		x"40",	--739
		x"00",	--740
		x"00",	--741
		x"3f",	--742
		x"40",	--743
		x"00",	--744
		x"00",	--745
		x"3f",	--746
		x"42",	--747
		x"00",	--748
		x"3f",	--749
		x"40",	--750
		x"00",	--751
		x"00",	--752
		x"3f",	--753
		x"40",	--754
		x"00",	--755
		x"00",	--756
		x"3f",	--757
		x"40",	--758
		x"00",	--759
		x"00",	--760
		x"3f",	--761
		x"40",	--762
		x"00",	--763
		x"00",	--764
		x"3f",	--765
		x"43",	--766
		x"42",	--767
		x"02",	--768
		x"12",	--769
		x"8a",	--770
		x"43",	--771
		x"42",	--772
		x"02",	--773
		x"12",	--774
		x"8a",	--775
		x"12",	--776
		x"d4",	--777
		x"12",	--778
		x"9b",	--779
		x"53",	--780
		x"41",	--781
		x"93",	--782
		x"02",	--783
		x"24",	--784
		x"42",	--785
		x"02",	--786
		x"12",	--787
		x"89",	--788
		x"42",	--789
		x"02",	--790
		x"12",	--791
		x"89",	--792
		x"41",	--793
		x"43",	--794
		x"40",	--795
		x"85",	--796
		x"12",	--797
		x"98",	--798
		x"4f",	--799
		x"02",	--800
		x"3f",	--801
		x"4f",	--802
		x"02",	--803
		x"4e",	--804
		x"02",	--805
		x"41",	--806
		x"4f",	--807
		x"02",	--808
		x"41",	--809
		x"12",	--810
		x"12",	--811
		x"83",	--812
		x"4e",	--813
		x"90",	--814
		x"00",	--815
		x"38",	--816
		x"20",	--817
		x"41",	--818
		x"4b",	--819
		x"00",	--820
		x"12",	--821
		x"88",	--822
		x"4f",	--823
		x"41",	--824
		x"4b",	--825
		x"00",	--826
		x"12",	--827
		x"88",	--828
		x"4f",	--829
		x"12",	--830
		x"12",	--831
		x"12",	--832
		x"d4",	--833
		x"12",	--834
		x"9b",	--835
		x"50",	--836
		x"00",	--837
		x"4a",	--838
		x"42",	--839
		x"02",	--840
		x"12",	--841
		x"8a",	--842
		x"4b",	--843
		x"42",	--844
		x"02",	--845
		x"12",	--846
		x"8a",	--847
		x"43",	--848
		x"53",	--849
		x"41",	--850
		x"41",	--851
		x"41",	--852
		x"41",	--853
		x"4b",	--854
		x"00",	--855
		x"12",	--856
		x"87",	--857
		x"43",	--858
		x"4f",	--859
		x"42",	--860
		x"02",	--861
		x"12",	--862
		x"98",	--863
		x"3f",	--864
		x"12",	--865
		x"d4",	--866
		x"12",	--867
		x"9b",	--868
		x"4b",	--869
		x"00",	--870
		x"12",	--871
		x"d4",	--872
		x"12",	--873
		x"9b",	--874
		x"52",	--875
		x"43",	--876
		x"3f",	--877
		x"40",	--878
		x"00",	--879
		x"42",	--880
		x"02",	--881
		x"12",	--882
		x"8a",	--883
		x"40",	--884
		x"ff",	--885
		x"42",	--886
		x"02",	--887
		x"12",	--888
		x"8a",	--889
		x"43",	--890
		x"40",	--891
		x"00",	--892
		x"42",	--893
		x"02",	--894
		x"12",	--895
		x"98",	--896
		x"41",	--897
		x"40",	--898
		x"ff",	--899
		x"42",	--900
		x"02",	--901
		x"12",	--902
		x"8a",	--903
		x"40",	--904
		x"00",	--905
		x"42",	--906
		x"02",	--907
		x"12",	--908
		x"8a",	--909
		x"43",	--910
		x"40",	--911
		x"00",	--912
		x"42",	--913
		x"02",	--914
		x"12",	--915
		x"98",	--916
		x"41",	--917
		x"40",	--918
		x"ff",	--919
		x"42",	--920
		x"02",	--921
		x"12",	--922
		x"8a",	--923
		x"40",	--924
		x"ff",	--925
		x"42",	--926
		x"02",	--927
		x"12",	--928
		x"8a",	--929
		x"43",	--930
		x"40",	--931
		x"00",	--932
		x"42",	--933
		x"02",	--934
		x"12",	--935
		x"98",	--936
		x"41",	--937
		x"40",	--938
		x"00",	--939
		x"42",	--940
		x"02",	--941
		x"12",	--942
		x"8a",	--943
		x"40",	--944
		x"00",	--945
		x"42",	--946
		x"02",	--947
		x"12",	--948
		x"8a",	--949
		x"43",	--950
		x"40",	--951
		x"00",	--952
		x"42",	--953
		x"02",	--954
		x"12",	--955
		x"98",	--956
		x"41",	--957
		x"12",	--958
		x"d4",	--959
		x"12",	--960
		x"9b",	--961
		x"53",	--962
		x"43",	--963
		x"41",	--964
		x"40",	--965
		x"80",	--966
		x"01",	--967
		x"40",	--968
		x"00",	--969
		x"01",	--970
		x"40",	--971
		x"02",	--972
		x"01",	--973
		x"12",	--974
		x"d4",	--975
		x"12",	--976
		x"9b",	--977
		x"43",	--978
		x"01",	--979
		x"40",	--980
		x"d5",	--981
		x"00",	--982
		x"12",	--983
		x"9b",	--984
		x"53",	--985
		x"43",	--986
		x"41",	--987
		x"12",	--988
		x"12",	--989
		x"43",	--990
		x"00",	--991
		x"4f",	--992
		x"93",	--993
		x"24",	--994
		x"53",	--995
		x"43",	--996
		x"43",	--997
		x"3c",	--998
		x"90",	--999
		x"00",	--1000
		x"2c",	--1001
		x"5c",	--1002
		x"5c",	--1003
		x"5c",	--1004
		x"5c",	--1005
		x"11",	--1006
		x"5d",	--1007
		x"50",	--1008
		x"ff",	--1009
		x"43",	--1010
		x"4f",	--1011
		x"93",	--1012
		x"24",	--1013
		x"90",	--1014
		x"00",	--1015
		x"24",	--1016
		x"4d",	--1017
		x"50",	--1018
		x"ff",	--1019
		x"93",	--1020
		x"23",	--1021
		x"90",	--1022
		x"00",	--1023
		x"2c",	--1024
		x"5c",	--1025
		x"4c",	--1026
		x"5b",	--1027
		x"5b",	--1028
		x"5b",	--1029
		x"11",	--1030
		x"5d",	--1031
		x"50",	--1032
		x"ff",	--1033
		x"4f",	--1034
		x"93",	--1035
		x"23",	--1036
		x"43",	--1037
		x"00",	--1038
		x"4c",	--1039
		x"41",	--1040
		x"41",	--1041
		x"41",	--1042
		x"43",	--1043
		x"3f",	--1044
		x"4d",	--1045
		x"50",	--1046
		x"ff",	--1047
		x"90",	--1048
		x"00",	--1049
		x"2c",	--1050
		x"5c",	--1051
		x"5c",	--1052
		x"5c",	--1053
		x"5c",	--1054
		x"11",	--1055
		x"5d",	--1056
		x"50",	--1057
		x"ff",	--1058
		x"43",	--1059
		x"3f",	--1060
		x"4d",	--1061
		x"50",	--1062
		x"ff",	--1063
		x"90",	--1064
		x"00",	--1065
		x"2c",	--1066
		x"5c",	--1067
		x"5c",	--1068
		x"5c",	--1069
		x"5c",	--1070
		x"11",	--1071
		x"5d",	--1072
		x"50",	--1073
		x"ff",	--1074
		x"43",	--1075
		x"3f",	--1076
		x"11",	--1077
		x"12",	--1078
		x"12",	--1079
		x"d5",	--1080
		x"12",	--1081
		x"9b",	--1082
		x"52",	--1083
		x"43",	--1084
		x"4c",	--1085
		x"41",	--1086
		x"41",	--1087
		x"41",	--1088
		x"43",	--1089
		x"3f",	--1090
		x"12",	--1091
		x"12",	--1092
		x"43",	--1093
		x"00",	--1094
		x"4f",	--1095
		x"93",	--1096
		x"24",	--1097
		x"53",	--1098
		x"43",	--1099
		x"43",	--1100
		x"3c",	--1101
		x"4b",	--1102
		x"50",	--1103
		x"ff",	--1104
		x"90",	--1105
		x"00",	--1106
		x"2c",	--1107
		x"5c",	--1108
		x"4c",	--1109
		x"5d",	--1110
		x"5d",	--1111
		x"5d",	--1112
		x"11",	--1113
		x"5b",	--1114
		x"50",	--1115
		x"ff",	--1116
		x"4f",	--1117
		x"93",	--1118
		x"24",	--1119
		x"90",	--1120
		x"00",	--1121
		x"23",	--1122
		x"43",	--1123
		x"4f",	--1124
		x"93",	--1125
		x"23",	--1126
		x"12",	--1127
		x"c2",	--1128
		x"43",	--1129
		x"4a",	--1130
		x"01",	--1131
		x"4c",	--1132
		x"01",	--1133
		x"42",	--1134
		x"01",	--1135
		x"41",	--1136
		x"43",	--1137
		x"00",	--1138
		x"41",	--1139
		x"41",	--1140
		x"41",	--1141
		x"11",	--1142
		x"12",	--1143
		x"12",	--1144
		x"d5",	--1145
		x"12",	--1146
		x"9b",	--1147
		x"52",	--1148
		x"43",	--1149
		x"41",	--1150
		x"41",	--1151
		x"41",	--1152
		x"43",	--1153
		x"3f",	--1154
		x"12",	--1155
		x"12",	--1156
		x"12",	--1157
		x"4f",	--1158
		x"4f",	--1159
		x"00",	--1160
		x"12",	--1161
		x"99",	--1162
		x"4e",	--1163
		x"4f",	--1164
		x"89",	--1165
		x"00",	--1166
		x"79",	--1167
		x"00",	--1168
		x"12",	--1169
		x"c2",	--1170
		x"4a",	--1171
		x"00",	--1172
		x"4b",	--1173
		x"00",	--1174
		x"4e",	--1175
		x"4f",	--1176
		x"49",	--1177
		x"12",	--1178
		x"90",	--1179
		x"43",	--1180
		x"40",	--1181
		x"3f",	--1182
		x"12",	--1183
		x"bd",	--1184
		x"4e",	--1185
		x"4f",	--1186
		x"40",	--1187
		x"66",	--1188
		x"40",	--1189
		x"3f",	--1190
		x"12",	--1191
		x"c1",	--1192
		x"93",	--1193
		x"24",	--1194
		x"34",	--1195
		x"40",	--1196
		x"cc",	--1197
		x"40",	--1198
		x"3d",	--1199
		x"4a",	--1200
		x"4b",	--1201
		x"12",	--1202
		x"c2",	--1203
		x"93",	--1204
		x"34",	--1205
		x"40",	--1206
		x"cc",	--1207
		x"40",	--1208
		x"3d",	--1209
		x"4a",	--1210
		x"4b",	--1211
		x"49",	--1212
		x"00",	--1213
		x"12",	--1214
		x"96",	--1215
		x"41",	--1216
		x"41",	--1217
		x"41",	--1218
		x"41",	--1219
		x"40",	--1220
		x"66",	--1221
		x"40",	--1222
		x"3f",	--1223
		x"3f",	--1224
		x"12",	--1225
		x"12",	--1226
		x"4f",	--1227
		x"4c",	--1228
		x"4e",	--1229
		x"00",	--1230
		x"4d",	--1231
		x"00",	--1232
		x"12",	--1233
		x"00",	--1234
		x"12",	--1235
		x"00",	--1236
		x"12",	--1237
		x"00",	--1238
		x"12",	--1239
		x"00",	--1240
		x"12",	--1241
		x"00",	--1242
		x"12",	--1243
		x"00",	--1244
		x"41",	--1245
		x"00",	--1246
		x"41",	--1247
		x"00",	--1248
		x"12",	--1249
		x"8f",	--1250
		x"50",	--1251
		x"00",	--1252
		x"4a",	--1253
		x"00",	--1254
		x"4b",	--1255
		x"40",	--1256
		x"89",	--1257
		x"12",	--1258
		x"98",	--1259
		x"4f",	--1260
		x"00",	--1261
		x"41",	--1262
		x"41",	--1263
		x"41",	--1264
		x"12",	--1265
		x"4f",	--1266
		x"4f",	--1267
		x"00",	--1268
		x"12",	--1269
		x"99",	--1270
		x"4e",	--1271
		x"00",	--1272
		x"4f",	--1273
		x"00",	--1274
		x"43",	--1275
		x"4b",	--1276
		x"00",	--1277
		x"4b",	--1278
		x"00",	--1279
		x"12",	--1280
		x"98",	--1281
		x"41",	--1282
		x"41",	--1283
		x"12",	--1284
		x"4f",	--1285
		x"43",	--1286
		x"40",	--1287
		x"3f",	--1288
		x"4f",	--1289
		x"00",	--1290
		x"12",	--1291
		x"96",	--1292
		x"4b",	--1293
		x"00",	--1294
		x"12",	--1295
		x"98",	--1296
		x"41",	--1297
		x"41",	--1298
		x"12",	--1299
		x"4f",	--1300
		x"4e",	--1301
		x"10",	--1302
		x"11",	--1303
		x"10",	--1304
		x"11",	--1305
		x"4d",	--1306
		x"12",	--1307
		x"c2",	--1308
		x"4e",	--1309
		x"4f",	--1310
		x"4b",	--1311
		x"12",	--1312
		x"90",	--1313
		x"41",	--1314
		x"41",	--1315
		x"12",	--1316
		x"12",	--1317
		x"43",	--1318
		x"40",	--1319
		x"3f",	--1320
		x"4a",	--1321
		x"4b",	--1322
		x"42",	--1323
		x"02",	--1324
		x"12",	--1325
		x"96",	--1326
		x"4a",	--1327
		x"4b",	--1328
		x"42",	--1329
		x"02",	--1330
		x"12",	--1331
		x"96",	--1332
		x"12",	--1333
		x"d5",	--1334
		x"12",	--1335
		x"9b",	--1336
		x"53",	--1337
		x"41",	--1338
		x"41",	--1339
		x"41",	--1340
		x"4f",	--1341
		x"02",	--1342
		x"4e",	--1343
		x"02",	--1344
		x"41",	--1345
		x"12",	--1346
		x"12",	--1347
		x"83",	--1348
		x"4f",	--1349
		x"4e",	--1350
		x"93",	--1351
		x"02",	--1352
		x"24",	--1353
		x"90",	--1354
		x"00",	--1355
		x"38",	--1356
		x"20",	--1357
		x"41",	--1358
		x"4b",	--1359
		x"00",	--1360
		x"12",	--1361
		x"87",	--1362
		x"4f",	--1363
		x"41",	--1364
		x"4b",	--1365
		x"00",	--1366
		x"12",	--1367
		x"87",	--1368
		x"4f",	--1369
		x"12",	--1370
		x"12",	--1371
		x"12",	--1372
		x"d5",	--1373
		x"12",	--1374
		x"9b",	--1375
		x"50",	--1376
		x"00",	--1377
		x"4a",	--1378
		x"43",	--1379
		x"12",	--1380
		x"c3",	--1381
		x"43",	--1382
		x"40",	--1383
		x"42",	--1384
		x"12",	--1385
		x"bf",	--1386
		x"4e",	--1387
		x"4f",	--1388
		x"43",	--1389
		x"40",	--1390
		x"3f",	--1391
		x"12",	--1392
		x"bd",	--1393
		x"4e",	--1394
		x"4f",	--1395
		x"42",	--1396
		x"02",	--1397
		x"12",	--1398
		x"96",	--1399
		x"4b",	--1400
		x"43",	--1401
		x"12",	--1402
		x"c3",	--1403
		x"43",	--1404
		x"40",	--1405
		x"42",	--1406
		x"12",	--1407
		x"bf",	--1408
		x"4e",	--1409
		x"4f",	--1410
		x"42",	--1411
		x"02",	--1412
		x"12",	--1413
		x"96",	--1414
		x"43",	--1415
		x"53",	--1416
		x"41",	--1417
		x"41",	--1418
		x"41",	--1419
		x"41",	--1420
		x"4b",	--1421
		x"00",	--1422
		x"12",	--1423
		x"87",	--1424
		x"43",	--1425
		x"4f",	--1426
		x"42",	--1427
		x"02",	--1428
		x"12",	--1429
		x"98",	--1430
		x"3f",	--1431
		x"43",	--1432
		x"40",	--1433
		x"8a",	--1434
		x"12",	--1435
		x"98",	--1436
		x"4f",	--1437
		x"02",	--1438
		x"3f",	--1439
		x"12",	--1440
		x"d5",	--1441
		x"12",	--1442
		x"9b",	--1443
		x"40",	--1444
		x"d5",	--1445
		x"00",	--1446
		x"12",	--1447
		x"9b",	--1448
		x"4b",	--1449
		x"00",	--1450
		x"12",	--1451
		x"d5",	--1452
		x"12",	--1453
		x"9b",	--1454
		x"52",	--1455
		x"43",	--1456
		x"3f",	--1457
		x"12",	--1458
		x"12",	--1459
		x"42",	--1460
		x"02",	--1461
		x"12",	--1462
		x"99",	--1463
		x"4e",	--1464
		x"4f",	--1465
		x"42",	--1466
		x"02",	--1467
		x"12",	--1468
		x"99",	--1469
		x"12",	--1470
		x"12",	--1471
		x"e3",	--1472
		x"e3",	--1473
		x"53",	--1474
		x"63",	--1475
		x"12",	--1476
		x"12",	--1477
		x"12",	--1478
		x"d5",	--1479
		x"12",	--1480
		x"02",	--1481
		x"12",	--1482
		x"c9",	--1483
		x"50",	--1484
		x"00",	--1485
		x"12",	--1486
		x"02",	--1487
		x"12",	--1488
		x"d5",	--1489
		x"12",	--1490
		x"9b",	--1491
		x"52",	--1492
		x"41",	--1493
		x"41",	--1494
		x"41",	--1495
		x"4f",	--1496
		x"02",	--1497
		x"4e",	--1498
		x"02",	--1499
		x"41",	--1500
		x"4f",	--1501
		x"02",	--1502
		x"4e",	--1503
		x"02",	--1504
		x"41",	--1505
		x"12",	--1506
		x"12",	--1507
		x"12",	--1508
		x"12",	--1509
		x"83",	--1510
		x"4f",	--1511
		x"4e",	--1512
		x"43",	--1513
		x"00",	--1514
		x"93",	--1515
		x"24",	--1516
		x"93",	--1517
		x"02",	--1518
		x"24",	--1519
		x"43",	--1520
		x"02",	--1521
		x"41",	--1522
		x"4b",	--1523
		x"00",	--1524
		x"12",	--1525
		x"87",	--1526
		x"4f",	--1527
		x"90",	--1528
		x"00",	--1529
		x"34",	--1530
		x"43",	--1531
		x"49",	--1532
		x"48",	--1533
		x"42",	--1534
		x"02",	--1535
		x"12",	--1536
		x"98",	--1537
		x"43",	--1538
		x"53",	--1539
		x"41",	--1540
		x"41",	--1541
		x"41",	--1542
		x"41",	--1543
		x"41",	--1544
		x"93",	--1545
		x"02",	--1546
		x"24",	--1547
		x"43",	--1548
		x"02",	--1549
		x"42",	--1550
		x"02",	--1551
		x"12",	--1552
		x"98",	--1553
		x"43",	--1554
		x"53",	--1555
		x"41",	--1556
		x"41",	--1557
		x"41",	--1558
		x"41",	--1559
		x"41",	--1560
		x"41",	--1561
		x"4b",	--1562
		x"00",	--1563
		x"12",	--1564
		x"87",	--1565
		x"4f",	--1566
		x"90",	--1567
		x"00",	--1568
		x"3b",	--1569
		x"41",	--1570
		x"4b",	--1571
		x"00",	--1572
		x"12",	--1573
		x"87",	--1574
		x"4f",	--1575
		x"41",	--1576
		x"4b",	--1577
		x"00",	--1578
		x"12",	--1579
		x"87",	--1580
		x"4f",	--1581
		x"12",	--1582
		x"12",	--1583
		x"12",	--1584
		x"d5",	--1585
		x"12",	--1586
		x"9b",	--1587
		x"50",	--1588
		x"00",	--1589
		x"4a",	--1590
		x"43",	--1591
		x"12",	--1592
		x"c3",	--1593
		x"43",	--1594
		x"40",	--1595
		x"42",	--1596
		x"12",	--1597
		x"bf",	--1598
		x"4e",	--1599
		x"4f",	--1600
		x"42",	--1601
		x"02",	--1602
		x"12",	--1603
		x"96",	--1604
		x"4b",	--1605
		x"43",	--1606
		x"12",	--1607
		x"c3",	--1608
		x"43",	--1609
		x"40",	--1610
		x"42",	--1611
		x"12",	--1612
		x"bf",	--1613
		x"4e",	--1614
		x"4f",	--1615
		x"42",	--1616
		x"02",	--1617
		x"12",	--1618
		x"96",	--1619
		x"3f",	--1620
		x"43",	--1621
		x"12",	--1622
		x"8b",	--1623
		x"43",	--1624
		x"53",	--1625
		x"41",	--1626
		x"41",	--1627
		x"41",	--1628
		x"41",	--1629
		x"41",	--1630
		x"43",	--1631
		x"40",	--1632
		x"8b",	--1633
		x"12",	--1634
		x"98",	--1635
		x"4f",	--1636
		x"02",	--1637
		x"3f",	--1638
		x"12",	--1639
		x"12",	--1640
		x"12",	--1641
		x"12",	--1642
		x"4f",	--1643
		x"40",	--1644
		x"02",	--1645
		x"43",	--1646
		x"43",	--1647
		x"4b",	--1648
		x"48",	--1649
		x"12",	--1650
		x"98",	--1651
		x"9a",	--1652
		x"2c",	--1653
		x"43",	--1654
		x"4b",	--1655
		x"f0",	--1656
		x"00",	--1657
		x"24",	--1658
		x"5e",	--1659
		x"53",	--1660
		x"23",	--1661
		x"5e",	--1662
		x"53",	--1663
		x"53",	--1664
		x"90",	--1665
		x"00",	--1666
		x"23",	--1667
		x"49",	--1668
		x"41",	--1669
		x"41",	--1670
		x"41",	--1671
		x"41",	--1672
		x"41",	--1673
		x"12",	--1674
		x"12",	--1675
		x"93",	--1676
		x"02",	--1677
		x"20",	--1678
		x"41",	--1679
		x"41",	--1680
		x"41",	--1681
		x"42",	--1682
		x"02",	--1683
		x"12",	--1684
		x"8c",	--1685
		x"4f",	--1686
		x"43",	--1687
		x"4b",	--1688
		x"42",	--1689
		x"02",	--1690
		x"12",	--1691
		x"98",	--1692
		x"12",	--1693
		x"12",	--1694
		x"d5",	--1695
		x"12",	--1696
		x"9b",	--1697
		x"52",	--1698
		x"53",	--1699
		x"90",	--1700
		x"00",	--1701
		x"23",	--1702
		x"12",	--1703
		x"d5",	--1704
		x"12",	--1705
		x"9b",	--1706
		x"53",	--1707
		x"42",	--1708
		x"02",	--1709
		x"93",	--1710
		x"20",	--1711
		x"93",	--1712
		x"24",	--1713
		x"b0",	--1714
		x"00",	--1715
		x"20",	--1716
		x"b3",	--1717
		x"20",	--1718
		x"b3",	--1719
		x"20",	--1720
		x"b2",	--1721
		x"24",	--1722
		x"43",	--1723
		x"02",	--1724
		x"43",	--1725
		x"42",	--1726
		x"02",	--1727
		x"12",	--1728
		x"8a",	--1729
		x"43",	--1730
		x"42",	--1731
		x"02",	--1732
		x"12",	--1733
		x"8a",	--1734
		x"40",	--1735
		x"00",	--1736
		x"02",	--1737
		x"40",	--1738
		x"00",	--1739
		x"02",	--1740
		x"12",	--1741
		x"d6",	--1742
		x"12",	--1743
		x"9b",	--1744
		x"53",	--1745
		x"3f",	--1746
		x"93",	--1747
		x"02",	--1748
		x"20",	--1749
		x"42",	--1750
		x"02",	--1751
		x"93",	--1752
		x"24",	--1753
		x"93",	--1754
		x"24",	--1755
		x"93",	--1756
		x"24",	--1757
		x"90",	--1758
		x"00",	--1759
		x"24",	--1760
		x"53",	--1761
		x"4e",	--1762
		x"02",	--1763
		x"3f",	--1764
		x"43",	--1765
		x"02",	--1766
		x"3f",	--1767
		x"43",	--1768
		x"42",	--1769
		x"02",	--1770
		x"12",	--1771
		x"8a",	--1772
		x"43",	--1773
		x"42",	--1774
		x"02",	--1775
		x"12",	--1776
		x"8a",	--1777
		x"12",	--1778
		x"d6",	--1779
		x"12",	--1780
		x"9b",	--1781
		x"53",	--1782
		x"53",	--1783
		x"02",	--1784
		x"93",	--1785
		x"23",	--1786
		x"43",	--1787
		x"02",	--1788
		x"43",	--1789
		x"02",	--1790
		x"43",	--1791
		x"02",	--1792
		x"3f",	--1793
		x"43",	--1794
		x"42",	--1795
		x"02",	--1796
		x"12",	--1797
		x"8a",	--1798
		x"43",	--1799
		x"42",	--1800
		x"02",	--1801
		x"12",	--1802
		x"8a",	--1803
		x"12",	--1804
		x"12",	--1805
		x"d6",	--1806
		x"12",	--1807
		x"9b",	--1808
		x"52",	--1809
		x"3f",	--1810
		x"40",	--1811
		x"00",	--1812
		x"42",	--1813
		x"02",	--1814
		x"12",	--1815
		x"8a",	--1816
		x"40",	--1817
		x"00",	--1818
		x"42",	--1819
		x"02",	--1820
		x"12",	--1821
		x"8a",	--1822
		x"12",	--1823
		x"d6",	--1824
		x"12",	--1825
		x"9b",	--1826
		x"53",	--1827
		x"42",	--1828
		x"02",	--1829
		x"3f",	--1830
		x"40",	--1831
		x"00",	--1832
		x"42",	--1833
		x"02",	--1834
		x"12",	--1835
		x"8a",	--1836
		x"40",	--1837
		x"ff",	--1838
		x"42",	--1839
		x"02",	--1840
		x"12",	--1841
		x"8a",	--1842
		x"3f",	--1843
		x"12",	--1844
		x"d5",	--1845
		x"12",	--1846
		x"9b",	--1847
		x"53",	--1848
		x"3f",	--1849
		x"43",	--1850
		x"02",	--1851
		x"43",	--1852
		x"42",	--1853
		x"02",	--1854
		x"12",	--1855
		x"8a",	--1856
		x"43",	--1857
		x"42",	--1858
		x"02",	--1859
		x"12",	--1860
		x"8a",	--1861
		x"40",	--1862
		x"00",	--1863
		x"02",	--1864
		x"40",	--1865
		x"00",	--1866
		x"02",	--1867
		x"12",	--1868
		x"d5",	--1869
		x"12",	--1870
		x"9b",	--1871
		x"53",	--1872
		x"3f",	--1873
		x"40",	--1874
		x"00",	--1875
		x"02",	--1876
		x"43",	--1877
		x"42",	--1878
		x"02",	--1879
		x"12",	--1880
		x"8a",	--1881
		x"43",	--1882
		x"42",	--1883
		x"02",	--1884
		x"12",	--1885
		x"8a",	--1886
		x"40",	--1887
		x"00",	--1888
		x"02",	--1889
		x"40",	--1890
		x"00",	--1891
		x"02",	--1892
		x"12",	--1893
		x"d5",	--1894
		x"12",	--1895
		x"9b",	--1896
		x"53",	--1897
		x"3f",	--1898
		x"40",	--1899
		x"00",	--1900
		x"42",	--1901
		x"02",	--1902
		x"12",	--1903
		x"8a",	--1904
		x"40",	--1905
		x"00",	--1906
		x"42",	--1907
		x"02",	--1908
		x"12",	--1909
		x"8a",	--1910
		x"12",	--1911
		x"d6",	--1912
		x"12",	--1913
		x"9b",	--1914
		x"53",	--1915
		x"42",	--1916
		x"02",	--1917
		x"3f",	--1918
		x"40",	--1919
		x"ff",	--1920
		x"42",	--1921
		x"02",	--1922
		x"12",	--1923
		x"8a",	--1924
		x"40",	--1925
		x"ff",	--1926
		x"42",	--1927
		x"02",	--1928
		x"12",	--1929
		x"8a",	--1930
		x"12",	--1931
		x"d6",	--1932
		x"12",	--1933
		x"9b",	--1934
		x"53",	--1935
		x"42",	--1936
		x"02",	--1937
		x"3f",	--1938
		x"4f",	--1939
		x"02",	--1940
		x"4e",	--1941
		x"02",	--1942
		x"41",	--1943
		x"4f",	--1944
		x"02",	--1945
		x"41",	--1946
		x"12",	--1947
		x"4f",	--1948
		x"43",	--1949
		x"40",	--1950
		x"8d",	--1951
		x"12",	--1952
		x"98",	--1953
		x"4f",	--1954
		x"02",	--1955
		x"43",	--1956
		x"4b",	--1957
		x"12",	--1958
		x"98",	--1959
		x"41",	--1960
		x"41",	--1961
		x"43",	--1962
		x"93",	--1963
		x"02",	--1964
		x"24",	--1965
		x"43",	--1966
		x"4f",	--1967
		x"02",	--1968
		x"93",	--1969
		x"20",	--1970
		x"43",	--1971
		x"42",	--1972
		x"02",	--1973
		x"12",	--1974
		x"8a",	--1975
		x"43",	--1976
		x"42",	--1977
		x"02",	--1978
		x"12",	--1979
		x"8a",	--1980
		x"12",	--1981
		x"d6",	--1982
		x"12",	--1983
		x"9b",	--1984
		x"53",	--1985
		x"43",	--1986
		x"41",	--1987
		x"12",	--1988
		x"d6",	--1989
		x"12",	--1990
		x"9b",	--1991
		x"53",	--1992
		x"43",	--1993
		x"41",	--1994
		x"4d",	--1995
		x"00",	--1996
		x"4e",	--1997
		x"00",	--1998
		x"41",	--1999
		x"00",	--2000
		x"00",	--2001
		x"41",	--2002
		x"00",	--2003
		x"00",	--2004
		x"41",	--2005
		x"00",	--2006
		x"00",	--2007
		x"41",	--2008
		x"00",	--2009
		x"00",	--2010
		x"41",	--2011
		x"00",	--2012
		x"00",	--2013
		x"41",	--2014
		x"00",	--2015
		x"00",	--2016
		x"43",	--2017
		x"00",	--2018
		x"43",	--2019
		x"00",	--2020
		x"43",	--2021
		x"00",	--2022
		x"43",	--2023
		x"00",	--2024
		x"43",	--2025
		x"00",	--2026
		x"43",	--2027
		x"00",	--2028
		x"43",	--2029
		x"00",	--2030
		x"43",	--2031
		x"00",	--2032
		x"41",	--2033
		x"43",	--2034
		x"00",	--2035
		x"43",	--2036
		x"00",	--2037
		x"43",	--2038
		x"00",	--2039
		x"43",	--2040
		x"00",	--2041
		x"43",	--2042
		x"00",	--2043
		x"43",	--2044
		x"00",	--2045
		x"41",	--2046
		x"4d",	--2047
		x"00",	--2048
		x"4e",	--2049
		x"00",	--2050
		x"41",	--2051
		x"4d",	--2052
		x"00",	--2053
		x"4e",	--2054
		x"00",	--2055
		x"41",	--2056
		x"4d",	--2057
		x"00",	--2058
		x"4e",	--2059
		x"00",	--2060
		x"41",	--2061
		x"4d",	--2062
		x"00",	--2063
		x"4e",	--2064
		x"00",	--2065
		x"41",	--2066
		x"4d",	--2067
		x"00",	--2068
		x"4e",	--2069
		x"00",	--2070
		x"41",	--2071
		x"12",	--2072
		x"12",	--2073
		x"12",	--2074
		x"12",	--2075
		x"12",	--2076
		x"12",	--2077
		x"12",	--2078
		x"4f",	--2079
		x"4d",	--2080
		x"4e",	--2081
		x"4f",	--2082
		x"00",	--2083
		x"4f",	--2084
		x"00",	--2085
		x"4f",	--2086
		x"00",	--2087
		x"4f",	--2088
		x"00",	--2089
		x"4a",	--2090
		x"4b",	--2091
		x"46",	--2092
		x"47",	--2093
		x"12",	--2094
		x"c2",	--2095
		x"49",	--2096
		x"00",	--2097
		x"49",	--2098
		x"00",	--2099
		x"93",	--2100
		x"34",	--2101
		x"46",	--2102
		x"47",	--2103
		x"12",	--2104
		x"bd",	--2105
		x"4e",	--2106
		x"4f",	--2107
		x"4e",	--2108
		x"00",	--2109
		x"4f",	--2110
		x"00",	--2111
		x"4e",	--2112
		x"4f",	--2113
		x"4a",	--2114
		x"4b",	--2115
		x"12",	--2116
		x"c2",	--2117
		x"93",	--2118
		x"34",	--2119
		x"4a",	--2120
		x"00",	--2121
		x"4b",	--2122
		x"00",	--2123
		x"44",	--2124
		x"45",	--2125
		x"4a",	--2126
		x"4b",	--2127
		x"12",	--2128
		x"bd",	--2129
		x"4e",	--2130
		x"4f",	--2131
		x"49",	--2132
		x"00",	--2133
		x"49",	--2134
		x"00",	--2135
		x"12",	--2136
		x"bd",	--2137
		x"4e",	--2138
		x"4f",	--2139
		x"4e",	--2140
		x"00",	--2141
		x"4f",	--2142
		x"00",	--2143
		x"49",	--2144
		x"49",	--2145
		x"00",	--2146
		x"4a",	--2147
		x"4b",	--2148
		x"12",	--2149
		x"bd",	--2150
		x"4e",	--2151
		x"4f",	--2152
		x"49",	--2153
		x"00",	--2154
		x"49",	--2155
		x"00",	--2156
		x"46",	--2157
		x"47",	--2158
		x"12",	--2159
		x"bd",	--2160
		x"44",	--2161
		x"45",	--2162
		x"12",	--2163
		x"bd",	--2164
		x"4e",	--2165
		x"4f",	--2166
		x"49",	--2167
		x"00",	--2168
		x"49",	--2169
		x"00",	--2170
		x"4a",	--2171
		x"4b",	--2172
		x"12",	--2173
		x"bd",	--2174
		x"49",	--2175
		x"00",	--2176
		x"49",	--2177
		x"00",	--2178
		x"12",	--2179
		x"bd",	--2180
		x"46",	--2181
		x"47",	--2182
		x"12",	--2183
		x"bd",	--2184
		x"41",	--2185
		x"41",	--2186
		x"41",	--2187
		x"41",	--2188
		x"41",	--2189
		x"41",	--2190
		x"41",	--2191
		x"41",	--2192
		x"46",	--2193
		x"47",	--2194
		x"12",	--2195
		x"bd",	--2196
		x"4e",	--2197
		x"4f",	--2198
		x"4e",	--2199
		x"00",	--2200
		x"4f",	--2201
		x"00",	--2202
		x"4e",	--2203
		x"4f",	--2204
		x"4a",	--2205
		x"4b",	--2206
		x"12",	--2207
		x"c1",	--2208
		x"93",	--2209
		x"24",	--2210
		x"37",	--2211
		x"46",	--2212
		x"47",	--2213
		x"3f",	--2214
		x"12",	--2215
		x"12",	--2216
		x"83",	--2217
		x"4f",	--2218
		x"4e",	--2219
		x"12",	--2220
		x"d6",	--2221
		x"12",	--2222
		x"9b",	--2223
		x"53",	--2224
		x"90",	--2225
		x"00",	--2226
		x"38",	--2227
		x"41",	--2228
		x"4b",	--2229
		x"00",	--2230
		x"12",	--2231
		x"87",	--2232
		x"4f",	--2233
		x"41",	--2234
		x"4b",	--2235
		x"00",	--2236
		x"12",	--2237
		x"87",	--2238
		x"4f",	--2239
		x"12",	--2240
		x"12",	--2241
		x"12",	--2242
		x"d6",	--2243
		x"12",	--2244
		x"9b",	--2245
		x"50",	--2246
		x"00",	--2247
		x"4b",	--2248
		x"00",	--2249
		x"43",	--2250
		x"53",	--2251
		x"41",	--2252
		x"41",	--2253
		x"41",	--2254
		x"12",	--2255
		x"d6",	--2256
		x"12",	--2257
		x"9b",	--2258
		x"40",	--2259
		x"d6",	--2260
		x"00",	--2261
		x"12",	--2262
		x"9b",	--2263
		x"4b",	--2264
		x"00",	--2265
		x"12",	--2266
		x"d6",	--2267
		x"12",	--2268
		x"9b",	--2269
		x"52",	--2270
		x"43",	--2271
		x"3f",	--2272
		x"12",	--2273
		x"83",	--2274
		x"4e",	--2275
		x"93",	--2276
		x"24",	--2277
		x"38",	--2278
		x"12",	--2279
		x"d6",	--2280
		x"12",	--2281
		x"9b",	--2282
		x"53",	--2283
		x"41",	--2284
		x"4b",	--2285
		x"00",	--2286
		x"12",	--2287
		x"87",	--2288
		x"12",	--2289
		x"12",	--2290
		x"12",	--2291
		x"d6",	--2292
		x"12",	--2293
		x"9b",	--2294
		x"50",	--2295
		x"00",	--2296
		x"43",	--2297
		x"53",	--2298
		x"41",	--2299
		x"41",	--2300
		x"12",	--2301
		x"d6",	--2302
		x"12",	--2303
		x"9b",	--2304
		x"40",	--2305
		x"d6",	--2306
		x"00",	--2307
		x"12",	--2308
		x"9b",	--2309
		x"4b",	--2310
		x"00",	--2311
		x"12",	--2312
		x"d6",	--2313
		x"12",	--2314
		x"9b",	--2315
		x"52",	--2316
		x"43",	--2317
		x"3f",	--2318
		x"12",	--2319
		x"12",	--2320
		x"12",	--2321
		x"12",	--2322
		x"12",	--2323
		x"12",	--2324
		x"4e",	--2325
		x"4f",	--2326
		x"4c",	--2327
		x"4d",	--2328
		x"12",	--2329
		x"bd",	--2330
		x"4e",	--2331
		x"4f",	--2332
		x"40",	--2333
		x"0f",	--2334
		x"40",	--2335
		x"c0",	--2336
		x"12",	--2337
		x"c2",	--2338
		x"93",	--2339
		x"24",	--2340
		x"38",	--2341
		x"40",	--2342
		x"0f",	--2343
		x"40",	--2344
		x"40",	--2345
		x"4a",	--2346
		x"4b",	--2347
		x"12",	--2348
		x"c1",	--2349
		x"93",	--2350
		x"24",	--2351
		x"34",	--2352
		x"4a",	--2353
		x"4b",	--2354
		x"41",	--2355
		x"41",	--2356
		x"41",	--2357
		x"41",	--2358
		x"41",	--2359
		x"41",	--2360
		x"41",	--2361
		x"40",	--2362
		x"0f",	--2363
		x"40",	--2364
		x"40",	--2365
		x"4a",	--2366
		x"4b",	--2367
		x"12",	--2368
		x"bd",	--2369
		x"4e",	--2370
		x"4f",	--2371
		x"3f",	--2372
		x"40",	--2373
		x"0f",	--2374
		x"40",	--2375
		x"40",	--2376
		x"46",	--2377
		x"47",	--2378
		x"12",	--2379
		x"bd",	--2380
		x"48",	--2381
		x"49",	--2382
		x"12",	--2383
		x"bd",	--2384
		x"4e",	--2385
		x"4f",	--2386
		x"3f",	--2387
		x"12",	--2388
		x"4f",	--2389
		x"43",	--2390
		x"00",	--2391
		x"43",	--2392
		x"00",	--2393
		x"43",	--2394
		x"00",	--2395
		x"43",	--2396
		x"00",	--2397
		x"43",	--2398
		x"00",	--2399
		x"43",	--2400
		x"00",	--2401
		x"4d",	--2402
		x"00",	--2403
		x"4e",	--2404
		x"00",	--2405
		x"41",	--2406
		x"00",	--2407
		x"00",	--2408
		x"41",	--2409
		x"00",	--2410
		x"00",	--2411
		x"41",	--2412
		x"00",	--2413
		x"00",	--2414
		x"43",	--2415
		x"00",	--2416
		x"43",	--2417
		x"00",	--2418
		x"43",	--2419
		x"00",	--2420
		x"43",	--2421
		x"00",	--2422
		x"4f",	--2423
		x"40",	--2424
		x"95",	--2425
		x"12",	--2426
		x"98",	--2427
		x"4f",	--2428
		x"00",	--2429
		x"41",	--2430
		x"41",	--2431
		x"4e",	--2432
		x"00",	--2433
		x"4d",	--2434
		x"00",	--2435
		x"41",	--2436
		x"12",	--2437
		x"12",	--2438
		x"12",	--2439
		x"12",	--2440
		x"12",	--2441
		x"12",	--2442
		x"12",	--2443
		x"50",	--2444
		x"ff",	--2445
		x"4f",	--2446
		x"4d",	--2447
		x"00",	--2448
		x"4e",	--2449
		x"00",	--2450
		x"40",	--2451
		x"0f",	--2452
		x"40",	--2453
		x"40",	--2454
		x"4f",	--2455
		x"4f",	--2456
		x"00",	--2457
		x"12",	--2458
		x"bd",	--2459
		x"4e",	--2460
		x"4f",	--2461
		x"47",	--2462
		x"00",	--2463
		x"4e",	--2464
		x"10",	--2465
		x"11",	--2466
		x"10",	--2467
		x"11",	--2468
		x"12",	--2469
		x"c2",	--2470
		x"4e",	--2471
		x"4f",	--2472
		x"4a",	--2473
		x"4b",	--2474
		x"12",	--2475
		x"bf",	--2476
		x"4e",	--2477
		x"4f",	--2478
		x"41",	--2479
		x"00",	--2480
		x"41",	--2481
		x"00",	--2482
		x"87",	--2483
		x"00",	--2484
		x"77",	--2485
		x"00",	--2486
		x"41",	--2487
		x"00",	--2488
		x"41",	--2489
		x"00",	--2490
		x"87",	--2491
		x"00",	--2492
		x"77",	--2493
		x"00",	--2494
		x"48",	--2495
		x"49",	--2496
		x"12",	--2497
		x"c2",	--2498
		x"4a",	--2499
		x"4b",	--2500
		x"12",	--2501
		x"bd",	--2502
		x"4e",	--2503
		x"00",	--2504
		x"4f",	--2505
		x"00",	--2506
		x"44",	--2507
		x"45",	--2508
		x"12",	--2509
		x"c2",	--2510
		x"4a",	--2511
		x"4b",	--2512
		x"12",	--2513
		x"bd",	--2514
		x"4e",	--2515
		x"4f",	--2516
		x"4e",	--2517
		x"4f",	--2518
		x"41",	--2519
		x"41",	--2520
		x"00",	--2521
		x"12",	--2522
		x"bd",	--2523
		x"4e",	--2524
		x"00",	--2525
		x"4f",	--2526
		x"00",	--2527
		x"93",	--2528
		x"20",	--2529
		x"93",	--2530
		x"20",	--2531
		x"93",	--2532
		x"20",	--2533
		x"40",	--2534
		x"95",	--2535
		x"47",	--2536
		x"00",	--2537
		x"47",	--2538
		x"00",	--2539
		x"41",	--2540
		x"41",	--2541
		x"00",	--2542
		x"4a",	--2543
		x"4b",	--2544
		x"12",	--2545
		x"bd",	--2546
		x"4e",	--2547
		x"4f",	--2548
		x"48",	--2549
		x"49",	--2550
		x"41",	--2551
		x"00",	--2552
		x"41",	--2553
		x"00",	--2554
		x"12",	--2555
		x"bd",	--2556
		x"4a",	--2557
		x"4b",	--2558
		x"12",	--2559
		x"bf",	--2560
		x"4e",	--2561
		x"4f",	--2562
		x"48",	--2563
		x"49",	--2564
		x"48",	--2565
		x"49",	--2566
		x"12",	--2567
		x"bd",	--2568
		x"4e",	--2569
		x"4f",	--2570
		x"4a",	--2571
		x"4b",	--2572
		x"12",	--2573
		x"bf",	--2574
		x"12",	--2575
		x"a0",	--2576
		x"4e",	--2577
		x"00",	--2578
		x"4f",	--2579
		x"00",	--2580
		x"47",	--2581
		x"00",	--2582
		x"47",	--2583
		x"00",	--2584
		x"4a",	--2585
		x"4b",	--2586
		x"12",	--2587
		x"a1",	--2588
		x"44",	--2589
		x"45",	--2590
		x"12",	--2591
		x"bd",	--2592
		x"4e",	--2593
		x"4f",	--2594
		x"47",	--2595
		x"00",	--2596
		x"47",	--2597
		x"00",	--2598
		x"12",	--2599
		x"bd",	--2600
		x"4e",	--2601
		x"00",	--2602
		x"4f",	--2603
		x"00",	--2604
		x"4a",	--2605
		x"4b",	--2606
		x"12",	--2607
		x"b6",	--2608
		x"44",	--2609
		x"45",	--2610
		x"12",	--2611
		x"bd",	--2612
		x"47",	--2613
		x"00",	--2614
		x"47",	--2615
		x"00",	--2616
		x"12",	--2617
		x"bd",	--2618
		x"4e",	--2619
		x"4f",	--2620
		x"41",	--2621
		x"41",	--2622
		x"00",	--2623
		x"4a",	--2624
		x"4b",	--2625
		x"12",	--2626
		x"92",	--2627
		x"4e",	--2628
		x"4f",	--2629
		x"4e",	--2630
		x"00",	--2631
		x"4f",	--2632
		x"00",	--2633
		x"12",	--2634
		x"a1",	--2635
		x"44",	--2636
		x"45",	--2637
		x"12",	--2638
		x"bd",	--2639
		x"41",	--2640
		x"00",	--2641
		x"41",	--2642
		x"00",	--2643
		x"12",	--2644
		x"bd",	--2645
		x"4e",	--2646
		x"00",	--2647
		x"4f",	--2648
		x"00",	--2649
		x"4a",	--2650
		x"4b",	--2651
		x"12",	--2652
		x"b6",	--2653
		x"44",	--2654
		x"45",	--2655
		x"12",	--2656
		x"bd",	--2657
		x"4e",	--2658
		x"4f",	--2659
		x"48",	--2660
		x"49",	--2661
		x"12",	--2662
		x"bd",	--2663
		x"4e",	--2664
		x"00",	--2665
		x"4f",	--2666
		x"00",	--2667
		x"41",	--2668
		x"00",	--2669
		x"00",	--2670
		x"41",	--2671
		x"00",	--2672
		x"00",	--2673
		x"41",	--2674
		x"00",	--2675
		x"00",	--2676
		x"41",	--2677
		x"00",	--2678
		x"00",	--2679
		x"50",	--2680
		x"00",	--2681
		x"41",	--2682
		x"41",	--2683
		x"41",	--2684
		x"41",	--2685
		x"41",	--2686
		x"41",	--2687
		x"41",	--2688
		x"41",	--2689
		x"94",	--2690
		x"23",	--2691
		x"95",	--2692
		x"23",	--2693
		x"43",	--2694
		x"40",	--2695
		x"3f",	--2696
		x"41",	--2697
		x"00",	--2698
		x"41",	--2699
		x"00",	--2700
		x"12",	--2701
		x"bd",	--2702
		x"4e",	--2703
		x"4f",	--2704
		x"47",	--2705
		x"00",	--2706
		x"47",	--2707
		x"00",	--2708
		x"48",	--2709
		x"49",	--2710
		x"12",	--2711
		x"b6",	--2712
		x"4a",	--2713
		x"4b",	--2714
		x"12",	--2715
		x"bd",	--2716
		x"4e",	--2717
		x"4f",	--2718
		x"47",	--2719
		x"00",	--2720
		x"47",	--2721
		x"00",	--2722
		x"12",	--2723
		x"bd",	--2724
		x"4e",	--2725
		x"00",	--2726
		x"4f",	--2727
		x"00",	--2728
		x"48",	--2729
		x"49",	--2730
		x"12",	--2731
		x"a1",	--2732
		x"4a",	--2733
		x"4b",	--2734
		x"12",	--2735
		x"bd",	--2736
		x"4e",	--2737
		x"4f",	--2738
		x"47",	--2739
		x"00",	--2740
		x"47",	--2741
		x"00",	--2742
		x"12",	--2743
		x"bd",	--2744
		x"4e",	--2745
		x"00",	--2746
		x"4f",	--2747
		x"00",	--2748
		x"3f",	--2749
		x"93",	--2750
		x"27",	--2751
		x"40",	--2752
		x"93",	--2753
		x"12",	--2754
		x"12",	--2755
		x"12",	--2756
		x"4f",	--2757
		x"4f",	--2758
		x"00",	--2759
		x"12",	--2760
		x"99",	--2761
		x"4e",	--2762
		x"4f",	--2763
		x"49",	--2764
		x"00",	--2765
		x"12",	--2766
		x"99",	--2767
		x"4a",	--2768
		x"4b",	--2769
		x"e3",	--2770
		x"e3",	--2771
		x"53",	--2772
		x"63",	--2773
		x"12",	--2774
		x"12",	--2775
		x"4e",	--2776
		x"4f",	--2777
		x"49",	--2778
		x"12",	--2779
		x"93",	--2780
		x"52",	--2781
		x"41",	--2782
		x"41",	--2783
		x"41",	--2784
		x"41",	--2785
		x"43",	--2786
		x"4f",	--2787
		x"00",	--2788
		x"12",	--2789
		x"98",	--2790
		x"41",	--2791
		x"4f",	--2792
		x"00",	--2793
		x"12",	--2794
		x"98",	--2795
		x"41",	--2796
		x"12",	--2797
		x"12",	--2798
		x"4e",	--2799
		x"4c",	--2800
		x"4e",	--2801
		x"00",	--2802
		x"4d",	--2803
		x"00",	--2804
		x"4c",	--2805
		x"00",	--2806
		x"4d",	--2807
		x"43",	--2808
		x"40",	--2809
		x"36",	--2810
		x"40",	--2811
		x"01",	--2812
		x"12",	--2813
		x"d2",	--2814
		x"4e",	--2815
		x"00",	--2816
		x"12",	--2817
		x"c2",	--2818
		x"43",	--2819
		x"4a",	--2820
		x"01",	--2821
		x"40",	--2822
		x"00",	--2823
		x"01",	--2824
		x"42",	--2825
		x"01",	--2826
		x"00",	--2827
		x"41",	--2828
		x"43",	--2829
		x"41",	--2830
		x"41",	--2831
		x"41",	--2832
		x"12",	--2833
		x"12",	--2834
		x"12",	--2835
		x"43",	--2836
		x"00",	--2837
		x"40",	--2838
		x"3f",	--2839
		x"00",	--2840
		x"4f",	--2841
		x"4b",	--2842
		x"00",	--2843
		x"43",	--2844
		x"12",	--2845
		x"c3",	--2846
		x"43",	--2847
		x"40",	--2848
		x"3f",	--2849
		x"12",	--2850
		x"bd",	--2851
		x"4e",	--2852
		x"4f",	--2853
		x"4b",	--2854
		x"00",	--2855
		x"43",	--2856
		x"12",	--2857
		x"c3",	--2858
		x"4e",	--2859
		x"4f",	--2860
		x"48",	--2861
		x"49",	--2862
		x"12",	--2863
		x"bd",	--2864
		x"12",	--2865
		x"ba",	--2866
		x"4e",	--2867
		x"00",	--2868
		x"43",	--2869
		x"00",	--2870
		x"41",	--2871
		x"41",	--2872
		x"41",	--2873
		x"41",	--2874
		x"12",	--2875
		x"12",	--2876
		x"12",	--2877
		x"4d",	--2878
		x"4e",	--2879
		x"4d",	--2880
		x"00",	--2881
		x"4e",	--2882
		x"00",	--2883
		x"4f",	--2884
		x"49",	--2885
		x"00",	--2886
		x"43",	--2887
		x"12",	--2888
		x"c3",	--2889
		x"4e",	--2890
		x"4f",	--2891
		x"4a",	--2892
		x"4b",	--2893
		x"12",	--2894
		x"bd",	--2895
		x"4e",	--2896
		x"4f",	--2897
		x"49",	--2898
		x"00",	--2899
		x"43",	--2900
		x"12",	--2901
		x"c3",	--2902
		x"4e",	--2903
		x"4f",	--2904
		x"4a",	--2905
		x"4b",	--2906
		x"12",	--2907
		x"bd",	--2908
		x"12",	--2909
		x"ba",	--2910
		x"4e",	--2911
		x"00",	--2912
		x"41",	--2913
		x"41",	--2914
		x"41",	--2915
		x"41",	--2916
		x"4f",	--2917
		x"4e",	--2918
		x"00",	--2919
		x"41",	--2920
		x"12",	--2921
		x"12",	--2922
		x"93",	--2923
		x"02",	--2924
		x"38",	--2925
		x"40",	--2926
		x"02",	--2927
		x"43",	--2928
		x"12",	--2929
		x"4b",	--2930
		x"ff",	--2931
		x"11",	--2932
		x"12",	--2933
		x"12",	--2934
		x"d6",	--2935
		x"12",	--2936
		x"9b",	--2937
		x"50",	--2938
		x"00",	--2939
		x"53",	--2940
		x"50",	--2941
		x"00",	--2942
		x"92",	--2943
		x"02",	--2944
		x"3b",	--2945
		x"43",	--2946
		x"41",	--2947
		x"41",	--2948
		x"41",	--2949
		x"42",	--2950
		x"02",	--2951
		x"90",	--2952
		x"00",	--2953
		x"34",	--2954
		x"4e",	--2955
		x"5f",	--2956
		x"5e",	--2957
		x"5f",	--2958
		x"50",	--2959
		x"02",	--2960
		x"40",	--2961
		x"00",	--2962
		x"00",	--2963
		x"40",	--2964
		x"96",	--2965
		x"00",	--2966
		x"40",	--2967
		x"02",	--2968
		x"00",	--2969
		x"53",	--2970
		x"4e",	--2971
		x"02",	--2972
		x"41",	--2973
		x"12",	--2974
		x"42",	--2975
		x"02",	--2976
		x"90",	--2977
		x"00",	--2978
		x"34",	--2979
		x"4b",	--2980
		x"5c",	--2981
		x"5b",	--2982
		x"5c",	--2983
		x"50",	--2984
		x"02",	--2985
		x"4f",	--2986
		x"00",	--2987
		x"4e",	--2988
		x"00",	--2989
		x"4d",	--2990
		x"00",	--2991
		x"53",	--2992
		x"4b",	--2993
		x"02",	--2994
		x"43",	--2995
		x"41",	--2996
		x"41",	--2997
		x"43",	--2998
		x"3f",	--2999
		x"12",	--3000
		x"50",	--3001
		x"ff",	--3002
		x"42",	--3003
		x"02",	--3004
		x"93",	--3005
		x"38",	--3006
		x"92",	--3007
		x"02",	--3008
		x"24",	--3009
		x"40",	--3010
		x"02",	--3011
		x"43",	--3012
		x"3c",	--3013
		x"50",	--3014
		x"00",	--3015
		x"9f",	--3016
		x"ff",	--3017
		x"24",	--3018
		x"53",	--3019
		x"9b",	--3020
		x"23",	--3021
		x"12",	--3022
		x"d6",	--3023
		x"12",	--3024
		x"9b",	--3025
		x"53",	--3026
		x"43",	--3027
		x"50",	--3028
		x"00",	--3029
		x"41",	--3030
		x"41",	--3031
		x"43",	--3032
		x"4e",	--3033
		x"00",	--3034
		x"4e",	--3035
		x"93",	--3036
		x"24",	--3037
		x"53",	--3038
		x"43",	--3039
		x"3c",	--3040
		x"4e",	--3041
		x"93",	--3042
		x"24",	--3043
		x"53",	--3044
		x"92",	--3045
		x"34",	--3046
		x"90",	--3047
		x"00",	--3048
		x"23",	--3049
		x"43",	--3050
		x"ff",	--3051
		x"4f",	--3052
		x"5d",	--3053
		x"51",	--3054
		x"4e",	--3055
		x"00",	--3056
		x"53",	--3057
		x"4e",	--3058
		x"93",	--3059
		x"23",	--3060
		x"4c",	--3061
		x"5e",	--3062
		x"5e",	--3063
		x"5c",	--3064
		x"50",	--3065
		x"02",	--3066
		x"41",	--3067
		x"12",	--3068
		x"00",	--3069
		x"50",	--3070
		x"00",	--3071
		x"41",	--3072
		x"41",	--3073
		x"43",	--3074
		x"3f",	--3075
		x"4e",	--3076
		x"00",	--3077
		x"43",	--3078
		x"41",	--3079
		x"5e",	--3080
		x"5f",	--3081
		x"4e",	--3082
		x"41",	--3083
		x"12",	--3084
		x"12",	--3085
		x"5e",	--3086
		x"5f",	--3087
		x"4e",	--3088
		x"43",	--3089
		x"4c",	--3090
		x"4d",	--3091
		x"5e",	--3092
		x"6f",	--3093
		x"4e",	--3094
		x"4f",	--3095
		x"5a",	--3096
		x"6b",	--3097
		x"5a",	--3098
		x"6b",	--3099
		x"40",	--3100
		x"00",	--3101
		x"43",	--3102
		x"5a",	--3103
		x"6b",	--3104
		x"12",	--3105
		x"d2",	--3106
		x"4e",	--3107
		x"41",	--3108
		x"41",	--3109
		x"41",	--3110
		x"d0",	--3111
		x"02",	--3112
		x"01",	--3113
		x"40",	--3114
		x"0b",	--3115
		x"01",	--3116
		x"43",	--3117
		x"41",	--3118
		x"12",	--3119
		x"4f",	--3120
		x"42",	--3121
		x"02",	--3122
		x"90",	--3123
		x"00",	--3124
		x"34",	--3125
		x"4f",	--3126
		x"5c",	--3127
		x"4c",	--3128
		x"5d",	--3129
		x"5d",	--3130
		x"5d",	--3131
		x"8c",	--3132
		x"50",	--3133
		x"03",	--3134
		x"43",	--3135
		x"00",	--3136
		x"43",	--3137
		x"00",	--3138
		x"43",	--3139
		x"00",	--3140
		x"4b",	--3141
		x"00",	--3142
		x"4e",	--3143
		x"00",	--3144
		x"4f",	--3145
		x"53",	--3146
		x"4e",	--3147
		x"02",	--3148
		x"41",	--3149
		x"41",	--3150
		x"43",	--3151
		x"3f",	--3152
		x"5f",	--3153
		x"4f",	--3154
		x"5c",	--3155
		x"5c",	--3156
		x"5c",	--3157
		x"8f",	--3158
		x"50",	--3159
		x"03",	--3160
		x"43",	--3161
		x"00",	--3162
		x"4e",	--3163
		x"00",	--3164
		x"43",	--3165
		x"00",	--3166
		x"4d",	--3167
		x"00",	--3168
		x"43",	--3169
		x"00",	--3170
		x"43",	--3171
		x"41",	--3172
		x"5f",	--3173
		x"4f",	--3174
		x"5e",	--3175
		x"5e",	--3176
		x"5e",	--3177
		x"8f",	--3178
		x"43",	--3179
		x"03",	--3180
		x"43",	--3181
		x"41",	--3182
		x"12",	--3183
		x"12",	--3184
		x"12",	--3185
		x"12",	--3186
		x"12",	--3187
		x"12",	--3188
		x"12",	--3189
		x"12",	--3190
		x"12",	--3191
		x"93",	--3192
		x"02",	--3193
		x"38",	--3194
		x"40",	--3195
		x"03",	--3196
		x"4a",	--3197
		x"53",	--3198
		x"4a",	--3199
		x"52",	--3200
		x"4a",	--3201
		x"50",	--3202
		x"00",	--3203
		x"43",	--3204
		x"3c",	--3205
		x"53",	--3206
		x"4f",	--3207
		x"00",	--3208
		x"53",	--3209
		x"50",	--3210
		x"00",	--3211
		x"50",	--3212
		x"00",	--3213
		x"50",	--3214
		x"00",	--3215
		x"50",	--3216
		x"00",	--3217
		x"92",	--3218
		x"02",	--3219
		x"34",	--3220
		x"93",	--3221
		x"00",	--3222
		x"27",	--3223
		x"4b",	--3224
		x"9b",	--3225
		x"00",	--3226
		x"2b",	--3227
		x"43",	--3228
		x"00",	--3229
		x"4b",	--3230
		x"00",	--3231
		x"12",	--3232
		x"00",	--3233
		x"93",	--3234
		x"00",	--3235
		x"27",	--3236
		x"47",	--3237
		x"53",	--3238
		x"4f",	--3239
		x"00",	--3240
		x"98",	--3241
		x"2b",	--3242
		x"43",	--3243
		x"00",	--3244
		x"3f",	--3245
		x"f0",	--3246
		x"ff",	--3247
		x"01",	--3248
		x"41",	--3249
		x"41",	--3250
		x"41",	--3251
		x"41",	--3252
		x"41",	--3253
		x"41",	--3254
		x"41",	--3255
		x"41",	--3256
		x"41",	--3257
		x"13",	--3258
		x"4e",	--3259
		x"00",	--3260
		x"43",	--3261
		x"41",	--3262
		x"4f",	--3263
		x"4f",	--3264
		x"4f",	--3265
		x"00",	--3266
		x"41",	--3267
		x"43",	--3268
		x"00",	--3269
		x"41",	--3270
		x"4e",	--3271
		x"00",	--3272
		x"40",	--3273
		x"99",	--3274
		x"12",	--3275
		x"98",	--3276
		x"4f",	--3277
		x"02",	--3278
		x"43",	--3279
		x"41",	--3280
		x"4d",	--3281
		x"4f",	--3282
		x"4e",	--3283
		x"00",	--3284
		x"43",	--3285
		x"4c",	--3286
		x"42",	--3287
		x"02",	--3288
		x"12",	--3289
		x"98",	--3290
		x"41",	--3291
		x"42",	--3292
		x"00",	--3293
		x"f2",	--3294
		x"23",	--3295
		x"4f",	--3296
		x"00",	--3297
		x"43",	--3298
		x"41",	--3299
		x"f0",	--3300
		x"00",	--3301
		x"4f",	--3302
		x"d7",	--3303
		x"11",	--3304
		x"12",	--3305
		x"99",	--3306
		x"41",	--3307
		x"12",	--3308
		x"4f",	--3309
		x"4f",	--3310
		x"11",	--3311
		x"11",	--3312
		x"11",	--3313
		x"11",	--3314
		x"4e",	--3315
		x"12",	--3316
		x"99",	--3317
		x"4b",	--3318
		x"12",	--3319
		x"99",	--3320
		x"41",	--3321
		x"41",	--3322
		x"12",	--3323
		x"12",	--3324
		x"4f",	--3325
		x"40",	--3326
		x"00",	--3327
		x"4a",	--3328
		x"4b",	--3329
		x"f0",	--3330
		x"00",	--3331
		x"24",	--3332
		x"11",	--3333
		x"53",	--3334
		x"23",	--3335
		x"f3",	--3336
		x"24",	--3337
		x"40",	--3338
		x"00",	--3339
		x"12",	--3340
		x"99",	--3341
		x"53",	--3342
		x"93",	--3343
		x"23",	--3344
		x"41",	--3345
		x"41",	--3346
		x"41",	--3347
		x"40",	--3348
		x"00",	--3349
		x"3f",	--3350
		x"12",	--3351
		x"4f",	--3352
		x"4f",	--3353
		x"10",	--3354
		x"11",	--3355
		x"4e",	--3356
		x"12",	--3357
		x"99",	--3358
		x"4b",	--3359
		x"12",	--3360
		x"99",	--3361
		x"41",	--3362
		x"41",	--3363
		x"12",	--3364
		x"12",	--3365
		x"4e",	--3366
		x"4f",	--3367
		x"4f",	--3368
		x"10",	--3369
		x"11",	--3370
		x"4d",	--3371
		x"12",	--3372
		x"99",	--3373
		x"4b",	--3374
		x"12",	--3375
		x"99",	--3376
		x"4b",	--3377
		x"4a",	--3378
		x"10",	--3379
		x"10",	--3380
		x"ec",	--3381
		x"ec",	--3382
		x"4d",	--3383
		x"12",	--3384
		x"99",	--3385
		x"4a",	--3386
		x"12",	--3387
		x"99",	--3388
		x"41",	--3389
		x"41",	--3390
		x"41",	--3391
		x"12",	--3392
		x"12",	--3393
		x"12",	--3394
		x"4f",	--3395
		x"93",	--3396
		x"24",	--3397
		x"4e",	--3398
		x"53",	--3399
		x"43",	--3400
		x"4a",	--3401
		x"5b",	--3402
		x"4d",	--3403
		x"11",	--3404
		x"12",	--3405
		x"99",	--3406
		x"99",	--3407
		x"24",	--3408
		x"53",	--3409
		x"b0",	--3410
		x"00",	--3411
		x"20",	--3412
		x"40",	--3413
		x"00",	--3414
		x"12",	--3415
		x"99",	--3416
		x"3f",	--3417
		x"40",	--3418
		x"00",	--3419
		x"12",	--3420
		x"99",	--3421
		x"3f",	--3422
		x"41",	--3423
		x"41",	--3424
		x"41",	--3425
		x"41",	--3426
		x"12",	--3427
		x"12",	--3428
		x"12",	--3429
		x"4f",	--3430
		x"93",	--3431
		x"24",	--3432
		x"4e",	--3433
		x"53",	--3434
		x"43",	--3435
		x"4a",	--3436
		x"11",	--3437
		x"12",	--3438
		x"99",	--3439
		x"99",	--3440
		x"24",	--3441
		x"53",	--3442
		x"b0",	--3443
		x"00",	--3444
		x"23",	--3445
		x"40",	--3446
		x"00",	--3447
		x"12",	--3448
		x"99",	--3449
		x"4a",	--3450
		x"11",	--3451
		x"12",	--3452
		x"99",	--3453
		x"99",	--3454
		x"23",	--3455
		x"41",	--3456
		x"41",	--3457
		x"41",	--3458
		x"41",	--3459
		x"12",	--3460
		x"12",	--3461
		x"12",	--3462
		x"50",	--3463
		x"ff",	--3464
		x"4f",	--3465
		x"93",	--3466
		x"38",	--3467
		x"90",	--3468
		x"00",	--3469
		x"38",	--3470
		x"43",	--3471
		x"41",	--3472
		x"59",	--3473
		x"40",	--3474
		x"00",	--3475
		x"4b",	--3476
		x"12",	--3477
		x"d2",	--3478
		x"50",	--3479
		x"00",	--3480
		x"4f",	--3481
		x"00",	--3482
		x"53",	--3483
		x"40",	--3484
		x"00",	--3485
		x"4b",	--3486
		x"12",	--3487
		x"d1",	--3488
		x"4f",	--3489
		x"90",	--3490
		x"00",	--3491
		x"37",	--3492
		x"49",	--3493
		x"53",	--3494
		x"51",	--3495
		x"40",	--3496
		x"00",	--3497
		x"4b",	--3498
		x"12",	--3499
		x"d2",	--3500
		x"50",	--3501
		x"00",	--3502
		x"4f",	--3503
		x"00",	--3504
		x"53",	--3505
		x"41",	--3506
		x"5a",	--3507
		x"4f",	--3508
		x"11",	--3509
		x"12",	--3510
		x"99",	--3511
		x"93",	--3512
		x"23",	--3513
		x"50",	--3514
		x"00",	--3515
		x"41",	--3516
		x"41",	--3517
		x"41",	--3518
		x"41",	--3519
		x"40",	--3520
		x"00",	--3521
		x"12",	--3522
		x"99",	--3523
		x"e3",	--3524
		x"53",	--3525
		x"3f",	--3526
		x"43",	--3527
		x"43",	--3528
		x"3f",	--3529
		x"12",	--3530
		x"12",	--3531
		x"12",	--3532
		x"41",	--3533
		x"52",	--3534
		x"4b",	--3535
		x"49",	--3536
		x"93",	--3537
		x"20",	--3538
		x"3c",	--3539
		x"11",	--3540
		x"12",	--3541
		x"99",	--3542
		x"49",	--3543
		x"4a",	--3544
		x"53",	--3545
		x"4a",	--3546
		x"00",	--3547
		x"93",	--3548
		x"24",	--3549
		x"90",	--3550
		x"00",	--3551
		x"23",	--3552
		x"49",	--3553
		x"53",	--3554
		x"49",	--3555
		x"00",	--3556
		x"50",	--3557
		x"ff",	--3558
		x"90",	--3559
		x"00",	--3560
		x"2f",	--3561
		x"4f",	--3562
		x"5f",	--3563
		x"4f",	--3564
		x"d7",	--3565
		x"41",	--3566
		x"41",	--3567
		x"41",	--3568
		x"41",	--3569
		x"4b",	--3570
		x"52",	--3571
		x"4b",	--3572
		x"00",	--3573
		x"4b",	--3574
		x"12",	--3575
		x"9a",	--3576
		x"49",	--3577
		x"3f",	--3578
		x"4b",	--3579
		x"53",	--3580
		x"4b",	--3581
		x"12",	--3582
		x"9a",	--3583
		x"49",	--3584
		x"3f",	--3585
		x"4b",	--3586
		x"53",	--3587
		x"4f",	--3588
		x"49",	--3589
		x"93",	--3590
		x"27",	--3591
		x"53",	--3592
		x"11",	--3593
		x"12",	--3594
		x"99",	--3595
		x"49",	--3596
		x"93",	--3597
		x"23",	--3598
		x"3f",	--3599
		x"4b",	--3600
		x"52",	--3601
		x"4b",	--3602
		x"00",	--3603
		x"4b",	--3604
		x"12",	--3605
		x"9a",	--3606
		x"49",	--3607
		x"3f",	--3608
		x"4b",	--3609
		x"53",	--3610
		x"4b",	--3611
		x"4e",	--3612
		x"10",	--3613
		x"11",	--3614
		x"10",	--3615
		x"11",	--3616
		x"12",	--3617
		x"9a",	--3618
		x"49",	--3619
		x"3f",	--3620
		x"4b",	--3621
		x"53",	--3622
		x"4b",	--3623
		x"12",	--3624
		x"9b",	--3625
		x"49",	--3626
		x"3f",	--3627
		x"4b",	--3628
		x"53",	--3629
		x"4b",	--3630
		x"12",	--3631
		x"99",	--3632
		x"49",	--3633
		x"3f",	--3634
		x"4b",	--3635
		x"53",	--3636
		x"4b",	--3637
		x"12",	--3638
		x"99",	--3639
		x"49",	--3640
		x"3f",	--3641
		x"4b",	--3642
		x"53",	--3643
		x"4b",	--3644
		x"12",	--3645
		x"99",	--3646
		x"49",	--3647
		x"3f",	--3648
		x"40",	--3649
		x"00",	--3650
		x"12",	--3651
		x"99",	--3652
		x"3f",	--3653
		x"12",	--3654
		x"12",	--3655
		x"42",	--3656
		x"02",	--3657
		x"42",	--3658
		x"00",	--3659
		x"05",	--3660
		x"42",	--3661
		x"02",	--3662
		x"90",	--3663
		x"00",	--3664
		x"34",	--3665
		x"53",	--3666
		x"02",	--3667
		x"42",	--3668
		x"02",	--3669
		x"42",	--3670
		x"02",	--3671
		x"9f",	--3672
		x"20",	--3673
		x"53",	--3674
		x"02",	--3675
		x"40",	--3676
		x"00",	--3677
		x"00",	--3678
		x"41",	--3679
		x"41",	--3680
		x"c0",	--3681
		x"00",	--3682
		x"00",	--3683
		x"13",	--3684
		x"43",	--3685
		x"02",	--3686
		x"3f",	--3687
		x"4e",	--3688
		x"4f",	--3689
		x"40",	--3690
		x"36",	--3691
		x"40",	--3692
		x"01",	--3693
		x"12",	--3694
		x"d2",	--3695
		x"53",	--3696
		x"4e",	--3697
		x"00",	--3698
		x"40",	--3699
		x"00",	--3700
		x"00",	--3701
		x"41",	--3702
		x"42",	--3703
		x"02",	--3704
		x"42",	--3705
		x"02",	--3706
		x"9f",	--3707
		x"38",	--3708
		x"42",	--3709
		x"02",	--3710
		x"82",	--3711
		x"02",	--3712
		x"41",	--3713
		x"42",	--3714
		x"02",	--3715
		x"42",	--3716
		x"02",	--3717
		x"40",	--3718
		x"00",	--3719
		x"8d",	--3720
		x"8e",	--3721
		x"41",	--3722
		x"42",	--3723
		x"02",	--3724
		x"4f",	--3725
		x"05",	--3726
		x"42",	--3727
		x"02",	--3728
		x"42",	--3729
		x"02",	--3730
		x"9e",	--3731
		x"24",	--3732
		x"42",	--3733
		x"02",	--3734
		x"90",	--3735
		x"00",	--3736
		x"38",	--3737
		x"43",	--3738
		x"02",	--3739
		x"41",	--3740
		x"53",	--3741
		x"02",	--3742
		x"41",	--3743
		x"43",	--3744
		x"41",	--3745
		x"12",	--3746
		x"12",	--3747
		x"12",	--3748
		x"12",	--3749
		x"12",	--3750
		x"12",	--3751
		x"12",	--3752
		x"12",	--3753
		x"82",	--3754
		x"4e",	--3755
		x"4f",	--3756
		x"4e",	--3757
		x"00",	--3758
		x"4f",	--3759
		x"00",	--3760
		x"4e",	--3761
		x"4f",	--3762
		x"f3",	--3763
		x"f0",	--3764
		x"7f",	--3765
		x"90",	--3766
		x"50",	--3767
		x"38",	--3768
		x"90",	--3769
		x"7f",	--3770
		x"38",	--3771
		x"20",	--3772
		x"93",	--3773
		x"28",	--3774
		x"44",	--3775
		x"45",	--3776
		x"44",	--3777
		x"45",	--3778
		x"12",	--3779
		x"bd",	--3780
		x"40",	--3781
		x"a0",	--3782
		x"93",	--3783
		x"00",	--3784
		x"34",	--3785
		x"40",	--3786
		x"a0",	--3787
		x"20",	--3788
		x"93",	--3789
		x"00",	--3790
		x"2c",	--3791
		x"40",	--3792
		x"a0",	--3793
		x"40",	--3794
		x"0f",	--3795
		x"40",	--3796
		x"3f",	--3797
		x"40",	--3798
		x"a0",	--3799
		x"90",	--3800
		x"3e",	--3801
		x"38",	--3802
		x"4e",	--3803
		x"4f",	--3804
		x"f0",	--3805
		x"7f",	--3806
		x"90",	--3807
		x"3f",	--3808
		x"38",	--3809
		x"3c",	--3810
		x"90",	--3811
		x"31",	--3812
		x"34",	--3813
		x"40",	--3814
		x"f2",	--3815
		x"40",	--3816
		x"71",	--3817
		x"12",	--3818
		x"bd",	--3819
		x"43",	--3820
		x"40",	--3821
		x"3f",	--3822
		x"12",	--3823
		x"c1",	--3824
		x"93",	--3825
		x"24",	--3826
		x"38",	--3827
		x"40",	--3828
		x"a0",	--3829
		x"43",	--3830
		x"43",	--3831
		x"3c",	--3832
		x"90",	--3833
		x"40",	--3834
		x"38",	--3835
		x"3c",	--3836
		x"90",	--3837
		x"3f",	--3838
		x"38",	--3839
		x"43",	--3840
		x"40",	--3841
		x"3f",	--3842
		x"4a",	--3843
		x"4b",	--3844
		x"12",	--3845
		x"bd",	--3846
		x"4e",	--3847
		x"4f",	--3848
		x"43",	--3849
		x"40",	--3850
		x"3f",	--3851
		x"4a",	--3852
		x"4b",	--3853
		x"12",	--3854
		x"bd",	--3855
		x"4e",	--3856
		x"4f",	--3857
		x"48",	--3858
		x"49",	--3859
		x"12",	--3860
		x"bf",	--3861
		x"4e",	--3862
		x"4f",	--3863
		x"43",	--3864
		x"43",	--3865
		x"3c",	--3866
		x"4a",	--3867
		x"4b",	--3868
		x"4a",	--3869
		x"4b",	--3870
		x"12",	--3871
		x"bd",	--3872
		x"43",	--3873
		x"40",	--3874
		x"3f",	--3875
		x"12",	--3876
		x"bd",	--3877
		x"4e",	--3878
		x"4f",	--3879
		x"43",	--3880
		x"40",	--3881
		x"40",	--3882
		x"4a",	--3883
		x"4b",	--3884
		x"12",	--3885
		x"bd",	--3886
		x"4e",	--3887
		x"4f",	--3888
		x"48",	--3889
		x"49",	--3890
		x"12",	--3891
		x"bf",	--3892
		x"4e",	--3893
		x"4f",	--3894
		x"43",	--3895
		x"43",	--3896
		x"3c",	--3897
		x"4a",	--3898
		x"4b",	--3899
		x"43",	--3900
		x"40",	--3901
		x"bf",	--3902
		x"12",	--3903
		x"bf",	--3904
		x"4e",	--3905
		x"4f",	--3906
		x"40",	--3907
		x"00",	--3908
		x"43",	--3909
		x"3c",	--3910
		x"43",	--3911
		x"40",	--3912
		x"3f",	--3913
		x"4a",	--3914
		x"4b",	--3915
		x"12",	--3916
		x"bd",	--3917
		x"4e",	--3918
		x"4f",	--3919
		x"43",	--3920
		x"40",	--3921
		x"3f",	--3922
		x"4a",	--3923
		x"4b",	--3924
		x"12",	--3925
		x"bd",	--3926
		x"43",	--3927
		x"40",	--3928
		x"3f",	--3929
		x"12",	--3930
		x"bd",	--3931
		x"4e",	--3932
		x"4f",	--3933
		x"48",	--3934
		x"49",	--3935
		x"12",	--3936
		x"bf",	--3937
		x"4e",	--3938
		x"4f",	--3939
		x"43",	--3940
		x"43",	--3941
		x"44",	--3942
		x"45",	--3943
		x"44",	--3944
		x"45",	--3945
		x"12",	--3946
		x"bd",	--3947
		x"4e",	--3948
		x"4f",	--3949
		x"4e",	--3950
		x"4f",	--3951
		x"12",	--3952
		x"bd",	--3953
		x"4e",	--3954
		x"4f",	--3955
		x"40",	--3956
		x"69",	--3957
		x"40",	--3958
		x"3c",	--3959
		x"12",	--3960
		x"bd",	--3961
		x"40",	--3962
		x"da",	--3963
		x"40",	--3964
		x"3d",	--3965
		x"12",	--3966
		x"bd",	--3967
		x"4e",	--3968
		x"4f",	--3969
		x"4a",	--3970
		x"4b",	--3971
		x"12",	--3972
		x"bd",	--3973
		x"40",	--3974
		x"6b",	--3975
		x"40",	--3976
		x"3d",	--3977
		x"12",	--3978
		x"bd",	--3979
		x"4e",	--3980
		x"4f",	--3981
		x"4a",	--3982
		x"4b",	--3983
		x"12",	--3984
		x"bd",	--3985
		x"40",	--3986
		x"2e",	--3987
		x"40",	--3988
		x"3d",	--3989
		x"12",	--3990
		x"bd",	--3991
		x"4e",	--3992
		x"4f",	--3993
		x"4a",	--3994
		x"4b",	--3995
		x"12",	--3996
		x"bd",	--3997
		x"40",	--3998
		x"49",	--3999
		x"40",	--4000
		x"3e",	--4001
		x"12",	--4002
		x"bd",	--4003
		x"4e",	--4004
		x"4f",	--4005
		x"4a",	--4006
		x"4b",	--4007
		x"12",	--4008
		x"bd",	--4009
		x"40",	--4010
		x"aa",	--4011
		x"40",	--4012
		x"3e",	--4013
		x"12",	--4014
		x"bd",	--4015
		x"4e",	--4016
		x"4f",	--4017
		x"48",	--4018
		x"49",	--4019
		x"12",	--4020
		x"bd",	--4021
		x"4e",	--4022
		x"00",	--4023
		x"4f",	--4024
		x"00",	--4025
		x"40",	--4026
		x"a2",	--4027
		x"40",	--4028
		x"bd",	--4029
		x"4a",	--4030
		x"4b",	--4031
		x"12",	--4032
		x"bd",	--4033
		x"40",	--4034
		x"f1",	--4035
		x"40",	--4036
		x"3d",	--4037
		x"12",	--4038
		x"bd",	--4039
		x"4e",	--4040
		x"4f",	--4041
		x"4a",	--4042
		x"4b",	--4043
		x"12",	--4044
		x"bd",	--4045
		x"40",	--4046
		x"87",	--4047
		x"40",	--4048
		x"3d",	--4049
		x"12",	--4050
		x"bd",	--4051
		x"4e",	--4052
		x"4f",	--4053
		x"4a",	--4054
		x"4b",	--4055
		x"12",	--4056
		x"bd",	--4057
		x"40",	--4058
		x"8e",	--4059
		x"40",	--4060
		x"3d",	--4061
		x"12",	--4062
		x"bd",	--4063
		x"4e",	--4064
		x"4f",	--4065
		x"4a",	--4066
		x"4b",	--4067
		x"12",	--4068
		x"bd",	--4069
		x"40",	--4070
		x"cc",	--4071
		x"40",	--4072
		x"3e",	--4073
		x"12",	--4074
		x"bd",	--4075
		x"4e",	--4076
		x"4f",	--4077
		x"4a",	--4078
		x"4b",	--4079
		x"12",	--4080
		x"bd",	--4081
		x"4e",	--4082
		x"4f",	--4083
		x"93",	--4084
		x"20",	--4085
		x"93",	--4086
		x"20",	--4087
		x"4e",	--4088
		x"4f",	--4089
		x"41",	--4090
		x"00",	--4091
		x"41",	--4092
		x"00",	--4093
		x"12",	--4094
		x"bd",	--4095
		x"4e",	--4096
		x"4f",	--4097
		x"44",	--4098
		x"45",	--4099
		x"12",	--4100
		x"bd",	--4101
		x"4e",	--4102
		x"4f",	--4103
		x"44",	--4104
		x"45",	--4105
		x"12",	--4106
		x"bd",	--4107
		x"4e",	--4108
		x"4f",	--4109
		x"3c",	--4110
		x"46",	--4111
		x"5b",	--4112
		x"5b",	--4113
		x"4b",	--4114
		x"50",	--4115
		x"d7",	--4116
		x"48",	--4117
		x"49",	--4118
		x"41",	--4119
		x"00",	--4120
		x"41",	--4121
		x"00",	--4122
		x"12",	--4123
		x"bd",	--4124
		x"4e",	--4125
		x"4f",	--4126
		x"44",	--4127
		x"45",	--4128
		x"12",	--4129
		x"bd",	--4130
		x"4b",	--4131
		x"d7",	--4132
		x"4b",	--4133
		x"d7",	--4134
		x"12",	--4135
		x"bd",	--4136
		x"44",	--4137
		x"45",	--4138
		x"12",	--4139
		x"bd",	--4140
		x"4e",	--4141
		x"4f",	--4142
		x"47",	--4143
		x"47",	--4144
		x"00",	--4145
		x"12",	--4146
		x"bd",	--4147
		x"4e",	--4148
		x"4f",	--4149
		x"93",	--4150
		x"00",	--4151
		x"34",	--4152
		x"e0",	--4153
		x"80",	--4154
		x"3c",	--4155
		x"40",	--4156
		x"0f",	--4157
		x"40",	--4158
		x"bf",	--4159
		x"44",	--4160
		x"45",	--4161
		x"52",	--4162
		x"41",	--4163
		x"41",	--4164
		x"41",	--4165
		x"41",	--4166
		x"41",	--4167
		x"41",	--4168
		x"41",	--4169
		x"41",	--4170
		x"41",	--4171
		x"12",	--4172
		x"9d",	--4173
		x"41",	--4174
		x"12",	--4175
		x"12",	--4176
		x"82",	--4177
		x"4e",	--4178
		x"4f",	--4179
		x"f3",	--4180
		x"f0",	--4181
		x"7f",	--4182
		x"90",	--4183
		x"3f",	--4184
		x"38",	--4185
		x"90",	--4186
		x"3f",	--4187
		x"34",	--4188
		x"90",	--4189
		x"0f",	--4190
		x"2c",	--4191
		x"12",	--4192
		x"43",	--4193
		x"43",	--4194
		x"3c",	--4195
		x"90",	--4196
		x"7f",	--4197
		x"38",	--4198
		x"4e",	--4199
		x"4f",	--4200
		x"12",	--4201
		x"bd",	--4202
		x"3c",	--4203
		x"41",	--4204
		x"12",	--4205
		x"a3",	--4206
		x"4e",	--4207
		x"4f",	--4208
		x"f0",	--4209
		x"00",	--4210
		x"f3",	--4211
		x"41",	--4212
		x"00",	--4213
		x"41",	--4214
		x"00",	--4215
		x"41",	--4216
		x"41",	--4217
		x"00",	--4218
		x"93",	--4219
		x"20",	--4220
		x"93",	--4221
		x"24",	--4222
		x"93",	--4223
		x"20",	--4224
		x"93",	--4225
		x"24",	--4226
		x"41",	--4227
		x"41",	--4228
		x"00",	--4229
		x"93",	--4230
		x"20",	--4231
		x"93",	--4232
		x"20",	--4233
		x"12",	--4234
		x"12",	--4235
		x"b6",	--4236
		x"53",	--4237
		x"3c",	--4238
		x"12",	--4239
		x"a1",	--4240
		x"3c",	--4241
		x"12",	--4242
		x"12",	--4243
		x"b6",	--4244
		x"53",	--4245
		x"3c",	--4246
		x"12",	--4247
		x"a1",	--4248
		x"e0",	--4249
		x"80",	--4250
		x"52",	--4251
		x"41",	--4252
		x"41",	--4253
		x"41",	--4254
		x"12",	--4255
		x"a0",	--4256
		x"41",	--4257
		x"12",	--4258
		x"12",	--4259
		x"12",	--4260
		x"12",	--4261
		x"12",	--4262
		x"12",	--4263
		x"12",	--4264
		x"12",	--4265
		x"82",	--4266
		x"4e",	--4267
		x"4f",	--4268
		x"4c",	--4269
		x"4d",	--4270
		x"4e",	--4271
		x"4f",	--4272
		x"f3",	--4273
		x"f0",	--4274
		x"7f",	--4275
		x"90",	--4276
		x"32",	--4277
		x"34",	--4278
		x"12",	--4279
		x"c3",	--4280
		x"93",	--4281
		x"24",	--4282
		x"46",	--4283
		x"47",	--4284
		x"46",	--4285
		x"47",	--4286
		x"12",	--4287
		x"bd",	--4288
		x"4e",	--4289
		x"4f",	--4290
		x"40",	--4291
		x"d7",	--4292
		x"40",	--4293
		x"ad",	--4294
		x"12",	--4295
		x"bd",	--4296
		x"40",	--4297
		x"74",	--4298
		x"40",	--4299
		x"31",	--4300
		x"12",	--4301
		x"bd",	--4302
		x"4e",	--4303
		x"4f",	--4304
		x"48",	--4305
		x"49",	--4306
		x"12",	--4307
		x"bd",	--4308
		x"40",	--4309
		x"f2",	--4310
		x"40",	--4311
		x"34",	--4312
		x"12",	--4313
		x"bd",	--4314
		x"4e",	--4315
		x"4f",	--4316
		x"48",	--4317
		x"49",	--4318
		x"12",	--4319
		x"bd",	--4320
		x"40",	--4321
		x"0d",	--4322
		x"40",	--4323
		x"37",	--4324
		x"12",	--4325
		x"bd",	--4326
		x"4e",	--4327
		x"4f",	--4328
		x"48",	--4329
		x"49",	--4330
		x"12",	--4331
		x"bd",	--4332
		x"40",	--4333
		x"0b",	--4334
		x"40",	--4335
		x"3a",	--4336
		x"12",	--4337
		x"bd",	--4338
		x"4e",	--4339
		x"4f",	--4340
		x"48",	--4341
		x"49",	--4342
		x"12",	--4343
		x"bd",	--4344
		x"40",	--4345
		x"aa",	--4346
		x"40",	--4347
		x"3d",	--4348
		x"12",	--4349
		x"bd",	--4350
		x"4e",	--4351
		x"4f",	--4352
		x"48",	--4353
		x"49",	--4354
		x"12",	--4355
		x"bd",	--4356
		x"4e",	--4357
		x"00",	--4358
		x"4f",	--4359
		x"00",	--4360
		x"90",	--4361
		x"3e",	--4362
		x"38",	--4363
		x"90",	--4364
		x"3e",	--4365
		x"34",	--4366
		x"90",	--4367
		x"99",	--4368
		x"2c",	--4369
		x"43",	--4370
		x"40",	--4371
		x"3f",	--4372
		x"48",	--4373
		x"49",	--4374
		x"12",	--4375
		x"bd",	--4376
		x"4e",	--4377
		x"4f",	--4378
		x"41",	--4379
		x"41",	--4380
		x"00",	--4381
		x"48",	--4382
		x"49",	--4383
		x"12",	--4384
		x"bd",	--4385
		x"4e",	--4386
		x"4f",	--4387
		x"44",	--4388
		x"45",	--4389
		x"46",	--4390
		x"47",	--4391
		x"12",	--4392
		x"bd",	--4393
		x"4e",	--4394
		x"4f",	--4395
		x"48",	--4396
		x"49",	--4397
		x"12",	--4398
		x"bd",	--4399
		x"4e",	--4400
		x"4f",	--4401
		x"4a",	--4402
		x"4b",	--4403
		x"12",	--4404
		x"bd",	--4405
		x"4e",	--4406
		x"4f",	--4407
		x"43",	--4408
		x"40",	--4409
		x"3f",	--4410
		x"3c",	--4411
		x"90",	--4412
		x"3f",	--4413
		x"38",	--4414
		x"90",	--4415
		x"3f",	--4416
		x"34",	--4417
		x"93",	--4418
		x"2c",	--4419
		x"53",	--4420
		x"60",	--4421
		x"ff",	--4422
		x"3c",	--4423
		x"43",	--4424
		x"40",	--4425
		x"3e",	--4426
		x"4a",	--4427
		x"4b",	--4428
		x"43",	--4429
		x"40",	--4430
		x"3f",	--4431
		x"12",	--4432
		x"bd",	--4433
		x"4e",	--4434
		x"00",	--4435
		x"4f",	--4436
		x"00",	--4437
		x"43",	--4438
		x"40",	--4439
		x"3f",	--4440
		x"48",	--4441
		x"49",	--4442
		x"12",	--4443
		x"bd",	--4444
		x"4a",	--4445
		x"4b",	--4446
		x"12",	--4447
		x"bd",	--4448
		x"4e",	--4449
		x"4f",	--4450
		x"41",	--4451
		x"41",	--4452
		x"00",	--4453
		x"48",	--4454
		x"49",	--4455
		x"12",	--4456
		x"bd",	--4457
		x"4e",	--4458
		x"4f",	--4459
		x"44",	--4460
		x"45",	--4461
		x"46",	--4462
		x"47",	--4463
		x"12",	--4464
		x"bd",	--4465
		x"4e",	--4466
		x"4f",	--4467
		x"48",	--4468
		x"49",	--4469
		x"12",	--4470
		x"bd",	--4471
		x"4e",	--4472
		x"4f",	--4473
		x"4a",	--4474
		x"4b",	--4475
		x"12",	--4476
		x"bd",	--4477
		x"4e",	--4478
		x"4f",	--4479
		x"41",	--4480
		x"00",	--4481
		x"41",	--4482
		x"00",	--4483
		x"12",	--4484
		x"bd",	--4485
		x"3c",	--4486
		x"43",	--4487
		x"40",	--4488
		x"3f",	--4489
		x"52",	--4490
		x"41",	--4491
		x"41",	--4492
		x"41",	--4493
		x"41",	--4494
		x"41",	--4495
		x"41",	--4496
		x"41",	--4497
		x"41",	--4498
		x"41",	--4499
		x"12",	--4500
		x"12",	--4501
		x"12",	--4502
		x"12",	--4503
		x"12",	--4504
		x"12",	--4505
		x"12",	--4506
		x"12",	--4507
		x"50",	--4508
		x"ff",	--4509
		x"4d",	--4510
		x"00",	--4511
		x"4e",	--4512
		x"00",	--4513
		x"4f",	--4514
		x"00",	--4515
		x"4e",	--4516
		x"4f",	--4517
		x"f3",	--4518
		x"f0",	--4519
		x"7f",	--4520
		x"90",	--4521
		x"3f",	--4522
		x"38",	--4523
		x"90",	--4524
		x"3f",	--4525
		x"34",	--4526
		x"90",	--4527
		x"0f",	--4528
		x"2c",	--4529
		x"41",	--4530
		x"00",	--4531
		x"4e",	--4532
		x"00",	--4533
		x"4f",	--4534
		x"00",	--4535
		x"43",	--4536
		x"00",	--4537
		x"43",	--4538
		x"00",	--4539
		x"40",	--4540
		x"a7",	--4541
		x"90",	--4542
		x"40",	--4543
		x"38",	--4544
		x"90",	--4545
		x"40",	--4546
		x"34",	--4547
		x"90",	--4548
		x"cb",	--4549
		x"2c",	--4550
		x"93",	--4551
		x"00",	--4552
		x"38",	--4553
		x"20",	--4554
		x"93",	--4555
		x"00",	--4556
		x"28",	--4557
		x"40",	--4558
		x"0f",	--4559
		x"40",	--4560
		x"3f",	--4561
		x"12",	--4562
		x"bd",	--4563
		x"4e",	--4564
		x"4f",	--4565
		x"f0",	--4566
		x"ff",	--4567
		x"f3",	--4568
		x"90",	--4569
		x"0f",	--4570
		x"20",	--4571
		x"90",	--4572
		x"3f",	--4573
		x"24",	--4574
		x"40",	--4575
		x"44",	--4576
		x"40",	--4577
		x"37",	--4578
		x"48",	--4579
		x"49",	--4580
		x"12",	--4581
		x"bd",	--4582
		x"4e",	--4583
		x"4f",	--4584
		x"41",	--4585
		x"00",	--4586
		x"4c",	--4587
		x"00",	--4588
		x"4d",	--4589
		x"00",	--4590
		x"48",	--4591
		x"49",	--4592
		x"12",	--4593
		x"bd",	--4594
		x"40",	--4595
		x"44",	--4596
		x"40",	--4597
		x"37",	--4598
		x"3c",	--4599
		x"40",	--4600
		x"44",	--4601
		x"40",	--4602
		x"37",	--4603
		x"12",	--4604
		x"bd",	--4605
		x"4e",	--4606
		x"4f",	--4607
		x"40",	--4608
		x"a3",	--4609
		x"40",	--4610
		x"2e",	--4611
		x"12",	--4612
		x"bd",	--4613
		x"4e",	--4614
		x"4f",	--4615
		x"41",	--4616
		x"00",	--4617
		x"4c",	--4618
		x"00",	--4619
		x"4d",	--4620
		x"00",	--4621
		x"4a",	--4622
		x"4b",	--4623
		x"12",	--4624
		x"bd",	--4625
		x"40",	--4626
		x"a3",	--4627
		x"40",	--4628
		x"2e",	--4629
		x"12",	--4630
		x"bd",	--4631
		x"41",	--4632
		x"00",	--4633
		x"4e",	--4634
		x"00",	--4635
		x"4f",	--4636
		x"00",	--4637
		x"43",	--4638
		x"43",	--4639
		x"40",	--4640
		x"a8",	--4641
		x"40",	--4642
		x"0f",	--4643
		x"40",	--4644
		x"3f",	--4645
		x"12",	--4646
		x"bd",	--4647
		x"4e",	--4648
		x"4f",	--4649
		x"f0",	--4650
		x"ff",	--4651
		x"f3",	--4652
		x"90",	--4653
		x"0f",	--4654
		x"20",	--4655
		x"90",	--4656
		x"3f",	--4657
		x"24",	--4658
		x"40",	--4659
		x"44",	--4660
		x"40",	--4661
		x"37",	--4662
		x"48",	--4663
		x"49",	--4664
		x"12",	--4665
		x"bd",	--4666
		x"4e",	--4667
		x"4f",	--4668
		x"41",	--4669
		x"00",	--4670
		x"4c",	--4671
		x"00",	--4672
		x"4d",	--4673
		x"00",	--4674
		x"48",	--4675
		x"49",	--4676
		x"12",	--4677
		x"bd",	--4678
		x"40",	--4679
		x"44",	--4680
		x"40",	--4681
		x"37",	--4682
		x"3c",	--4683
		x"40",	--4684
		x"44",	--4685
		x"40",	--4686
		x"37",	--4687
		x"12",	--4688
		x"bd",	--4689
		x"4e",	--4690
		x"4f",	--4691
		x"40",	--4692
		x"a3",	--4693
		x"40",	--4694
		x"2e",	--4695
		x"12",	--4696
		x"bd",	--4697
		x"4e",	--4698
		x"4f",	--4699
		x"41",	--4700
		x"00",	--4701
		x"4c",	--4702
		x"00",	--4703
		x"4d",	--4704
		x"00",	--4705
		x"4a",	--4706
		x"4b",	--4707
		x"12",	--4708
		x"bd",	--4709
		x"40",	--4710
		x"a3",	--4711
		x"40",	--4712
		x"2e",	--4713
		x"12",	--4714
		x"bd",	--4715
		x"41",	--4716
		x"00",	--4717
		x"4e",	--4718
		x"00",	--4719
		x"4f",	--4720
		x"00",	--4721
		x"43",	--4722
		x"43",	--4723
		x"40",	--4724
		x"a8",	--4725
		x"90",	--4726
		x"43",	--4727
		x"38",	--4728
		x"90",	--4729
		x"43",	--4730
		x"38",	--4731
		x"40",	--4732
		x"a7",	--4733
		x"90",	--4734
		x"0f",	--4735
		x"28",	--4736
		x"40",	--4737
		x"a7",	--4738
		x"4e",	--4739
		x"4f",	--4740
		x"f0",	--4741
		x"7f",	--4742
		x"40",	--4743
		x"f9",	--4744
		x"40",	--4745
		x"3f",	--4746
		x"48",	--4747
		x"49",	--4748
		x"12",	--4749
		x"bd",	--4750
		x"43",	--4751
		x"40",	--4752
		x"3f",	--4753
		x"12",	--4754
		x"bd",	--4755
		x"12",	--4756
		x"c3",	--4757
		x"4e",	--4758
		x"4f",	--4759
		x"12",	--4760
		x"c2",	--4761
		x"4e",	--4762
		x"00",	--4763
		x"4f",	--4764
		x"00",	--4765
		x"40",	--4766
		x"0f",	--4767
		x"40",	--4768
		x"3f",	--4769
		x"12",	--4770
		x"bd",	--4771
		x"4e",	--4772
		x"4f",	--4773
		x"48",	--4774
		x"49",	--4775
		x"12",	--4776
		x"bd",	--4777
		x"4e",	--4778
		x"4f",	--4779
		x"40",	--4780
		x"44",	--4781
		x"40",	--4782
		x"37",	--4783
		x"41",	--4784
		x"00",	--4785
		x"41",	--4786
		x"00",	--4787
		x"12",	--4788
		x"bd",	--4789
		x"4e",	--4790
		x"00",	--4791
		x"4f",	--4792
		x"00",	--4793
		x"93",	--4794
		x"38",	--4795
		x"93",	--4796
		x"34",	--4797
		x"90",	--4798
		x"00",	--4799
		x"2c",	--4800
		x"4a",	--4801
		x"4b",	--4802
		x"f0",	--4803
		x"ff",	--4804
		x"f3",	--4805
		x"46",	--4806
		x"53",	--4807
		x"5f",	--4808
		x"5f",	--4809
		x"50",	--4810
		x"d7",	--4811
		x"9f",	--4812
		x"20",	--4813
		x"9f",	--4814
		x"00",	--4815
		x"24",	--4816
		x"41",	--4817
		x"00",	--4818
		x"41",	--4819
		x"00",	--4820
		x"40",	--4821
		x"a7",	--4822
		x"41",	--4823
		x"00",	--4824
		x"41",	--4825
		x"00",	--4826
		x"44",	--4827
		x"45",	--4828
		x"12",	--4829
		x"bd",	--4830
		x"4e",	--4831
		x"4f",	--4832
		x"41",	--4833
		x"00",	--4834
		x"48",	--4835
		x"00",	--4836
		x"49",	--4837
		x"00",	--4838
		x"4b",	--4839
		x"00",	--4840
		x"4b",	--4841
		x"10",	--4842
		x"11",	--4843
		x"10",	--4844
		x"11",	--4845
		x"4d",	--4846
		x"00",	--4847
		x"40",	--4848
		x"00",	--4849
		x"4f",	--4850
		x"41",	--4851
		x"00",	--4852
		x"41",	--4853
		x"00",	--4854
		x"11",	--4855
		x"10",	--4856
		x"53",	--4857
		x"23",	--4858
		x"4e",	--4859
		x"00",	--4860
		x"4f",	--4861
		x"00",	--4862
		x"4c",	--4863
		x"43",	--4864
		x"40",	--4865
		x"00",	--4866
		x"c3",	--4867
		x"10",	--4868
		x"10",	--4869
		x"53",	--4870
		x"23",	--4871
		x"f0",	--4872
		x"00",	--4873
		x"f3",	--4874
		x"41",	--4875
		x"00",	--4876
		x"41",	--4877
		x"00",	--4878
		x"8a",	--4879
		x"7b",	--4880
		x"93",	--4881
		x"38",	--4882
		x"20",	--4883
		x"90",	--4884
		x"00",	--4885
		x"28",	--4886
		x"40",	--4887
		x"44",	--4888
		x"40",	--4889
		x"37",	--4890
		x"41",	--4891
		x"00",	--4892
		x"41",	--4893
		x"00",	--4894
		x"12",	--4895
		x"bd",	--4896
		x"4e",	--4897
		x"4f",	--4898
		x"4e",	--4899
		x"4f",	--4900
		x"44",	--4901
		x"45",	--4902
		x"12",	--4903
		x"bd",	--4904
		x"4e",	--4905
		x"00",	--4906
		x"4f",	--4907
		x"00",	--4908
		x"4e",	--4909
		x"4f",	--4910
		x"44",	--4911
		x"45",	--4912
		x"12",	--4913
		x"bd",	--4914
		x"48",	--4915
		x"49",	--4916
		x"12",	--4917
		x"bd",	--4918
		x"4e",	--4919
		x"4f",	--4920
		x"40",	--4921
		x"a3",	--4922
		x"40",	--4923
		x"2e",	--4924
		x"41",	--4925
		x"00",	--4926
		x"41",	--4927
		x"00",	--4928
		x"12",	--4929
		x"bd",	--4930
		x"48",	--4931
		x"49",	--4932
		x"12",	--4933
		x"bd",	--4934
		x"4e",	--4935
		x"00",	--4936
		x"4f",	--4937
		x"00",	--4938
		x"4e",	--4939
		x"4f",	--4940
		x"41",	--4941
		x"00",	--4942
		x"41",	--4943
		x"00",	--4944
		x"12",	--4945
		x"bd",	--4946
		x"4e",	--4947
		x"4f",	--4948
		x"41",	--4949
		x"00",	--4950
		x"4a",	--4951
		x"00",	--4952
		x"4b",	--4953
		x"00",	--4954
		x"4f",	--4955
		x"43",	--4956
		x"40",	--4957
		x"00",	--4958
		x"c3",	--4959
		x"10",	--4960
		x"10",	--4961
		x"53",	--4962
		x"23",	--4963
		x"f0",	--4964
		x"00",	--4965
		x"f3",	--4966
		x"41",	--4967
		x"00",	--4968
		x"41",	--4969
		x"00",	--4970
		x"8a",	--4971
		x"7b",	--4972
		x"4d",	--4973
		x"4e",	--4974
		x"93",	--4975
		x"38",	--4976
		x"20",	--4977
		x"90",	--4978
		x"00",	--4979
		x"28",	--4980
		x"40",	--4981
		x"a3",	--4982
		x"40",	--4983
		x"2e",	--4984
		x"41",	--4985
		x"00",	--4986
		x"41",	--4987
		x"00",	--4988
		x"12",	--4989
		x"bd",	--4990
		x"4e",	--4991
		x"4f",	--4992
		x"4e",	--4993
		x"4f",	--4994
		x"41",	--4995
		x"00",	--4996
		x"41",	--4997
		x"00",	--4998
		x"12",	--4999
		x"bd",	--5000
		x"4e",	--5001
		x"4f",	--5002
		x"4e",	--5003
		x"4f",	--5004
		x"41",	--5005
		x"00",	--5006
		x"41",	--5007
		x"00",	--5008
		x"12",	--5009
		x"bd",	--5010
		x"4a",	--5011
		x"4b",	--5012
		x"12",	--5013
		x"bd",	--5014
		x"4e",	--5015
		x"4f",	--5016
		x"40",	--5017
		x"31",	--5018
		x"40",	--5019
		x"24",	--5020
		x"41",	--5021
		x"00",	--5022
		x"41",	--5023
		x"00",	--5024
		x"12",	--5025
		x"bd",	--5026
		x"4a",	--5027
		x"4b",	--5028
		x"12",	--5029
		x"bd",	--5030
		x"4e",	--5031
		x"00",	--5032
		x"4f",	--5033
		x"00",	--5034
		x"4e",	--5035
		x"4f",	--5036
		x"44",	--5037
		x"45",	--5038
		x"12",	--5039
		x"bd",	--5040
		x"41",	--5041
		x"00",	--5042
		x"4e",	--5043
		x"00",	--5044
		x"4f",	--5045
		x"00",	--5046
		x"3c",	--5047
		x"41",	--5048
		x"00",	--5049
		x"41",	--5050
		x"00",	--5051
		x"41",	--5052
		x"00",	--5053
		x"4e",	--5054
		x"4e",	--5055
		x"00",	--5056
		x"48",	--5057
		x"49",	--5058
		x"44",	--5059
		x"45",	--5060
		x"12",	--5061
		x"bd",	--5062
		x"41",	--5063
		x"00",	--5064
		x"41",	--5065
		x"00",	--5066
		x"12",	--5067
		x"bd",	--5068
		x"4e",	--5069
		x"4f",	--5070
		x"41",	--5071
		x"00",	--5072
		x"4a",	--5073
		x"00",	--5074
		x"4b",	--5075
		x"00",	--5076
		x"93",	--5077
		x"00",	--5078
		x"34",	--5079
		x"48",	--5080
		x"49",	--5081
		x"e0",	--5082
		x"80",	--5083
		x"4d",	--5084
		x"00",	--5085
		x"4e",	--5086
		x"00",	--5087
		x"4a",	--5088
		x"4b",	--5089
		x"e0",	--5090
		x"80",	--5091
		x"4d",	--5092
		x"00",	--5093
		x"4e",	--5094
		x"00",	--5095
		x"3c",	--5096
		x"90",	--5097
		x"7f",	--5098
		x"38",	--5099
		x"4e",	--5100
		x"4f",	--5101
		x"12",	--5102
		x"bd",	--5103
		x"41",	--5104
		x"00",	--5105
		x"4e",	--5106
		x"00",	--5107
		x"4f",	--5108
		x"00",	--5109
		x"4e",	--5110
		x"00",	--5111
		x"4f",	--5112
		x"00",	--5113
		x"43",	--5114
		x"43",	--5115
		x"3c",	--5116
		x"4b",	--5117
		x"4b",	--5118
		x"10",	--5119
		x"11",	--5120
		x"10",	--5121
		x"11",	--5122
		x"40",	--5123
		x"00",	--5124
		x"11",	--5125
		x"10",	--5126
		x"53",	--5127
		x"23",	--5128
		x"4c",	--5129
		x"50",	--5130
		x"ff",	--5131
		x"43",	--5132
		x"43",	--5133
		x"49",	--5134
		x"40",	--5135
		x"00",	--5136
		x"5c",	--5137
		x"6d",	--5138
		x"53",	--5139
		x"23",	--5140
		x"8c",	--5141
		x"7d",	--5142
		x"4a",	--5143
		x"4b",	--5144
		x"12",	--5145
		x"c3",	--5146
		x"12",	--5147
		x"c2",	--5148
		x"4e",	--5149
		x"4f",	--5150
		x"4e",	--5151
		x"00",	--5152
		x"4f",	--5153
		x"00",	--5154
		x"4a",	--5155
		x"4b",	--5156
		x"12",	--5157
		x"bd",	--5158
		x"43",	--5159
		x"40",	--5160
		x"43",	--5161
		x"12",	--5162
		x"bd",	--5163
		x"4e",	--5164
		x"4f",	--5165
		x"12",	--5166
		x"c3",	--5167
		x"12",	--5168
		x"c2",	--5169
		x"4e",	--5170
		x"4f",	--5171
		x"4e",	--5172
		x"00",	--5173
		x"4f",	--5174
		x"00",	--5175
		x"4a",	--5176
		x"4b",	--5177
		x"12",	--5178
		x"bd",	--5179
		x"43",	--5180
		x"40",	--5181
		x"43",	--5182
		x"12",	--5183
		x"bd",	--5184
		x"4e",	--5185
		x"00",	--5186
		x"4f",	--5187
		x"00",	--5188
		x"41",	--5189
		x"52",	--5190
		x"40",	--5191
		x"00",	--5192
		x"3c",	--5193
		x"53",	--5194
		x"82",	--5195
		x"43",	--5196
		x"43",	--5197
		x"48",	--5198
		x"00",	--5199
		x"48",	--5200
		x"00",	--5201
		x"12",	--5202
		x"c1",	--5203
		x"93",	--5204
		x"27",	--5205
		x"12",	--5206
		x"d8",	--5207
		x"12",	--5208
		x"4a",	--5209
		x"49",	--5210
		x"41",	--5211
		x"00",	--5212
		x"41",	--5213
		x"52",	--5214
		x"12",	--5215
		x"a9",	--5216
		x"52",	--5217
		x"4f",	--5218
		x"10",	--5219
		x"11",	--5220
		x"10",	--5221
		x"11",	--5222
		x"4f",	--5223
		x"93",	--5224
		x"00",	--5225
		x"34",	--5226
		x"41",	--5227
		x"00",	--5228
		x"e0",	--5229
		x"80",	--5230
		x"00",	--5231
		x"e0",	--5232
		x"80",	--5233
		x"00",	--5234
		x"e3",	--5235
		x"e3",	--5236
		x"53",	--5237
		x"63",	--5238
		x"46",	--5239
		x"47",	--5240
		x"50",	--5241
		x"00",	--5242
		x"41",	--5243
		x"41",	--5244
		x"41",	--5245
		x"41",	--5246
		x"41",	--5247
		x"41",	--5248
		x"41",	--5249
		x"41",	--5250
		x"41",	--5251
		x"12",	--5252
		x"12",	--5253
		x"12",	--5254
		x"12",	--5255
		x"12",	--5256
		x"12",	--5257
		x"12",	--5258
		x"12",	--5259
		x"50",	--5260
		x"fe",	--5261
		x"4f",	--5262
		x"01",	--5263
		x"4e",	--5264
		x"01",	--5265
		x"4c",	--5266
		x"01",	--5267
		x"41",	--5268
		x"01",	--5269
		x"5a",	--5270
		x"43",	--5271
		x"01",	--5272
		x"43",	--5273
		x"01",	--5274
		x"4a",	--5275
		x"db",	--5276
		x"01",	--5277
		x"41",	--5278
		x"01",	--5279
		x"10",	--5280
		x"11",	--5281
		x"10",	--5282
		x"11",	--5283
		x"4a",	--5284
		x"01",	--5285
		x"4c",	--5286
		x"53",	--5287
		x"4a",	--5288
		x"01",	--5289
		x"10",	--5290
		x"11",	--5291
		x"10",	--5292
		x"11",	--5293
		x"4a",	--5294
		x"01",	--5295
		x"4d",	--5296
		x"50",	--5297
		x"ff",	--5298
		x"93",	--5299
		x"34",	--5300
		x"50",	--5301
		x"00",	--5302
		x"11",	--5303
		x"11",	--5304
		x"11",	--5305
		x"4a",	--5306
		x"10",	--5307
		x"11",	--5308
		x"10",	--5309
		x"11",	--5310
		x"4a",	--5311
		x"01",	--5312
		x"48",	--5313
		x"01",	--5314
		x"34",	--5315
		x"43",	--5316
		x"01",	--5317
		x"43",	--5318
		x"01",	--5319
		x"4d",	--5320
		x"10",	--5321
		x"11",	--5322
		x"10",	--5323
		x"11",	--5324
		x"4d",	--5325
		x"41",	--5326
		x"01",	--5327
		x"41",	--5328
		x"01",	--5329
		x"e3",	--5330
		x"e3",	--5331
		x"5a",	--5332
		x"6b",	--5333
		x"5a",	--5334
		x"6b",	--5335
		x"5a",	--5336
		x"6b",	--5337
		x"48",	--5338
		x"49",	--5339
		x"5a",	--5340
		x"6b",	--5341
		x"4d",	--5342
		x"01",	--5343
		x"4e",	--5344
		x"01",	--5345
		x"41",	--5346
		x"01",	--5347
		x"41",	--5348
		x"01",	--5349
		x"81",	--5350
		x"01",	--5351
		x"71",	--5352
		x"01",	--5353
		x"48",	--5354
		x"01",	--5355
		x"49",	--5356
		x"01",	--5357
		x"41",	--5358
		x"01",	--5359
		x"41",	--5360
		x"01",	--5361
		x"51",	--5362
		x"01",	--5363
		x"61",	--5364
		x"01",	--5365
		x"43",	--5366
		x"43",	--5367
		x"43",	--5368
		x"3c",	--5369
		x"41",	--5370
		x"01",	--5371
		x"41",	--5372
		x"01",	--5373
		x"56",	--5374
		x"67",	--5375
		x"93",	--5376
		x"38",	--5377
		x"41",	--5378
		x"01",	--5379
		x"5f",	--5380
		x"5f",	--5381
		x"51",	--5382
		x"01",	--5383
		x"59",	--5384
		x"4f",	--5385
		x"4f",	--5386
		x"00",	--5387
		x"12",	--5388
		x"c2",	--5389
		x"3c",	--5390
		x"43",	--5391
		x"43",	--5392
		x"40",	--5393
		x"00",	--5394
		x"51",	--5395
		x"59",	--5396
		x"4e",	--5397
		x"00",	--5398
		x"4f",	--5399
		x"00",	--5400
		x"53",	--5401
		x"63",	--5402
		x"52",	--5403
		x"97",	--5404
		x"38",	--5405
		x"95",	--5406
		x"3b",	--5407
		x"96",	--5408
		x"2f",	--5409
		x"43",	--5410
		x"01",	--5411
		x"43",	--5412
		x"01",	--5413
		x"41",	--5414
		x"3c",	--5415
		x"41",	--5416
		x"01",	--5417
		x"53",	--5418
		x"5f",	--5419
		x"5f",	--5420
		x"50",	--5421
		x"00",	--5422
		x"54",	--5423
		x"55",	--5424
		x"4f",	--5425
		x"4f",	--5426
		x"00",	--5427
		x"47",	--5428
		x"47",	--5429
		x"12",	--5430
		x"bd",	--5431
		x"4e",	--5432
		x"4f",	--5433
		x"4a",	--5434
		x"4b",	--5435
		x"12",	--5436
		x"bd",	--5437
		x"4e",	--5438
		x"4f",	--5439
		x"53",	--5440
		x"63",	--5441
		x"82",	--5442
		x"99",	--5443
		x"01",	--5444
		x"38",	--5445
		x"91",	--5446
		x"01",	--5447
		x"3b",	--5448
		x"98",	--5449
		x"01",	--5450
		x"2f",	--5451
		x"4a",	--5452
		x"00",	--5453
		x"4b",	--5454
		x"00",	--5455
		x"53",	--5456
		x"01",	--5457
		x"63",	--5458
		x"01",	--5459
		x"52",	--5460
		x"91",	--5461
		x"01",	--5462
		x"01",	--5463
		x"38",	--5464
		x"91",	--5465
		x"01",	--5466
		x"01",	--5467
		x"38",	--5468
		x"91",	--5469
		x"01",	--5470
		x"01",	--5471
		x"2c",	--5472
		x"41",	--5473
		x"01",	--5474
		x"01",	--5475
		x"41",	--5476
		x"01",	--5477
		x"01",	--5478
		x"41",	--5479
		x"01",	--5480
		x"41",	--5481
		x"01",	--5482
		x"53",	--5483
		x"63",	--5484
		x"49",	--5485
		x"01",	--5486
		x"4a",	--5487
		x"01",	--5488
		x"3c",	--5489
		x"41",	--5490
		x"01",	--5491
		x"43",	--5492
		x"43",	--5493
		x"43",	--5494
		x"43",	--5495
		x"43",	--5496
		x"3f",	--5497
		x"41",	--5498
		x"01",	--5499
		x"5f",	--5500
		x"5f",	--5501
		x"51",	--5502
		x"4f",	--5503
		x"4f",	--5504
		x"00",	--5505
		x"41",	--5506
		x"50",	--5507
		x"00",	--5508
		x"4a",	--5509
		x"01",	--5510
		x"41",	--5511
		x"01",	--5512
		x"41",	--5513
		x"01",	--5514
		x"43",	--5515
		x"01",	--5516
		x"46",	--5517
		x"47",	--5518
		x"53",	--5519
		x"63",	--5520
		x"44",	--5521
		x"01",	--5522
		x"45",	--5523
		x"01",	--5524
		x"4a",	--5525
		x"3c",	--5526
		x"43",	--5527
		x"40",	--5528
		x"3b",	--5529
		x"48",	--5530
		x"49",	--5531
		x"12",	--5532
		x"bd",	--5533
		x"12",	--5534
		x"c3",	--5535
		x"12",	--5536
		x"c2",	--5537
		x"4e",	--5538
		x"4f",	--5539
		x"43",	--5540
		x"40",	--5541
		x"43",	--5542
		x"12",	--5543
		x"bd",	--5544
		x"4e",	--5545
		x"4f",	--5546
		x"48",	--5547
		x"49",	--5548
		x"12",	--5549
		x"bd",	--5550
		x"12",	--5551
		x"c3",	--5552
		x"4e",	--5553
		x"00",	--5554
		x"4f",	--5555
		x"00",	--5556
		x"41",	--5557
		x"01",	--5558
		x"5f",	--5559
		x"5f",	--5560
		x"51",	--5561
		x"51",	--5562
		x"01",	--5563
		x"4f",	--5564
		x"00",	--5565
		x"4f",	--5566
		x"00",	--5567
		x"4a",	--5568
		x"4b",	--5569
		x"12",	--5570
		x"bd",	--5571
		x"4e",	--5572
		x"4f",	--5573
		x"53",	--5574
		x"63",	--5575
		x"52",	--5576
		x"82",	--5577
		x"01",	--5578
		x"93",	--5579
		x"38",	--5580
		x"93",	--5581
		x"37",	--5582
		x"93",	--5583
		x"2f",	--5584
		x"41",	--5585
		x"01",	--5586
		x"01",	--5587
		x"41",	--5588
		x"01",	--5589
		x"48",	--5590
		x"49",	--5591
		x"12",	--5592
		x"b7",	--5593
		x"4e",	--5594
		x"4f",	--5595
		x"43",	--5596
		x"40",	--5597
		x"3e",	--5598
		x"12",	--5599
		x"bd",	--5600
		x"12",	--5601
		x"b9",	--5602
		x"43",	--5603
		x"40",	--5604
		x"41",	--5605
		x"12",	--5606
		x"bd",	--5607
		x"4e",	--5608
		x"4f",	--5609
		x"4a",	--5610
		x"4b",	--5611
		x"12",	--5612
		x"bd",	--5613
		x"4e",	--5614
		x"4f",	--5615
		x"12",	--5616
		x"c3",	--5617
		x"4e",	--5618
		x"01",	--5619
		x"4f",	--5620
		x"01",	--5621
		x"12",	--5622
		x"c2",	--5623
		x"4e",	--5624
		x"4f",	--5625
		x"4a",	--5626
		x"4b",	--5627
		x"12",	--5628
		x"bd",	--5629
		x"4e",	--5630
		x"01",	--5631
		x"4f",	--5632
		x"01",	--5633
		x"93",	--5634
		x"01",	--5635
		x"38",	--5636
		x"20",	--5637
		x"93",	--5638
		x"01",	--5639
		x"28",	--5640
		x"41",	--5641
		x"01",	--5642
		x"41",	--5643
		x"01",	--5644
		x"53",	--5645
		x"63",	--5646
		x"4c",	--5647
		x"5b",	--5648
		x"5b",	--5649
		x"51",	--5650
		x"4b",	--5651
		x"00",	--5652
		x"4b",	--5653
		x"00",	--5654
		x"41",	--5655
		x"01",	--5656
		x"42",	--5657
		x"8e",	--5658
		x"46",	--5659
		x"47",	--5660
		x"49",	--5661
		x"f0",	--5662
		x"00",	--5663
		x"93",	--5664
		x"24",	--5665
		x"11",	--5666
		x"10",	--5667
		x"53",	--5668
		x"3f",	--5669
		x"5a",	--5670
		x"01",	--5671
		x"6b",	--5672
		x"01",	--5673
		x"f0",	--5674
		x"00",	--5675
		x"93",	--5676
		x"24",	--5677
		x"5a",	--5678
		x"6b",	--5679
		x"53",	--5680
		x"3f",	--5681
		x"46",	--5682
		x"47",	--5683
		x"8a",	--5684
		x"7b",	--5685
		x"4c",	--5686
		x"5f",	--5687
		x"5f",	--5688
		x"51",	--5689
		x"48",	--5690
		x"00",	--5691
		x"49",	--5692
		x"00",	--5693
		x"48",	--5694
		x"49",	--5695
		x"40",	--5696
		x"00",	--5697
		x"8e",	--5698
		x"f0",	--5699
		x"00",	--5700
		x"93",	--5701
		x"24",	--5702
		x"11",	--5703
		x"10",	--5704
		x"53",	--5705
		x"3f",	--5706
		x"93",	--5707
		x"01",	--5708
		x"20",	--5709
		x"93",	--5710
		x"01",	--5711
		x"20",	--5712
		x"41",	--5713
		x"01",	--5714
		x"53",	--5715
		x"5f",	--5716
		x"5f",	--5717
		x"51",	--5718
		x"4f",	--5719
		x"00",	--5720
		x"4f",	--5721
		x"00",	--5722
		x"10",	--5723
		x"10",	--5724
		x"e7",	--5725
		x"e7",	--5726
		x"11",	--5727
		x"3c",	--5728
		x"43",	--5729
		x"40",	--5730
		x"3f",	--5731
		x"41",	--5732
		x"01",	--5733
		x"41",	--5734
		x"01",	--5735
		x"12",	--5736
		x"c1",	--5737
		x"93",	--5738
		x"34",	--5739
		x"43",	--5740
		x"43",	--5741
		x"3c",	--5742
		x"93",	--5743
		x"38",	--5744
		x"20",	--5745
		x"93",	--5746
		x"28",	--5747
		x"3c",	--5748
		x"43",	--5749
		x"43",	--5750
		x"53",	--5751
		x"01",	--5752
		x"63",	--5753
		x"01",	--5754
		x"43",	--5755
		x"43",	--5756
		x"43",	--5757
		x"43",	--5758
		x"41",	--5759
		x"01",	--5760
		x"3c",	--5761
		x"4b",	--5762
		x"4b",	--5763
		x"00",	--5764
		x"93",	--5765
		x"20",	--5766
		x"93",	--5767
		x"20",	--5768
		x"93",	--5769
		x"20",	--5770
		x"93",	--5771
		x"24",	--5772
		x"40",	--5773
		x"01",	--5774
		x"43",	--5775
		x"4e",	--5776
		x"4f",	--5777
		x"8c",	--5778
		x"7d",	--5779
		x"49",	--5780
		x"00",	--5781
		x"4a",	--5782
		x"00",	--5783
		x"3c",	--5784
		x"40",	--5785
		x"00",	--5786
		x"43",	--5787
		x"4e",	--5788
		x"4f",	--5789
		x"8c",	--5790
		x"7d",	--5791
		x"48",	--5792
		x"00",	--5793
		x"49",	--5794
		x"00",	--5795
		x"43",	--5796
		x"43",	--5797
		x"53",	--5798
		x"63",	--5799
		x"52",	--5800
		x"91",	--5801
		x"01",	--5802
		x"3b",	--5803
		x"20",	--5804
		x"91",	--5805
		x"01",	--5806
		x"2b",	--5807
		x"93",	--5808
		x"01",	--5809
		x"38",	--5810
		x"20",	--5811
		x"93",	--5812
		x"01",	--5813
		x"28",	--5814
		x"93",	--5815
		x"01",	--5816
		x"20",	--5817
		x"93",	--5818
		x"01",	--5819
		x"24",	--5820
		x"93",	--5821
		x"01",	--5822
		x"20",	--5823
		x"93",	--5824
		x"01",	--5825
		x"24",	--5826
		x"3c",	--5827
		x"41",	--5828
		x"01",	--5829
		x"53",	--5830
		x"5f",	--5831
		x"5f",	--5832
		x"51",	--5833
		x"f0",	--5834
		x"00",	--5835
		x"00",	--5836
		x"f3",	--5837
		x"00",	--5838
		x"3c",	--5839
		x"41",	--5840
		x"01",	--5841
		x"53",	--5842
		x"5f",	--5843
		x"5f",	--5844
		x"51",	--5845
		x"f0",	--5846
		x"00",	--5847
		x"00",	--5848
		x"f3",	--5849
		x"00",	--5850
		x"93",	--5851
		x"20",	--5852
		x"93",	--5853
		x"20",	--5854
		x"41",	--5855
		x"01",	--5856
		x"41",	--5857
		x"01",	--5858
		x"43",	--5859
		x"40",	--5860
		x"3f",	--5861
		x"12",	--5862
		x"bd",	--5863
		x"4e",	--5864
		x"01",	--5865
		x"4f",	--5866
		x"01",	--5867
		x"93",	--5868
		x"20",	--5869
		x"93",	--5870
		x"24",	--5871
		x"41",	--5872
		x"01",	--5873
		x"43",	--5874
		x"40",	--5875
		x"3f",	--5876
		x"12",	--5877
		x"b7",	--5878
		x"4e",	--5879
		x"4f",	--5880
		x"41",	--5881
		x"01",	--5882
		x"41",	--5883
		x"01",	--5884
		x"12",	--5885
		x"bd",	--5886
		x"4e",	--5887
		x"01",	--5888
		x"4f",	--5889
		x"01",	--5890
		x"43",	--5891
		x"43",	--5892
		x"41",	--5893
		x"01",	--5894
		x"41",	--5895
		x"01",	--5896
		x"12",	--5897
		x"c1",	--5898
		x"93",	--5899
		x"20",	--5900
		x"41",	--5901
		x"01",	--5902
		x"41",	--5903
		x"01",	--5904
		x"53",	--5905
		x"63",	--5906
		x"41",	--5907
		x"01",	--5908
		x"41",	--5909
		x"01",	--5910
		x"43",	--5911
		x"43",	--5912
		x"01",	--5913
		x"43",	--5914
		x"01",	--5915
		x"3c",	--5916
		x"4a",	--5917
		x"5f",	--5918
		x"5f",	--5919
		x"40",	--5920
		x"00",	--5921
		x"51",	--5922
		x"5e",	--5923
		x"59",	--5924
		x"df",	--5925
		x"00",	--5926
		x"01",	--5927
		x"df",	--5928
		x"00",	--5929
		x"01",	--5930
		x"53",	--5931
		x"63",	--5932
		x"82",	--5933
		x"91",	--5934
		x"01",	--5935
		x"38",	--5936
		x"9d",	--5937
		x"01",	--5938
		x"3b",	--5939
		x"91",	--5940
		x"01",	--5941
		x"2f",	--5942
		x"93",	--5943
		x"01",	--5944
		x"20",	--5945
		x"93",	--5946
		x"01",	--5947
		x"24",	--5948
		x"3c",	--5949
		x"53",	--5950
		x"01",	--5951
		x"63",	--5952
		x"01",	--5953
		x"3c",	--5954
		x"43",	--5955
		x"43",	--5956
		x"01",	--5957
		x"43",	--5958
		x"01",	--5959
		x"82",	--5960
		x"41",	--5961
		x"01",	--5962
		x"5f",	--5963
		x"5f",	--5964
		x"40",	--5965
		x"00",	--5966
		x"51",	--5967
		x"58",	--5968
		x"5e",	--5969
		x"93",	--5970
		x"00",	--5971
		x"20",	--5972
		x"93",	--5973
		x"00",	--5974
		x"27",	--5975
		x"41",	--5976
		x"01",	--5977
		x"41",	--5978
		x"01",	--5979
		x"53",	--5980
		x"63",	--5981
		x"49",	--5982
		x"01",	--5983
		x"4a",	--5984
		x"01",	--5985
		x"43",	--5986
		x"01",	--5987
		x"43",	--5988
		x"49",	--5989
		x"01",	--5990
		x"41",	--5991
		x"01",	--5992
		x"41",	--5993
		x"01",	--5994
		x"59",	--5995
		x"6a",	--5996
		x"4d",	--5997
		x"01",	--5998
		x"4e",	--5999
		x"01",	--6000
		x"49",	--6001
		x"51",	--6002
		x"01",	--6003
		x"48",	--6004
		x"01",	--6005
		x"44",	--6006
		x"3c",	--6007
		x"52",	--6008
		x"01",	--6009
		x"41",	--6010
		x"01",	--6011
		x"5f",	--6012
		x"5f",	--6013
		x"41",	--6014
		x"50",	--6015
		x"00",	--6016
		x"5f",	--6017
		x"41",	--6018
		x"01",	--6019
		x"54",	--6020
		x"41",	--6021
		x"01",	--6022
		x"5f",	--6023
		x"5f",	--6024
		x"51",	--6025
		x"01",	--6026
		x"56",	--6027
		x"4f",	--6028
		x"4f",	--6029
		x"00",	--6030
		x"12",	--6031
		x"c2",	--6032
		x"4e",	--6033
		x"ff",	--6034
		x"4f",	--6035
		x"ff",	--6036
		x"41",	--6037
		x"01",	--6038
		x"41",	--6039
		x"01",	--6040
		x"41",	--6041
		x"01",	--6042
		x"43",	--6043
		x"43",	--6044
		x"43",	--6045
		x"56",	--6046
		x"3c",	--6047
		x"44",	--6048
		x"55",	--6049
		x"4f",	--6050
		x"4f",	--6051
		x"00",	--6052
		x"47",	--6053
		x"47",	--6054
		x"12",	--6055
		x"bd",	--6056
		x"4e",	--6057
		x"4f",	--6058
		x"48",	--6059
		x"49",	--6060
		x"12",	--6061
		x"bd",	--6062
		x"4e",	--6063
		x"4f",	--6064
		x"53",	--6065
		x"63",	--6066
		x"82",	--6067
		x"9b",	--6068
		x"01",	--6069
		x"38",	--6070
		x"91",	--6071
		x"01",	--6072
		x"3b",	--6073
		x"9a",	--6074
		x"01",	--6075
		x"2f",	--6076
		x"41",	--6077
		x"01",	--6078
		x"5f",	--6079
		x"5f",	--6080
		x"51",	--6081
		x"51",	--6082
		x"01",	--6083
		x"48",	--6084
		x"ff",	--6085
		x"49",	--6086
		x"ff",	--6087
		x"53",	--6088
		x"01",	--6089
		x"63",	--6090
		x"01",	--6091
		x"52",	--6092
		x"41",	--6093
		x"01",	--6094
		x"41",	--6095
		x"01",	--6096
		x"51",	--6097
		x"01",	--6098
		x"61",	--6099
		x"01",	--6100
		x"91",	--6101
		x"01",	--6102
		x"38",	--6103
		x"9f",	--6104
		x"01",	--6105
		x"3b",	--6106
		x"91",	--6107
		x"01",	--6108
		x"2f",	--6109
		x"4e",	--6110
		x"01",	--6111
		x"4f",	--6112
		x"01",	--6113
		x"40",	--6114
		x"aa",	--6115
		x"46",	--6116
		x"01",	--6117
		x"47",	--6118
		x"01",	--6119
		x"41",	--6120
		x"01",	--6121
		x"e3",	--6122
		x"47",	--6123
		x"53",	--6124
		x"41",	--6125
		x"01",	--6126
		x"41",	--6127
		x"01",	--6128
		x"12",	--6129
		x"b7",	--6130
		x"4e",	--6131
		x"4f",	--6132
		x"43",	--6133
		x"40",	--6134
		x"43",	--6135
		x"12",	--6136
		x"c1",	--6137
		x"93",	--6138
		x"34",	--6139
		x"3c",	--6140
		x"46",	--6141
		x"01",	--6142
		x"47",	--6143
		x"01",	--6144
		x"41",	--6145
		x"01",	--6146
		x"41",	--6147
		x"01",	--6148
		x"53",	--6149
		x"63",	--6150
		x"82",	--6151
		x"01",	--6152
		x"73",	--6153
		x"01",	--6154
		x"46",	--6155
		x"01",	--6156
		x"47",	--6157
		x"01",	--6158
		x"43",	--6159
		x"3c",	--6160
		x"53",	--6161
		x"01",	--6162
		x"63",	--6163
		x"01",	--6164
		x"82",	--6165
		x"01",	--6166
		x"73",	--6167
		x"01",	--6168
		x"82",	--6169
		x"46",	--6170
		x"5f",	--6171
		x"5f",	--6172
		x"40",	--6173
		x"00",	--6174
		x"51",	--6175
		x"59",	--6176
		x"5d",	--6177
		x"93",	--6178
		x"00",	--6179
		x"20",	--6180
		x"93",	--6181
		x"00",	--6182
		x"27",	--6183
		x"3c",	--6184
		x"43",	--6185
		x"40",	--6186
		x"3b",	--6187
		x"46",	--6188
		x"47",	--6189
		x"12",	--6190
		x"bd",	--6191
		x"12",	--6192
		x"c3",	--6193
		x"12",	--6194
		x"c2",	--6195
		x"4e",	--6196
		x"4f",	--6197
		x"41",	--6198
		x"01",	--6199
		x"5c",	--6200
		x"5c",	--6201
		x"41",	--6202
		x"5c",	--6203
		x"50",	--6204
		x"00",	--6205
		x"43",	--6206
		x"40",	--6207
		x"43",	--6208
		x"12",	--6209
		x"bd",	--6210
		x"4e",	--6211
		x"4f",	--6212
		x"46",	--6213
		x"47",	--6214
		x"12",	--6215
		x"bd",	--6216
		x"12",	--6217
		x"c3",	--6218
		x"4e",	--6219
		x"00",	--6220
		x"4f",	--6221
		x"00",	--6222
		x"53",	--6223
		x"01",	--6224
		x"63",	--6225
		x"01",	--6226
		x"52",	--6227
		x"01",	--6228
		x"63",	--6229
		x"01",	--6230
		x"41",	--6231
		x"01",	--6232
		x"5c",	--6233
		x"5c",	--6234
		x"41",	--6235
		x"5c",	--6236
		x"50",	--6237
		x"00",	--6238
		x"44",	--6239
		x"45",	--6240
		x"12",	--6241
		x"c3",	--6242
		x"4e",	--6243
		x"00",	--6244
		x"4f",	--6245
		x"00",	--6246
		x"3c",	--6247
		x"41",	--6248
		x"01",	--6249
		x"5c",	--6250
		x"5c",	--6251
		x"41",	--6252
		x"5c",	--6253
		x"50",	--6254
		x"00",	--6255
		x"46",	--6256
		x"47",	--6257
		x"12",	--6258
		x"c3",	--6259
		x"4e",	--6260
		x"00",	--6261
		x"4f",	--6262
		x"00",	--6263
		x"41",	--6264
		x"01",	--6265
		x"43",	--6266
		x"40",	--6267
		x"3f",	--6268
		x"12",	--6269
		x"b7",	--6270
		x"4e",	--6271
		x"4f",	--6272
		x"41",	--6273
		x"01",	--6274
		x"41",	--6275
		x"01",	--6276
		x"43",	--6277
		x"93",	--6278
		x"38",	--6279
		x"41",	--6280
		x"01",	--6281
		x"5f",	--6282
		x"5f",	--6283
		x"41",	--6284
		x"5f",	--6285
		x"5b",	--6286
		x"40",	--6287
		x"00",	--6288
		x"51",	--6289
		x"5d",	--6290
		x"5b",	--6291
		x"4f",	--6292
		x"4f",	--6293
		x"00",	--6294
		x"12",	--6295
		x"c2",	--6296
		x"4e",	--6297
		x"4f",	--6298
		x"46",	--6299
		x"47",	--6300
		x"12",	--6301
		x"bd",	--6302
		x"4e",	--6303
		x"00",	--6304
		x"4f",	--6305
		x"00",	--6306
		x"43",	--6307
		x"40",	--6308
		x"3b",	--6309
		x"46",	--6310
		x"47",	--6311
		x"12",	--6312
		x"bd",	--6313
		x"4e",	--6314
		x"4f",	--6315
		x"53",	--6316
		x"63",	--6317
		x"82",	--6318
		x"3f",	--6319
		x"41",	--6320
		x"01",	--6321
		x"01",	--6322
		x"41",	--6323
		x"01",	--6324
		x"01",	--6325
		x"43",	--6326
		x"43",	--6327
		x"43",	--6328
		x"3c",	--6329
		x"41",	--6330
		x"01",	--6331
		x"5f",	--6332
		x"5f",	--6333
		x"51",	--6334
		x"87",	--6335
		x"56",	--6336
		x"4f",	--6337
		x"4f",	--6338
		x"00",	--6339
		x"46",	--6340
		x"db",	--6341
		x"46",	--6342
		x"db",	--6343
		x"12",	--6344
		x"bd",	--6345
		x"4e",	--6346
		x"4f",	--6347
		x"48",	--6348
		x"49",	--6349
		x"12",	--6350
		x"bd",	--6351
		x"4e",	--6352
		x"4f",	--6353
		x"53",	--6354
		x"63",	--6355
		x"52",	--6356
		x"9b",	--6357
		x"01",	--6358
		x"38",	--6359
		x"20",	--6360
		x"9a",	--6361
		x"01",	--6362
		x"28",	--6363
		x"9b",	--6364
		x"38",	--6365
		x"95",	--6366
		x"3b",	--6367
		x"9a",	--6368
		x"2f",	--6369
		x"40",	--6370
		x"00",	--6371
		x"51",	--6372
		x"57",	--6373
		x"48",	--6374
		x"00",	--6375
		x"49",	--6376
		x"00",	--6377
		x"53",	--6378
		x"01",	--6379
		x"63",	--6380
		x"01",	--6381
		x"52",	--6382
		x"53",	--6383
		x"63",	--6384
		x"93",	--6385
		x"01",	--6386
		x"38",	--6387
		x"43",	--6388
		x"43",	--6389
		x"43",	--6390
		x"43",	--6391
		x"43",	--6392
		x"3f",	--6393
		x"90",	--6394
		x"00",	--6395
		x"01",	--6396
		x"34",	--6397
		x"93",	--6398
		x"01",	--6399
		x"34",	--6400
		x"93",	--6401
		x"01",	--6402
		x"24",	--6403
		x"40",	--6404
		x"b5",	--6405
		x"90",	--6406
		x"00",	--6407
		x"01",	--6408
		x"24",	--6409
		x"40",	--6410
		x"b5",	--6411
		x"3c",	--6412
		x"41",	--6413
		x"01",	--6414
		x"41",	--6415
		x"01",	--6416
		x"43",	--6417
		x"43",	--6418
		x"43",	--6419
		x"93",	--6420
		x"38",	--6421
		x"41",	--6422
		x"01",	--6423
		x"5f",	--6424
		x"5f",	--6425
		x"40",	--6426
		x"00",	--6427
		x"51",	--6428
		x"5e",	--6429
		x"55",	--6430
		x"4f",	--6431
		x"4f",	--6432
		x"00",	--6433
		x"4a",	--6434
		x"4b",	--6435
		x"12",	--6436
		x"bd",	--6437
		x"4e",	--6438
		x"4f",	--6439
		x"53",	--6440
		x"63",	--6441
		x"82",	--6442
		x"3f",	--6443
		x"93",	--6444
		x"01",	--6445
		x"20",	--6446
		x"93",	--6447
		x"01",	--6448
		x"24",	--6449
		x"e0",	--6450
		x"80",	--6451
		x"41",	--6452
		x"01",	--6453
		x"4a",	--6454
		x"00",	--6455
		x"4b",	--6456
		x"00",	--6457
		x"40",	--6458
		x"b5",	--6459
		x"41",	--6460
		x"01",	--6461
		x"41",	--6462
		x"01",	--6463
		x"43",	--6464
		x"43",	--6465
		x"43",	--6466
		x"93",	--6467
		x"38",	--6468
		x"41",	--6469
		x"01",	--6470
		x"5f",	--6471
		x"5f",	--6472
		x"40",	--6473
		x"00",	--6474
		x"51",	--6475
		x"59",	--6476
		x"55",	--6477
		x"4f",	--6478
		x"4f",	--6479
		x"00",	--6480
		x"4a",	--6481
		x"4b",	--6482
		x"12",	--6483
		x"bd",	--6484
		x"4e",	--6485
		x"4f",	--6486
		x"53",	--6487
		x"63",	--6488
		x"82",	--6489
		x"3f",	--6490
		x"4a",	--6491
		x"4b",	--6492
		x"93",	--6493
		x"01",	--6494
		x"20",	--6495
		x"93",	--6496
		x"01",	--6497
		x"24",	--6498
		x"e0",	--6499
		x"80",	--6500
		x"41",	--6501
		x"01",	--6502
		x"4a",	--6503
		x"00",	--6504
		x"4b",	--6505
		x"00",	--6506
		x"41",	--6507
		x"00",	--6508
		x"41",	--6509
		x"00",	--6510
		x"12",	--6511
		x"bd",	--6512
		x"41",	--6513
		x"50",	--6514
		x"00",	--6515
		x"43",	--6516
		x"43",	--6517
		x"3c",	--6518
		x"45",	--6519
		x"45",	--6520
		x"12",	--6521
		x"bd",	--6522
		x"53",	--6523
		x"63",	--6524
		x"97",	--6525
		x"01",	--6526
		x"38",	--6527
		x"91",	--6528
		x"01",	--6529
		x"3b",	--6530
		x"96",	--6531
		x"01",	--6532
		x"2f",	--6533
		x"4e",	--6534
		x"4f",	--6535
		x"93",	--6536
		x"01",	--6537
		x"20",	--6538
		x"93",	--6539
		x"01",	--6540
		x"24",	--6541
		x"e0",	--6542
		x"80",	--6543
		x"41",	--6544
		x"01",	--6545
		x"4a",	--6546
		x"00",	--6547
		x"4b",	--6548
		x"00",	--6549
		x"40",	--6550
		x"b5",	--6551
		x"41",	--6552
		x"01",	--6553
		x"5f",	--6554
		x"5f",	--6555
		x"40",	--6556
		x"00",	--6557
		x"51",	--6558
		x"5f",	--6559
		x"51",	--6560
		x"01",	--6561
		x"4a",	--6562
		x"01",	--6563
		x"4a",	--6564
		x"00",	--6565
		x"4a",	--6566
		x"00",	--6567
		x"41",	--6568
		x"01",	--6569
		x"5f",	--6570
		x"5f",	--6571
		x"40",	--6572
		x"00",	--6573
		x"51",	--6574
		x"5f",	--6575
		x"51",	--6576
		x"01",	--6577
		x"49",	--6578
		x"01",	--6579
		x"49",	--6580
		x"49",	--6581
		x"00",	--6582
		x"48",	--6583
		x"49",	--6584
		x"46",	--6585
		x"47",	--6586
		x"12",	--6587
		x"bd",	--6588
		x"4e",	--6589
		x"4f",	--6590
		x"4e",	--6591
		x"4f",	--6592
		x"46",	--6593
		x"47",	--6594
		x"12",	--6595
		x"bd",	--6596
		x"4e",	--6597
		x"4f",	--6598
		x"48",	--6599
		x"49",	--6600
		x"12",	--6601
		x"bd",	--6602
		x"41",	--6603
		x"01",	--6604
		x"4e",	--6605
		x"00",	--6606
		x"4f",	--6607
		x"00",	--6608
		x"41",	--6609
		x"01",	--6610
		x"4a",	--6611
		x"00",	--6612
		x"4b",	--6613
		x"00",	--6614
		x"53",	--6615
		x"63",	--6616
		x"82",	--6617
		x"01",	--6618
		x"3c",	--6619
		x"41",	--6620
		x"01",	--6621
		x"41",	--6622
		x"01",	--6623
		x"43",	--6624
		x"01",	--6625
		x"43",	--6626
		x"01",	--6627
		x"4c",	--6628
		x"4d",	--6629
		x"53",	--6630
		x"63",	--6631
		x"48",	--6632
		x"01",	--6633
		x"49",	--6634
		x"01",	--6635
		x"4c",	--6636
		x"4d",	--6637
		x"82",	--6638
		x"01",	--6639
		x"93",	--6640
		x"38",	--6641
		x"93",	--6642
		x"37",	--6643
		x"93",	--6644
		x"2f",	--6645
		x"41",	--6646
		x"01",	--6647
		x"41",	--6648
		x"01",	--6649
		x"43",	--6650
		x"01",	--6651
		x"43",	--6652
		x"01",	--6653
		x"4c",	--6654
		x"4d",	--6655
		x"53",	--6656
		x"63",	--6657
		x"49",	--6658
		x"01",	--6659
		x"4a",	--6660
		x"01",	--6661
		x"4c",	--6662
		x"4d",	--6663
		x"3c",	--6664
		x"41",	--6665
		x"01",	--6666
		x"5f",	--6667
		x"5f",	--6668
		x"40",	--6669
		x"00",	--6670
		x"51",	--6671
		x"5f",	--6672
		x"51",	--6673
		x"01",	--6674
		x"4a",	--6675
		x"01",	--6676
		x"4a",	--6677
		x"00",	--6678
		x"4a",	--6679
		x"00",	--6680
		x"41",	--6681
		x"01",	--6682
		x"5f",	--6683
		x"5f",	--6684
		x"40",	--6685
		x"00",	--6686
		x"51",	--6687
		x"5f",	--6688
		x"51",	--6689
		x"01",	--6690
		x"49",	--6691
		x"01",	--6692
		x"49",	--6693
		x"49",	--6694
		x"00",	--6695
		x"48",	--6696
		x"49",	--6697
		x"46",	--6698
		x"47",	--6699
		x"12",	--6700
		x"bd",	--6701
		x"4e",	--6702
		x"4f",	--6703
		x"4e",	--6704
		x"4f",	--6705
		x"46",	--6706
		x"47",	--6707
		x"12",	--6708
		x"bd",	--6709
		x"4e",	--6710
		x"4f",	--6711
		x"48",	--6712
		x"49",	--6713
		x"12",	--6714
		x"bd",	--6715
		x"41",	--6716
		x"01",	--6717
		x"4e",	--6718
		x"00",	--6719
		x"4f",	--6720
		x"00",	--6721
		x"41",	--6722
		x"01",	--6723
		x"4a",	--6724
		x"00",	--6725
		x"4b",	--6726
		x"00",	--6727
		x"53",	--6728
		x"63",	--6729
		x"82",	--6730
		x"01",	--6731
		x"82",	--6732
		x"01",	--6733
		x"93",	--6734
		x"38",	--6735
		x"93",	--6736
		x"37",	--6737
		x"93",	--6738
		x"2f",	--6739
		x"41",	--6740
		x"01",	--6741
		x"41",	--6742
		x"01",	--6743
		x"43",	--6744
		x"43",	--6745
		x"43",	--6746
		x"3c",	--6747
		x"41",	--6748
		x"01",	--6749
		x"5f",	--6750
		x"5f",	--6751
		x"40",	--6752
		x"00",	--6753
		x"51",	--6754
		x"5d",	--6755
		x"55",	--6756
		x"4f",	--6757
		x"4f",	--6758
		x"00",	--6759
		x"4a",	--6760
		x"4b",	--6761
		x"12",	--6762
		x"bd",	--6763
		x"4e",	--6764
		x"4f",	--6765
		x"53",	--6766
		x"63",	--6767
		x"82",	--6768
		x"93",	--6769
		x"38",	--6770
		x"93",	--6771
		x"37",	--6772
		x"93",	--6773
		x"2f",	--6774
		x"93",	--6775
		x"01",	--6776
		x"20",	--6777
		x"93",	--6778
		x"01",	--6779
		x"20",	--6780
		x"41",	--6781
		x"01",	--6782
		x"41",	--6783
		x"00",	--6784
		x"00",	--6785
		x"41",	--6786
		x"00",	--6787
		x"00",	--6788
		x"41",	--6789
		x"00",	--6790
		x"00",	--6791
		x"41",	--6792
		x"00",	--6793
		x"00",	--6794
		x"4a",	--6795
		x"00",	--6796
		x"4b",	--6797
		x"00",	--6798
		x"3c",	--6799
		x"41",	--6800
		x"00",	--6801
		x"41",	--6802
		x"00",	--6803
		x"e0",	--6804
		x"80",	--6805
		x"41",	--6806
		x"01",	--6807
		x"4d",	--6808
		x"00",	--6809
		x"4e",	--6810
		x"00",	--6811
		x"41",	--6812
		x"00",	--6813
		x"41",	--6814
		x"00",	--6815
		x"e0",	--6816
		x"80",	--6817
		x"4d",	--6818
		x"00",	--6819
		x"4e",	--6820
		x"00",	--6821
		x"4a",	--6822
		x"4b",	--6823
		x"e0",	--6824
		x"80",	--6825
		x"4d",	--6826
		x"00",	--6827
		x"4e",	--6828
		x"00",	--6829
		x"41",	--6830
		x"01",	--6831
		x"f0",	--6832
		x"00",	--6833
		x"50",	--6834
		x"01",	--6835
		x"41",	--6836
		x"41",	--6837
		x"41",	--6838
		x"41",	--6839
		x"41",	--6840
		x"41",	--6841
		x"41",	--6842
		x"41",	--6843
		x"41",	--6844
		x"12",	--6845
		x"12",	--6846
		x"82",	--6847
		x"4e",	--6848
		x"4f",	--6849
		x"f3",	--6850
		x"f0",	--6851
		x"7f",	--6852
		x"90",	--6853
		x"3f",	--6854
		x"38",	--6855
		x"90",	--6856
		x"3f",	--6857
		x"34",	--6858
		x"90",	--6859
		x"0f",	--6860
		x"2c",	--6861
		x"43",	--6862
		x"43",	--6863
		x"3c",	--6864
		x"90",	--6865
		x"7f",	--6866
		x"38",	--6867
		x"4e",	--6868
		x"4f",	--6869
		x"12",	--6870
		x"bd",	--6871
		x"3c",	--6872
		x"41",	--6873
		x"12",	--6874
		x"a3",	--6875
		x"4e",	--6876
		x"4f",	--6877
		x"f0",	--6878
		x"00",	--6879
		x"f3",	--6880
		x"41",	--6881
		x"00",	--6882
		x"41",	--6883
		x"00",	--6884
		x"41",	--6885
		x"41",	--6886
		x"00",	--6887
		x"93",	--6888
		x"20",	--6889
		x"93",	--6890
		x"24",	--6891
		x"93",	--6892
		x"20",	--6893
		x"93",	--6894
		x"24",	--6895
		x"41",	--6896
		x"41",	--6897
		x"00",	--6898
		x"93",	--6899
		x"20",	--6900
		x"93",	--6901
		x"20",	--6902
		x"12",	--6903
		x"a1",	--6904
		x"3c",	--6905
		x"12",	--6906
		x"12",	--6907
		x"b6",	--6908
		x"53",	--6909
		x"3c",	--6910
		x"12",	--6911
		x"a1",	--6912
		x"e0",	--6913
		x"80",	--6914
		x"3c",	--6915
		x"12",	--6916
		x"12",	--6917
		x"b6",	--6918
		x"53",	--6919
		x"52",	--6920
		x"41",	--6921
		x"41",	--6922
		x"41",	--6923
		x"12",	--6924
		x"b5",	--6925
		x"41",	--6926
		x"12",	--6927
		x"12",	--6928
		x"12",	--6929
		x"12",	--6930
		x"12",	--6931
		x"12",	--6932
		x"12",	--6933
		x"12",	--6934
		x"82",	--6935
		x"4e",	--6936
		x"4f",	--6937
		x"4c",	--6938
		x"00",	--6939
		x"4d",	--6940
		x"00",	--6941
		x"4e",	--6942
		x"4f",	--6943
		x"f3",	--6944
		x"f0",	--6945
		x"7f",	--6946
		x"90",	--6947
		x"32",	--6948
		x"34",	--6949
		x"12",	--6950
		x"c3",	--6951
		x"93",	--6952
		x"24",	--6953
		x"48",	--6954
		x"49",	--6955
		x"48",	--6956
		x"49",	--6957
		x"12",	--6958
		x"bd",	--6959
		x"4e",	--6960
		x"4f",	--6961
		x"48",	--6962
		x"49",	--6963
		x"12",	--6964
		x"bd",	--6965
		x"4e",	--6966
		x"4f",	--6967
		x"40",	--6968
		x"c9",	--6969
		x"40",	--6970
		x"2f",	--6971
		x"4a",	--6972
		x"4b",	--6973
		x"12",	--6974
		x"bd",	--6975
		x"40",	--6976
		x"2f",	--6977
		x"40",	--6978
		x"32",	--6979
		x"12",	--6980
		x"bd",	--6981
		x"4e",	--6982
		x"4f",	--6983
		x"4a",	--6984
		x"4b",	--6985
		x"12",	--6986
		x"bd",	--6987
		x"40",	--6988
		x"ef",	--6989
		x"40",	--6990
		x"36",	--6991
		x"12",	--6992
		x"bd",	--6993
		x"4e",	--6994
		x"4f",	--6995
		x"4a",	--6996
		x"4b",	--6997
		x"12",	--6998
		x"bd",	--6999
		x"40",	--7000
		x"0d",	--7001
		x"40",	--7002
		x"39",	--7003
		x"12",	--7004
		x"bd",	--7005
		x"4e",	--7006
		x"4f",	--7007
		x"4a",	--7008
		x"4b",	--7009
		x"12",	--7010
		x"bd",	--7011
		x"40",	--7012
		x"88",	--7013
		x"40",	--7014
		x"3c",	--7015
		x"12",	--7016
		x"bd",	--7017
		x"4e",	--7018
		x"4f",	--7019
		x"93",	--7020
		x"00",	--7021
		x"20",	--7022
		x"4e",	--7023
		x"4f",	--7024
		x"4a",	--7025
		x"4b",	--7026
		x"12",	--7027
		x"bd",	--7028
		x"40",	--7029
		x"aa",	--7030
		x"40",	--7031
		x"3e",	--7032
		x"12",	--7033
		x"bd",	--7034
		x"4e",	--7035
		x"4f",	--7036
		x"46",	--7037
		x"47",	--7038
		x"12",	--7039
		x"bd",	--7040
		x"4e",	--7041
		x"4f",	--7042
		x"48",	--7043
		x"49",	--7044
		x"12",	--7045
		x"bd",	--7046
		x"3c",	--7047
		x"43",	--7048
		x"40",	--7049
		x"3f",	--7050
		x"41",	--7051
		x"41",	--7052
		x"00",	--7053
		x"12",	--7054
		x"bd",	--7055
		x"4e",	--7056
		x"00",	--7057
		x"4f",	--7058
		x"00",	--7059
		x"44",	--7060
		x"45",	--7061
		x"46",	--7062
		x"47",	--7063
		x"12",	--7064
		x"bd",	--7065
		x"4e",	--7066
		x"4f",	--7067
		x"41",	--7068
		x"00",	--7069
		x"41",	--7070
		x"00",	--7071
		x"12",	--7072
		x"bd",	--7073
		x"4e",	--7074
		x"4f",	--7075
		x"4a",	--7076
		x"4b",	--7077
		x"12",	--7078
		x"bd",	--7079
		x"41",	--7080
		x"41",	--7081
		x"00",	--7082
		x"12",	--7083
		x"bd",	--7084
		x"4e",	--7085
		x"4f",	--7086
		x"40",	--7087
		x"aa",	--7088
		x"40",	--7089
		x"3e",	--7090
		x"46",	--7091
		x"47",	--7092
		x"12",	--7093
		x"bd",	--7094
		x"4e",	--7095
		x"4f",	--7096
		x"4a",	--7097
		x"4b",	--7098
		x"12",	--7099
		x"bd",	--7100
		x"4e",	--7101
		x"4f",	--7102
		x"48",	--7103
		x"49",	--7104
		x"12",	--7105
		x"bd",	--7106
		x"4e",	--7107
		x"4f",	--7108
		x"48",	--7109
		x"49",	--7110
		x"52",	--7111
		x"41",	--7112
		x"41",	--7113
		x"41",	--7114
		x"41",	--7115
		x"41",	--7116
		x"41",	--7117
		x"41",	--7118
		x"41",	--7119
		x"41",	--7120
		x"12",	--7121
		x"12",	--7122
		x"12",	--7123
		x"12",	--7124
		x"12",	--7125
		x"4d",	--7126
		x"4e",	--7127
		x"4f",	--7128
		x"48",	--7129
		x"49",	--7130
		x"f3",	--7131
		x"f0",	--7132
		x"7f",	--7133
		x"93",	--7134
		x"20",	--7135
		x"93",	--7136
		x"24",	--7137
		x"90",	--7138
		x"7f",	--7139
		x"28",	--7140
		x"4e",	--7141
		x"4f",	--7142
		x"12",	--7143
		x"bd",	--7144
		x"3c",	--7145
		x"90",	--7146
		x"00",	--7147
		x"28",	--7148
		x"4d",	--7149
		x"43",	--7150
		x"40",	--7151
		x"00",	--7152
		x"c3",	--7153
		x"10",	--7154
		x"10",	--7155
		x"53",	--7156
		x"23",	--7157
		x"3c",	--7158
		x"43",	--7159
		x"40",	--7160
		x"4c",	--7161
		x"12",	--7162
		x"bd",	--7163
		x"4e",	--7164
		x"4f",	--7165
		x"48",	--7166
		x"49",	--7167
		x"f3",	--7168
		x"f0",	--7169
		x"7f",	--7170
		x"4b",	--7171
		x"4b",	--7172
		x"10",	--7173
		x"11",	--7174
		x"10",	--7175
		x"11",	--7176
		x"40",	--7177
		x"00",	--7178
		x"11",	--7179
		x"10",	--7180
		x"53",	--7181
		x"23",	--7182
		x"50",	--7183
		x"ff",	--7184
		x"63",	--7185
		x"47",	--7186
		x"47",	--7187
		x"10",	--7188
		x"11",	--7189
		x"10",	--7190
		x"11",	--7191
		x"4e",	--7192
		x"5a",	--7193
		x"6b",	--7194
		x"93",	--7195
		x"38",	--7196
		x"20",	--7197
		x"90",	--7198
		x"00",	--7199
		x"28",	--7200
		x"40",	--7201
		x"f2",	--7202
		x"40",	--7203
		x"71",	--7204
		x"93",	--7205
		x"34",	--7206
		x"40",	--7207
		x"f2",	--7208
		x"40",	--7209
		x"f1",	--7210
		x"40",	--7211
		x"f2",	--7212
		x"40",	--7213
		x"71",	--7214
		x"4a",	--7215
		x"4b",	--7216
		x"3c",	--7217
		x"93",	--7218
		x"38",	--7219
		x"20",	--7220
		x"93",	--7221
		x"28",	--7222
		x"43",	--7223
		x"43",	--7224
		x"4c",	--7225
		x"40",	--7226
		x"00",	--7227
		x"5a",	--7228
		x"6b",	--7229
		x"53",	--7230
		x"23",	--7231
		x"f3",	--7232
		x"f0",	--7233
		x"80",	--7234
		x"da",	--7235
		x"db",	--7236
		x"48",	--7237
		x"49",	--7238
		x"3c",	--7239
		x"93",	--7240
		x"38",	--7241
		x"93",	--7242
		x"34",	--7243
		x"90",	--7244
		x"ff",	--7245
		x"2c",	--7246
		x"4f",	--7247
		x"f0",	--7248
		x"80",	--7249
		x"90",	--7250
		x"75",	--7251
		x"38",	--7252
		x"40",	--7253
		x"f2",	--7254
		x"40",	--7255
		x"71",	--7256
		x"93",	--7257
		x"24",	--7258
		x"40",	--7259
		x"f2",	--7260
		x"40",	--7261
		x"f1",	--7262
		x"40",	--7263
		x"f2",	--7264
		x"40",	--7265
		x"71",	--7266
		x"3c",	--7267
		x"40",	--7268
		x"42",	--7269
		x"40",	--7270
		x"0d",	--7271
		x"93",	--7272
		x"24",	--7273
		x"40",	--7274
		x"42",	--7275
		x"40",	--7276
		x"8d",	--7277
		x"40",	--7278
		x"42",	--7279
		x"40",	--7280
		x"0d",	--7281
		x"3c",	--7282
		x"43",	--7283
		x"43",	--7284
		x"4c",	--7285
		x"50",	--7286
		x"00",	--7287
		x"40",	--7288
		x"00",	--7289
		x"5a",	--7290
		x"6b",	--7291
		x"53",	--7292
		x"23",	--7293
		x"48",	--7294
		x"49",	--7295
		x"f3",	--7296
		x"f0",	--7297
		x"80",	--7298
		x"da",	--7299
		x"db",	--7300
		x"43",	--7301
		x"40",	--7302
		x"33",	--7303
		x"12",	--7304
		x"bd",	--7305
		x"41",	--7306
		x"41",	--7307
		x"41",	--7308
		x"41",	--7309
		x"41",	--7310
		x"41",	--7311
		x"12",	--7312
		x"b7",	--7313
		x"41",	--7314
		x"12",	--7315
		x"12",	--7316
		x"12",	--7317
		x"12",	--7318
		x"12",	--7319
		x"12",	--7320
		x"12",	--7321
		x"12",	--7322
		x"83",	--7323
		x"4e",	--7324
		x"4f",	--7325
		x"4e",	--7326
		x"4f",	--7327
		x"f3",	--7328
		x"f0",	--7329
		x"7f",	--7330
		x"49",	--7331
		x"43",	--7332
		x"40",	--7333
		x"00",	--7334
		x"c3",	--7335
		x"10",	--7336
		x"10",	--7337
		x"53",	--7338
		x"23",	--7339
		x"50",	--7340
		x"ff",	--7341
		x"63",	--7342
		x"93",	--7343
		x"38",	--7344
		x"93",	--7345
		x"34",	--7346
		x"90",	--7347
		x"00",	--7348
		x"2c",	--7349
		x"46",	--7350
		x"47",	--7351
		x"93",	--7352
		x"38",	--7353
		x"4c",	--7354
		x"00",	--7355
		x"43",	--7356
		x"40",	--7357
		x"00",	--7358
		x"41",	--7359
		x"f0",	--7360
		x"00",	--7361
		x"3c",	--7362
		x"40",	--7363
		x"f2",	--7364
		x"40",	--7365
		x"71",	--7366
		x"12",	--7367
		x"bd",	--7368
		x"43",	--7369
		x"43",	--7370
		x"12",	--7371
		x"c1",	--7372
		x"93",	--7373
		x"24",	--7374
		x"38",	--7375
		x"93",	--7376
		x"38",	--7377
		x"43",	--7378
		x"43",	--7379
		x"3c",	--7380
		x"93",	--7381
		x"20",	--7382
		x"93",	--7383
		x"24",	--7384
		x"43",	--7385
		x"40",	--7386
		x"bf",	--7387
		x"3c",	--7388
		x"11",	--7389
		x"10",	--7390
		x"53",	--7391
		x"93",	--7392
		x"23",	--7393
		x"48",	--7394
		x"49",	--7395
		x"f6",	--7396
		x"f7",	--7397
		x"93",	--7398
		x"20",	--7399
		x"93",	--7400
		x"24",	--7401
		x"40",	--7402
		x"f2",	--7403
		x"40",	--7404
		x"71",	--7405
		x"12",	--7406
		x"bd",	--7407
		x"43",	--7408
		x"43",	--7409
		x"12",	--7410
		x"c1",	--7411
		x"93",	--7412
		x"24",	--7413
		x"38",	--7414
		x"93",	--7415
		x"34",	--7416
		x"43",	--7417
		x"40",	--7418
		x"00",	--7419
		x"41",	--7420
		x"f0",	--7421
		x"00",	--7422
		x"93",	--7423
		x"24",	--7424
		x"11",	--7425
		x"10",	--7426
		x"53",	--7427
		x"3f",	--7428
		x"56",	--7429
		x"67",	--7430
		x"c8",	--7431
		x"c9",	--7432
		x"3c",	--7433
		x"90",	--7434
		x"7f",	--7435
		x"28",	--7436
		x"4e",	--7437
		x"4f",	--7438
		x"12",	--7439
		x"bd",	--7440
		x"3c",	--7441
		x"4a",	--7442
		x"4b",	--7443
		x"53",	--7444
		x"41",	--7445
		x"41",	--7446
		x"41",	--7447
		x"41",	--7448
		x"41",	--7449
		x"41",	--7450
		x"41",	--7451
		x"41",	--7452
		x"41",	--7453
		x"12",	--7454
		x"b9",	--7455
		x"41",	--7456
		x"12",	--7457
		x"12",	--7458
		x"4e",	--7459
		x"4f",	--7460
		x"43",	--7461
		x"40",	--7462
		x"4f",	--7463
		x"12",	--7464
		x"c1",	--7465
		x"93",	--7466
		x"34",	--7467
		x"4a",	--7468
		x"4b",	--7469
		x"12",	--7470
		x"c3",	--7471
		x"41",	--7472
		x"41",	--7473
		x"41",	--7474
		x"43",	--7475
		x"40",	--7476
		x"4f",	--7477
		x"4a",	--7478
		x"4b",	--7479
		x"12",	--7480
		x"bd",	--7481
		x"12",	--7482
		x"c3",	--7483
		x"53",	--7484
		x"60",	--7485
		x"80",	--7486
		x"41",	--7487
		x"41",	--7488
		x"41",	--7489
		x"12",	--7490
		x"12",	--7491
		x"12",	--7492
		x"12",	--7493
		x"12",	--7494
		x"12",	--7495
		x"12",	--7496
		x"12",	--7497
		x"50",	--7498
		x"ff",	--7499
		x"4d",	--7500
		x"4f",	--7501
		x"93",	--7502
		x"28",	--7503
		x"4e",	--7504
		x"93",	--7505
		x"28",	--7506
		x"92",	--7507
		x"20",	--7508
		x"40",	--7509
		x"bd",	--7510
		x"92",	--7511
		x"24",	--7512
		x"93",	--7513
		x"24",	--7514
		x"93",	--7515
		x"24",	--7516
		x"4f",	--7517
		x"00",	--7518
		x"00",	--7519
		x"4e",	--7520
		x"00",	--7521
		x"4f",	--7522
		x"00",	--7523
		x"4f",	--7524
		x"00",	--7525
		x"4e",	--7526
		x"00",	--7527
		x"4e",	--7528
		x"00",	--7529
		x"41",	--7530
		x"8b",	--7531
		x"4c",	--7532
		x"93",	--7533
		x"38",	--7534
		x"90",	--7535
		x"00",	--7536
		x"34",	--7537
		x"93",	--7538
		x"38",	--7539
		x"46",	--7540
		x"00",	--7541
		x"47",	--7542
		x"00",	--7543
		x"49",	--7544
		x"f0",	--7545
		x"00",	--7546
		x"24",	--7547
		x"46",	--7548
		x"47",	--7549
		x"c3",	--7550
		x"10",	--7551
		x"10",	--7552
		x"53",	--7553
		x"23",	--7554
		x"4a",	--7555
		x"00",	--7556
		x"4b",	--7557
		x"00",	--7558
		x"43",	--7559
		x"43",	--7560
		x"f0",	--7561
		x"00",	--7562
		x"24",	--7563
		x"5c",	--7564
		x"6d",	--7565
		x"53",	--7566
		x"23",	--7567
		x"53",	--7568
		x"63",	--7569
		x"f6",	--7570
		x"f7",	--7571
		x"43",	--7572
		x"43",	--7573
		x"93",	--7574
		x"20",	--7575
		x"93",	--7576
		x"24",	--7577
		x"41",	--7578
		x"00",	--7579
		x"41",	--7580
		x"00",	--7581
		x"da",	--7582
		x"db",	--7583
		x"4f",	--7584
		x"00",	--7585
		x"9e",	--7586
		x"00",	--7587
		x"20",	--7588
		x"4f",	--7589
		x"00",	--7590
		x"41",	--7591
		x"00",	--7592
		x"46",	--7593
		x"47",	--7594
		x"54",	--7595
		x"65",	--7596
		x"4e",	--7597
		x"00",	--7598
		x"4f",	--7599
		x"00",	--7600
		x"40",	--7601
		x"00",	--7602
		x"00",	--7603
		x"93",	--7604
		x"38",	--7605
		x"48",	--7606
		x"50",	--7607
		x"00",	--7608
		x"41",	--7609
		x"41",	--7610
		x"41",	--7611
		x"41",	--7612
		x"41",	--7613
		x"41",	--7614
		x"41",	--7615
		x"41",	--7616
		x"41",	--7617
		x"91",	--7618
		x"38",	--7619
		x"4b",	--7620
		x"00",	--7621
		x"43",	--7622
		x"43",	--7623
		x"4f",	--7624
		x"00",	--7625
		x"9e",	--7626
		x"00",	--7627
		x"27",	--7628
		x"93",	--7629
		x"24",	--7630
		x"46",	--7631
		x"47",	--7632
		x"84",	--7633
		x"75",	--7634
		x"93",	--7635
		x"38",	--7636
		x"43",	--7637
		x"00",	--7638
		x"41",	--7639
		x"00",	--7640
		x"4e",	--7641
		x"00",	--7642
		x"4f",	--7643
		x"00",	--7644
		x"4e",	--7645
		x"4f",	--7646
		x"53",	--7647
		x"63",	--7648
		x"90",	--7649
		x"3f",	--7650
		x"28",	--7651
		x"90",	--7652
		x"40",	--7653
		x"2c",	--7654
		x"93",	--7655
		x"2c",	--7656
		x"48",	--7657
		x"00",	--7658
		x"53",	--7659
		x"5e",	--7660
		x"6f",	--7661
		x"4b",	--7662
		x"53",	--7663
		x"4e",	--7664
		x"4f",	--7665
		x"53",	--7666
		x"63",	--7667
		x"90",	--7668
		x"3f",	--7669
		x"2b",	--7670
		x"24",	--7671
		x"4e",	--7672
		x"00",	--7673
		x"4f",	--7674
		x"00",	--7675
		x"4a",	--7676
		x"00",	--7677
		x"40",	--7678
		x"00",	--7679
		x"00",	--7680
		x"93",	--7681
		x"37",	--7682
		x"4e",	--7683
		x"4f",	--7684
		x"f3",	--7685
		x"f3",	--7686
		x"c3",	--7687
		x"10",	--7688
		x"10",	--7689
		x"4c",	--7690
		x"4d",	--7691
		x"de",	--7692
		x"df",	--7693
		x"4a",	--7694
		x"00",	--7695
		x"4b",	--7696
		x"00",	--7697
		x"53",	--7698
		x"00",	--7699
		x"48",	--7700
		x"3f",	--7701
		x"93",	--7702
		x"23",	--7703
		x"4f",	--7704
		x"00",	--7705
		x"4f",	--7706
		x"00",	--7707
		x"00",	--7708
		x"4f",	--7709
		x"00",	--7710
		x"00",	--7711
		x"4f",	--7712
		x"00",	--7713
		x"00",	--7714
		x"4e",	--7715
		x"00",	--7716
		x"ff",	--7717
		x"00",	--7718
		x"4e",	--7719
		x"00",	--7720
		x"4d",	--7721
		x"3f",	--7722
		x"43",	--7723
		x"43",	--7724
		x"3f",	--7725
		x"e3",	--7726
		x"53",	--7727
		x"90",	--7728
		x"00",	--7729
		x"37",	--7730
		x"3f",	--7731
		x"93",	--7732
		x"2b",	--7733
		x"3f",	--7734
		x"44",	--7735
		x"45",	--7736
		x"86",	--7737
		x"77",	--7738
		x"3f",	--7739
		x"4e",	--7740
		x"3f",	--7741
		x"43",	--7742
		x"00",	--7743
		x"41",	--7744
		x"00",	--7745
		x"e3",	--7746
		x"e3",	--7747
		x"53",	--7748
		x"63",	--7749
		x"4e",	--7750
		x"00",	--7751
		x"4f",	--7752
		x"00",	--7753
		x"3f",	--7754
		x"93",	--7755
		x"27",	--7756
		x"59",	--7757
		x"00",	--7758
		x"44",	--7759
		x"00",	--7760
		x"45",	--7761
		x"00",	--7762
		x"49",	--7763
		x"f0",	--7764
		x"00",	--7765
		x"24",	--7766
		x"4d",	--7767
		x"44",	--7768
		x"45",	--7769
		x"c3",	--7770
		x"10",	--7771
		x"10",	--7772
		x"53",	--7773
		x"23",	--7774
		x"4c",	--7775
		x"00",	--7776
		x"4d",	--7777
		x"00",	--7778
		x"43",	--7779
		x"43",	--7780
		x"f0",	--7781
		x"00",	--7782
		x"24",	--7783
		x"5c",	--7784
		x"6d",	--7785
		x"53",	--7786
		x"23",	--7787
		x"53",	--7788
		x"63",	--7789
		x"f4",	--7790
		x"f5",	--7791
		x"43",	--7792
		x"43",	--7793
		x"93",	--7794
		x"20",	--7795
		x"93",	--7796
		x"20",	--7797
		x"43",	--7798
		x"43",	--7799
		x"41",	--7800
		x"00",	--7801
		x"41",	--7802
		x"00",	--7803
		x"da",	--7804
		x"db",	--7805
		x"3f",	--7806
		x"43",	--7807
		x"43",	--7808
		x"3f",	--7809
		x"92",	--7810
		x"23",	--7811
		x"9e",	--7812
		x"00",	--7813
		x"00",	--7814
		x"27",	--7815
		x"40",	--7816
		x"db",	--7817
		x"3f",	--7818
		x"50",	--7819
		x"ff",	--7820
		x"4e",	--7821
		x"00",	--7822
		x"4f",	--7823
		x"00",	--7824
		x"4c",	--7825
		x"00",	--7826
		x"4d",	--7827
		x"00",	--7828
		x"41",	--7829
		x"50",	--7830
		x"00",	--7831
		x"41",	--7832
		x"52",	--7833
		x"12",	--7834
		x"c7",	--7835
		x"41",	--7836
		x"50",	--7837
		x"00",	--7838
		x"41",	--7839
		x"12",	--7840
		x"c7",	--7841
		x"41",	--7842
		x"52",	--7843
		x"41",	--7844
		x"50",	--7845
		x"00",	--7846
		x"41",	--7847
		x"50",	--7848
		x"00",	--7849
		x"12",	--7850
		x"ba",	--7851
		x"12",	--7852
		x"c5",	--7853
		x"50",	--7854
		x"00",	--7855
		x"41",	--7856
		x"50",	--7857
		x"ff",	--7858
		x"4e",	--7859
		x"00",	--7860
		x"4f",	--7861
		x"00",	--7862
		x"4c",	--7863
		x"00",	--7864
		x"4d",	--7865
		x"00",	--7866
		x"41",	--7867
		x"50",	--7868
		x"00",	--7869
		x"41",	--7870
		x"52",	--7871
		x"12",	--7872
		x"c7",	--7873
		x"41",	--7874
		x"50",	--7875
		x"00",	--7876
		x"41",	--7877
		x"12",	--7878
		x"c7",	--7879
		x"e3",	--7880
		x"00",	--7881
		x"41",	--7882
		x"52",	--7883
		x"41",	--7884
		x"50",	--7885
		x"00",	--7886
		x"41",	--7887
		x"50",	--7888
		x"00",	--7889
		x"12",	--7890
		x"ba",	--7891
		x"12",	--7892
		x"c5",	--7893
		x"50",	--7894
		x"00",	--7895
		x"41",	--7896
		x"12",	--7897
		x"12",	--7898
		x"12",	--7899
		x"12",	--7900
		x"12",	--7901
		x"12",	--7902
		x"12",	--7903
		x"12",	--7904
		x"50",	--7905
		x"ff",	--7906
		x"4e",	--7907
		x"00",	--7908
		x"4f",	--7909
		x"00",	--7910
		x"4c",	--7911
		x"00",	--7912
		x"4d",	--7913
		x"00",	--7914
		x"41",	--7915
		x"50",	--7916
		x"00",	--7917
		x"41",	--7918
		x"52",	--7919
		x"12",	--7920
		x"c7",	--7921
		x"41",	--7922
		x"50",	--7923
		x"00",	--7924
		x"41",	--7925
		x"12",	--7926
		x"c7",	--7927
		x"41",	--7928
		x"00",	--7929
		x"93",	--7930
		x"28",	--7931
		x"41",	--7932
		x"00",	--7933
		x"93",	--7934
		x"28",	--7935
		x"92",	--7936
		x"24",	--7937
		x"92",	--7938
		x"24",	--7939
		x"93",	--7940
		x"24",	--7941
		x"93",	--7942
		x"24",	--7943
		x"41",	--7944
		x"00",	--7945
		x"41",	--7946
		x"00",	--7947
		x"41",	--7948
		x"00",	--7949
		x"41",	--7950
		x"00",	--7951
		x"40",	--7952
		x"00",	--7953
		x"43",	--7954
		x"43",	--7955
		x"43",	--7956
		x"43",	--7957
		x"43",	--7958
		x"00",	--7959
		x"43",	--7960
		x"00",	--7961
		x"43",	--7962
		x"43",	--7963
		x"4c",	--7964
		x"00",	--7965
		x"3c",	--7966
		x"58",	--7967
		x"69",	--7968
		x"c3",	--7969
		x"10",	--7970
		x"10",	--7971
		x"53",	--7972
		x"00",	--7973
		x"24",	--7974
		x"b3",	--7975
		x"24",	--7976
		x"58",	--7977
		x"69",	--7978
		x"56",	--7979
		x"67",	--7980
		x"43",	--7981
		x"43",	--7982
		x"99",	--7983
		x"28",	--7984
		x"24",	--7985
		x"43",	--7986
		x"43",	--7987
		x"5c",	--7988
		x"6d",	--7989
		x"56",	--7990
		x"67",	--7991
		x"93",	--7992
		x"37",	--7993
		x"d3",	--7994
		x"d3",	--7995
		x"3f",	--7996
		x"98",	--7997
		x"2b",	--7998
		x"3f",	--7999
		x"4a",	--8000
		x"00",	--8001
		x"4b",	--8002
		x"00",	--8003
		x"4f",	--8004
		x"41",	--8005
		x"00",	--8006
		x"51",	--8007
		x"00",	--8008
		x"4a",	--8009
		x"53",	--8010
		x"46",	--8011
		x"00",	--8012
		x"43",	--8013
		x"91",	--8014
		x"00",	--8015
		x"00",	--8016
		x"24",	--8017
		x"4d",	--8018
		x"00",	--8019
		x"93",	--8020
		x"38",	--8021
		x"90",	--8022
		x"40",	--8023
		x"2c",	--8024
		x"41",	--8025
		x"00",	--8026
		x"53",	--8027
		x"41",	--8028
		x"00",	--8029
		x"41",	--8030
		x"00",	--8031
		x"4d",	--8032
		x"5e",	--8033
		x"6f",	--8034
		x"93",	--8035
		x"38",	--8036
		x"5a",	--8037
		x"6b",	--8038
		x"53",	--8039
		x"90",	--8040
		x"40",	--8041
		x"2b",	--8042
		x"4a",	--8043
		x"00",	--8044
		x"4b",	--8045
		x"00",	--8046
		x"4c",	--8047
		x"00",	--8048
		x"4e",	--8049
		x"4f",	--8050
		x"f0",	--8051
		x"00",	--8052
		x"f3",	--8053
		x"90",	--8054
		x"00",	--8055
		x"24",	--8056
		x"4e",	--8057
		x"00",	--8058
		x"4f",	--8059
		x"00",	--8060
		x"40",	--8061
		x"00",	--8062
		x"00",	--8063
		x"41",	--8064
		x"52",	--8065
		x"12",	--8066
		x"c5",	--8067
		x"50",	--8068
		x"00",	--8069
		x"41",	--8070
		x"41",	--8071
		x"41",	--8072
		x"41",	--8073
		x"41",	--8074
		x"41",	--8075
		x"41",	--8076
		x"41",	--8077
		x"41",	--8078
		x"d3",	--8079
		x"d3",	--8080
		x"3f",	--8081
		x"50",	--8082
		x"00",	--8083
		x"4a",	--8084
		x"b3",	--8085
		x"24",	--8086
		x"41",	--8087
		x"00",	--8088
		x"41",	--8089
		x"00",	--8090
		x"c3",	--8091
		x"10",	--8092
		x"10",	--8093
		x"4c",	--8094
		x"4d",	--8095
		x"d3",	--8096
		x"d0",	--8097
		x"80",	--8098
		x"46",	--8099
		x"00",	--8100
		x"47",	--8101
		x"00",	--8102
		x"c3",	--8103
		x"10",	--8104
		x"10",	--8105
		x"53",	--8106
		x"93",	--8107
		x"3b",	--8108
		x"48",	--8109
		x"00",	--8110
		x"3f",	--8111
		x"93",	--8112
		x"24",	--8113
		x"43",	--8114
		x"91",	--8115
		x"00",	--8116
		x"00",	--8117
		x"24",	--8118
		x"4f",	--8119
		x"00",	--8120
		x"41",	--8121
		x"50",	--8122
		x"00",	--8123
		x"3f",	--8124
		x"93",	--8125
		x"23",	--8126
		x"4e",	--8127
		x"4f",	--8128
		x"f0",	--8129
		x"00",	--8130
		x"f3",	--8131
		x"93",	--8132
		x"23",	--8133
		x"93",	--8134
		x"23",	--8135
		x"93",	--8136
		x"00",	--8137
		x"20",	--8138
		x"93",	--8139
		x"00",	--8140
		x"27",	--8141
		x"50",	--8142
		x"00",	--8143
		x"63",	--8144
		x"f0",	--8145
		x"ff",	--8146
		x"f3",	--8147
		x"3f",	--8148
		x"43",	--8149
		x"3f",	--8150
		x"43",	--8151
		x"3f",	--8152
		x"43",	--8153
		x"91",	--8154
		x"00",	--8155
		x"00",	--8156
		x"24",	--8157
		x"4f",	--8158
		x"00",	--8159
		x"41",	--8160
		x"50",	--8161
		x"00",	--8162
		x"3f",	--8163
		x"43",	--8164
		x"3f",	--8165
		x"93",	--8166
		x"23",	--8167
		x"40",	--8168
		x"db",	--8169
		x"3f",	--8170
		x"12",	--8171
		x"12",	--8172
		x"12",	--8173
		x"12",	--8174
		x"12",	--8175
		x"50",	--8176
		x"ff",	--8177
		x"4e",	--8178
		x"00",	--8179
		x"4f",	--8180
		x"00",	--8181
		x"4c",	--8182
		x"00",	--8183
		x"4d",	--8184
		x"00",	--8185
		x"41",	--8186
		x"50",	--8187
		x"00",	--8188
		x"41",	--8189
		x"52",	--8190
		x"12",	--8191
		x"c7",	--8192
		x"41",	--8193
		x"52",	--8194
		x"41",	--8195
		x"12",	--8196
		x"c7",	--8197
		x"41",	--8198
		x"00",	--8199
		x"93",	--8200
		x"28",	--8201
		x"41",	--8202
		x"00",	--8203
		x"93",	--8204
		x"28",	--8205
		x"e1",	--8206
		x"00",	--8207
		x"00",	--8208
		x"92",	--8209
		x"24",	--8210
		x"93",	--8211
		x"24",	--8212
		x"92",	--8213
		x"24",	--8214
		x"93",	--8215
		x"24",	--8216
		x"41",	--8217
		x"00",	--8218
		x"81",	--8219
		x"00",	--8220
		x"4d",	--8221
		x"00",	--8222
		x"41",	--8223
		x"00",	--8224
		x"41",	--8225
		x"00",	--8226
		x"41",	--8227
		x"00",	--8228
		x"41",	--8229
		x"00",	--8230
		x"99",	--8231
		x"2c",	--8232
		x"5e",	--8233
		x"6f",	--8234
		x"53",	--8235
		x"4d",	--8236
		x"00",	--8237
		x"40",	--8238
		x"00",	--8239
		x"43",	--8240
		x"40",	--8241
		x"40",	--8242
		x"43",	--8243
		x"43",	--8244
		x"3c",	--8245
		x"dc",	--8246
		x"dd",	--8247
		x"88",	--8248
		x"79",	--8249
		x"c3",	--8250
		x"10",	--8251
		x"10",	--8252
		x"5e",	--8253
		x"6f",	--8254
		x"53",	--8255
		x"24",	--8256
		x"99",	--8257
		x"2b",	--8258
		x"23",	--8259
		x"98",	--8260
		x"2b",	--8261
		x"3f",	--8262
		x"9f",	--8263
		x"2b",	--8264
		x"98",	--8265
		x"2f",	--8266
		x"3f",	--8267
		x"4a",	--8268
		x"4b",	--8269
		x"f0",	--8270
		x"00",	--8271
		x"f3",	--8272
		x"90",	--8273
		x"00",	--8274
		x"24",	--8275
		x"4a",	--8276
		x"00",	--8277
		x"4b",	--8278
		x"00",	--8279
		x"41",	--8280
		x"50",	--8281
		x"00",	--8282
		x"12",	--8283
		x"c5",	--8284
		x"50",	--8285
		x"00",	--8286
		x"41",	--8287
		x"41",	--8288
		x"41",	--8289
		x"41",	--8290
		x"41",	--8291
		x"41",	--8292
		x"42",	--8293
		x"00",	--8294
		x"41",	--8295
		x"50",	--8296
		x"00",	--8297
		x"3f",	--8298
		x"9e",	--8299
		x"23",	--8300
		x"40",	--8301
		x"db",	--8302
		x"3f",	--8303
		x"93",	--8304
		x"23",	--8305
		x"4a",	--8306
		x"4b",	--8307
		x"f0",	--8308
		x"00",	--8309
		x"f3",	--8310
		x"93",	--8311
		x"23",	--8312
		x"93",	--8313
		x"23",	--8314
		x"93",	--8315
		x"20",	--8316
		x"93",	--8317
		x"27",	--8318
		x"50",	--8319
		x"00",	--8320
		x"63",	--8321
		x"f0",	--8322
		x"ff",	--8323
		x"f3",	--8324
		x"3f",	--8325
		x"43",	--8326
		x"00",	--8327
		x"43",	--8328
		x"00",	--8329
		x"43",	--8330
		x"00",	--8331
		x"41",	--8332
		x"50",	--8333
		x"00",	--8334
		x"3f",	--8335
		x"41",	--8336
		x"52",	--8337
		x"3f",	--8338
		x"50",	--8339
		x"ff",	--8340
		x"4e",	--8341
		x"00",	--8342
		x"4f",	--8343
		x"00",	--8344
		x"4c",	--8345
		x"00",	--8346
		x"4d",	--8347
		x"00",	--8348
		x"41",	--8349
		x"50",	--8350
		x"00",	--8351
		x"41",	--8352
		x"52",	--8353
		x"12",	--8354
		x"c7",	--8355
		x"41",	--8356
		x"52",	--8357
		x"41",	--8358
		x"12",	--8359
		x"c7",	--8360
		x"93",	--8361
		x"00",	--8362
		x"28",	--8363
		x"93",	--8364
		x"00",	--8365
		x"28",	--8366
		x"41",	--8367
		x"52",	--8368
		x"41",	--8369
		x"50",	--8370
		x"00",	--8371
		x"12",	--8372
		x"c8",	--8373
		x"50",	--8374
		x"00",	--8375
		x"41",	--8376
		x"43",	--8377
		x"3f",	--8378
		x"50",	--8379
		x"ff",	--8380
		x"4e",	--8381
		x"00",	--8382
		x"4f",	--8383
		x"00",	--8384
		x"4c",	--8385
		x"00",	--8386
		x"4d",	--8387
		x"00",	--8388
		x"41",	--8389
		x"50",	--8390
		x"00",	--8391
		x"41",	--8392
		x"52",	--8393
		x"12",	--8394
		x"c7",	--8395
		x"41",	--8396
		x"52",	--8397
		x"41",	--8398
		x"12",	--8399
		x"c7",	--8400
		x"93",	--8401
		x"00",	--8402
		x"28",	--8403
		x"93",	--8404
		x"00",	--8405
		x"28",	--8406
		x"41",	--8407
		x"52",	--8408
		x"41",	--8409
		x"50",	--8410
		x"00",	--8411
		x"12",	--8412
		x"c8",	--8413
		x"50",	--8414
		x"00",	--8415
		x"41",	--8416
		x"43",	--8417
		x"3f",	--8418
		x"50",	--8419
		x"ff",	--8420
		x"4e",	--8421
		x"00",	--8422
		x"4f",	--8423
		x"00",	--8424
		x"4c",	--8425
		x"00",	--8426
		x"4d",	--8427
		x"00",	--8428
		x"41",	--8429
		x"50",	--8430
		x"00",	--8431
		x"41",	--8432
		x"52",	--8433
		x"12",	--8434
		x"c7",	--8435
		x"41",	--8436
		x"52",	--8437
		x"41",	--8438
		x"12",	--8439
		x"c7",	--8440
		x"93",	--8441
		x"00",	--8442
		x"28",	--8443
		x"93",	--8444
		x"00",	--8445
		x"28",	--8446
		x"41",	--8447
		x"52",	--8448
		x"41",	--8449
		x"50",	--8450
		x"00",	--8451
		x"12",	--8452
		x"c8",	--8453
		x"50",	--8454
		x"00",	--8455
		x"41",	--8456
		x"43",	--8457
		x"3f",	--8458
		x"50",	--8459
		x"ff",	--8460
		x"4e",	--8461
		x"00",	--8462
		x"4f",	--8463
		x"00",	--8464
		x"4c",	--8465
		x"00",	--8466
		x"4d",	--8467
		x"00",	--8468
		x"41",	--8469
		x"50",	--8470
		x"00",	--8471
		x"41",	--8472
		x"52",	--8473
		x"12",	--8474
		x"c7",	--8475
		x"41",	--8476
		x"52",	--8477
		x"41",	--8478
		x"12",	--8479
		x"c7",	--8480
		x"93",	--8481
		x"00",	--8482
		x"28",	--8483
		x"93",	--8484
		x"00",	--8485
		x"28",	--8486
		x"41",	--8487
		x"52",	--8488
		x"41",	--8489
		x"50",	--8490
		x"00",	--8491
		x"12",	--8492
		x"c8",	--8493
		x"50",	--8494
		x"00",	--8495
		x"41",	--8496
		x"43",	--8497
		x"3f",	--8498
		x"50",	--8499
		x"ff",	--8500
		x"4e",	--8501
		x"00",	--8502
		x"4f",	--8503
		x"00",	--8504
		x"4c",	--8505
		x"00",	--8506
		x"4d",	--8507
		x"00",	--8508
		x"41",	--8509
		x"50",	--8510
		x"00",	--8511
		x"41",	--8512
		x"52",	--8513
		x"12",	--8514
		x"c7",	--8515
		x"41",	--8516
		x"52",	--8517
		x"41",	--8518
		x"12",	--8519
		x"c7",	--8520
		x"93",	--8521
		x"00",	--8522
		x"28",	--8523
		x"93",	--8524
		x"00",	--8525
		x"28",	--8526
		x"41",	--8527
		x"52",	--8528
		x"41",	--8529
		x"50",	--8530
		x"00",	--8531
		x"12",	--8532
		x"c8",	--8533
		x"50",	--8534
		x"00",	--8535
		x"41",	--8536
		x"43",	--8537
		x"3f",	--8538
		x"12",	--8539
		x"12",	--8540
		x"82",	--8541
		x"40",	--8542
		x"00",	--8543
		x"00",	--8544
		x"4f",	--8545
		x"5d",	--8546
		x"43",	--8547
		x"6d",	--8548
		x"4d",	--8549
		x"4d",	--8550
		x"00",	--8551
		x"93",	--8552
		x"20",	--8553
		x"93",	--8554
		x"20",	--8555
		x"43",	--8556
		x"00",	--8557
		x"41",	--8558
		x"12",	--8559
		x"c5",	--8560
		x"52",	--8561
		x"41",	--8562
		x"41",	--8563
		x"41",	--8564
		x"40",	--8565
		x"00",	--8566
		x"00",	--8567
		x"93",	--8568
		x"20",	--8569
		x"4e",	--8570
		x"4f",	--8571
		x"4a",	--8572
		x"00",	--8573
		x"4b",	--8574
		x"00",	--8575
		x"4a",	--8576
		x"4b",	--8577
		x"12",	--8578
		x"c4",	--8579
		x"53",	--8580
		x"93",	--8581
		x"3b",	--8582
		x"4a",	--8583
		x"00",	--8584
		x"4b",	--8585
		x"00",	--8586
		x"4f",	--8587
		x"f0",	--8588
		x"00",	--8589
		x"20",	--8590
		x"40",	--8591
		x"00",	--8592
		x"8f",	--8593
		x"4e",	--8594
		x"00",	--8595
		x"3f",	--8596
		x"93",	--8597
		x"24",	--8598
		x"4e",	--8599
		x"4f",	--8600
		x"e3",	--8601
		x"e3",	--8602
		x"53",	--8603
		x"63",	--8604
		x"3f",	--8605
		x"51",	--8606
		x"00",	--8607
		x"00",	--8608
		x"61",	--8609
		x"00",	--8610
		x"00",	--8611
		x"53",	--8612
		x"23",	--8613
		x"3f",	--8614
		x"90",	--8615
		x"80",	--8616
		x"23",	--8617
		x"43",	--8618
		x"40",	--8619
		x"cf",	--8620
		x"3f",	--8621
		x"50",	--8622
		x"ff",	--8623
		x"4e",	--8624
		x"00",	--8625
		x"4f",	--8626
		x"00",	--8627
		x"41",	--8628
		x"52",	--8629
		x"41",	--8630
		x"12",	--8631
		x"c7",	--8632
		x"41",	--8633
		x"00",	--8634
		x"93",	--8635
		x"24",	--8636
		x"28",	--8637
		x"92",	--8638
		x"24",	--8639
		x"41",	--8640
		x"00",	--8641
		x"93",	--8642
		x"38",	--8643
		x"90",	--8644
		x"00",	--8645
		x"38",	--8646
		x"93",	--8647
		x"00",	--8648
		x"20",	--8649
		x"43",	--8650
		x"40",	--8651
		x"7f",	--8652
		x"50",	--8653
		x"00",	--8654
		x"41",	--8655
		x"41",	--8656
		x"00",	--8657
		x"41",	--8658
		x"00",	--8659
		x"40",	--8660
		x"00",	--8661
		x"8d",	--8662
		x"4c",	--8663
		x"f0",	--8664
		x"00",	--8665
		x"20",	--8666
		x"93",	--8667
		x"00",	--8668
		x"27",	--8669
		x"e3",	--8670
		x"e3",	--8671
		x"53",	--8672
		x"63",	--8673
		x"50",	--8674
		x"00",	--8675
		x"41",	--8676
		x"43",	--8677
		x"43",	--8678
		x"50",	--8679
		x"00",	--8680
		x"41",	--8681
		x"c3",	--8682
		x"10",	--8683
		x"10",	--8684
		x"53",	--8685
		x"23",	--8686
		x"3f",	--8687
		x"43",	--8688
		x"40",	--8689
		x"80",	--8690
		x"50",	--8691
		x"00",	--8692
		x"41",	--8693
		x"12",	--8694
		x"12",	--8695
		x"12",	--8696
		x"12",	--8697
		x"82",	--8698
		x"4e",	--8699
		x"4f",	--8700
		x"43",	--8701
		x"00",	--8702
		x"93",	--8703
		x"20",	--8704
		x"93",	--8705
		x"20",	--8706
		x"43",	--8707
		x"00",	--8708
		x"41",	--8709
		x"12",	--8710
		x"c5",	--8711
		x"52",	--8712
		x"41",	--8713
		x"41",	--8714
		x"41",	--8715
		x"41",	--8716
		x"41",	--8717
		x"40",	--8718
		x"00",	--8719
		x"00",	--8720
		x"40",	--8721
		x"00",	--8722
		x"00",	--8723
		x"4a",	--8724
		x"00",	--8725
		x"4b",	--8726
		x"00",	--8727
		x"4a",	--8728
		x"4b",	--8729
		x"12",	--8730
		x"c4",	--8731
		x"53",	--8732
		x"93",	--8733
		x"38",	--8734
		x"27",	--8735
		x"4a",	--8736
		x"00",	--8737
		x"4b",	--8738
		x"00",	--8739
		x"4f",	--8740
		x"f0",	--8741
		x"00",	--8742
		x"20",	--8743
		x"40",	--8744
		x"00",	--8745
		x"8f",	--8746
		x"4e",	--8747
		x"00",	--8748
		x"3f",	--8749
		x"51",	--8750
		x"00",	--8751
		x"00",	--8752
		x"61",	--8753
		x"00",	--8754
		x"00",	--8755
		x"53",	--8756
		x"23",	--8757
		x"3f",	--8758
		x"4f",	--8759
		x"e3",	--8760
		x"53",	--8761
		x"43",	--8762
		x"43",	--8763
		x"4e",	--8764
		x"f0",	--8765
		x"00",	--8766
		x"24",	--8767
		x"5c",	--8768
		x"6d",	--8769
		x"53",	--8770
		x"23",	--8771
		x"53",	--8772
		x"63",	--8773
		x"fa",	--8774
		x"fb",	--8775
		x"43",	--8776
		x"43",	--8777
		x"93",	--8778
		x"20",	--8779
		x"93",	--8780
		x"20",	--8781
		x"43",	--8782
		x"43",	--8783
		x"f0",	--8784
		x"00",	--8785
		x"20",	--8786
		x"48",	--8787
		x"49",	--8788
		x"da",	--8789
		x"db",	--8790
		x"4d",	--8791
		x"00",	--8792
		x"4e",	--8793
		x"00",	--8794
		x"40",	--8795
		x"00",	--8796
		x"8f",	--8797
		x"4e",	--8798
		x"00",	--8799
		x"3f",	--8800
		x"c3",	--8801
		x"10",	--8802
		x"10",	--8803
		x"53",	--8804
		x"23",	--8805
		x"3f",	--8806
		x"12",	--8807
		x"12",	--8808
		x"12",	--8809
		x"93",	--8810
		x"2c",	--8811
		x"90",	--8812
		x"01",	--8813
		x"28",	--8814
		x"40",	--8815
		x"00",	--8816
		x"43",	--8817
		x"42",	--8818
		x"4e",	--8819
		x"4f",	--8820
		x"49",	--8821
		x"93",	--8822
		x"20",	--8823
		x"50",	--8824
		x"db",	--8825
		x"4c",	--8826
		x"43",	--8827
		x"8e",	--8828
		x"7f",	--8829
		x"4a",	--8830
		x"41",	--8831
		x"41",	--8832
		x"41",	--8833
		x"41",	--8834
		x"90",	--8835
		x"01",	--8836
		x"28",	--8837
		x"42",	--8838
		x"43",	--8839
		x"40",	--8840
		x"00",	--8841
		x"4e",	--8842
		x"4f",	--8843
		x"49",	--8844
		x"93",	--8845
		x"27",	--8846
		x"c3",	--8847
		x"10",	--8848
		x"10",	--8849
		x"53",	--8850
		x"23",	--8851
		x"3f",	--8852
		x"40",	--8853
		x"00",	--8854
		x"43",	--8855
		x"40",	--8856
		x"00",	--8857
		x"3f",	--8858
		x"40",	--8859
		x"00",	--8860
		x"43",	--8861
		x"43",	--8862
		x"3f",	--8863
		x"12",	--8864
		x"12",	--8865
		x"12",	--8866
		x"12",	--8867
		x"12",	--8868
		x"4f",	--8869
		x"4f",	--8870
		x"00",	--8871
		x"4f",	--8872
		x"00",	--8873
		x"4d",	--8874
		x"00",	--8875
		x"4d",	--8876
		x"93",	--8877
		x"28",	--8878
		x"92",	--8879
		x"24",	--8880
		x"93",	--8881
		x"24",	--8882
		x"93",	--8883
		x"24",	--8884
		x"4d",	--8885
		x"00",	--8886
		x"90",	--8887
		x"ff",	--8888
		x"38",	--8889
		x"90",	--8890
		x"00",	--8891
		x"34",	--8892
		x"4e",	--8893
		x"4f",	--8894
		x"f0",	--8895
		x"00",	--8896
		x"f3",	--8897
		x"90",	--8898
		x"00",	--8899
		x"24",	--8900
		x"50",	--8901
		x"00",	--8902
		x"63",	--8903
		x"93",	--8904
		x"38",	--8905
		x"4b",	--8906
		x"50",	--8907
		x"00",	--8908
		x"c3",	--8909
		x"10",	--8910
		x"10",	--8911
		x"c3",	--8912
		x"10",	--8913
		x"10",	--8914
		x"c3",	--8915
		x"10",	--8916
		x"10",	--8917
		x"c3",	--8918
		x"10",	--8919
		x"10",	--8920
		x"c3",	--8921
		x"10",	--8922
		x"10",	--8923
		x"c3",	--8924
		x"10",	--8925
		x"10",	--8926
		x"c3",	--8927
		x"10",	--8928
		x"10",	--8929
		x"f3",	--8930
		x"f0",	--8931
		x"00",	--8932
		x"4d",	--8933
		x"3c",	--8934
		x"93",	--8935
		x"23",	--8936
		x"43",	--8937
		x"43",	--8938
		x"43",	--8939
		x"4d",	--8940
		x"5d",	--8941
		x"5d",	--8942
		x"5d",	--8943
		x"5d",	--8944
		x"5d",	--8945
		x"5d",	--8946
		x"5d",	--8947
		x"4f",	--8948
		x"f0",	--8949
		x"00",	--8950
		x"dd",	--8951
		x"4a",	--8952
		x"11",	--8953
		x"43",	--8954
		x"10",	--8955
		x"4c",	--8956
		x"df",	--8957
		x"4d",	--8958
		x"41",	--8959
		x"41",	--8960
		x"41",	--8961
		x"41",	--8962
		x"41",	--8963
		x"41",	--8964
		x"93",	--8965
		x"23",	--8966
		x"4e",	--8967
		x"4f",	--8968
		x"f0",	--8969
		x"00",	--8970
		x"f3",	--8971
		x"93",	--8972
		x"20",	--8973
		x"93",	--8974
		x"27",	--8975
		x"50",	--8976
		x"00",	--8977
		x"63",	--8978
		x"3f",	--8979
		x"c3",	--8980
		x"10",	--8981
		x"10",	--8982
		x"4b",	--8983
		x"50",	--8984
		x"00",	--8985
		x"3f",	--8986
		x"43",	--8987
		x"43",	--8988
		x"43",	--8989
		x"3f",	--8990
		x"d3",	--8991
		x"d0",	--8992
		x"00",	--8993
		x"f3",	--8994
		x"f0",	--8995
		x"00",	--8996
		x"43",	--8997
		x"3f",	--8998
		x"40",	--8999
		x"ff",	--9000
		x"8b",	--9001
		x"90",	--9002
		x"00",	--9003
		x"34",	--9004
		x"4e",	--9005
		x"4f",	--9006
		x"47",	--9007
		x"f0",	--9008
		x"00",	--9009
		x"24",	--9010
		x"c3",	--9011
		x"10",	--9012
		x"10",	--9013
		x"53",	--9014
		x"23",	--9015
		x"43",	--9016
		x"43",	--9017
		x"f0",	--9018
		x"00",	--9019
		x"24",	--9020
		x"58",	--9021
		x"69",	--9022
		x"53",	--9023
		x"23",	--9024
		x"53",	--9025
		x"63",	--9026
		x"fe",	--9027
		x"ff",	--9028
		x"43",	--9029
		x"43",	--9030
		x"93",	--9031
		x"20",	--9032
		x"93",	--9033
		x"20",	--9034
		x"43",	--9035
		x"43",	--9036
		x"4e",	--9037
		x"4f",	--9038
		x"dc",	--9039
		x"dd",	--9040
		x"48",	--9041
		x"49",	--9042
		x"f0",	--9043
		x"00",	--9044
		x"f3",	--9045
		x"90",	--9046
		x"00",	--9047
		x"24",	--9048
		x"50",	--9049
		x"00",	--9050
		x"63",	--9051
		x"48",	--9052
		x"49",	--9053
		x"c3",	--9054
		x"10",	--9055
		x"10",	--9056
		x"c3",	--9057
		x"10",	--9058
		x"10",	--9059
		x"c3",	--9060
		x"10",	--9061
		x"10",	--9062
		x"c3",	--9063
		x"10",	--9064
		x"10",	--9065
		x"c3",	--9066
		x"10",	--9067
		x"10",	--9068
		x"c3",	--9069
		x"10",	--9070
		x"10",	--9071
		x"c3",	--9072
		x"10",	--9073
		x"10",	--9074
		x"f3",	--9075
		x"f0",	--9076
		x"00",	--9077
		x"43",	--9078
		x"90",	--9079
		x"40",	--9080
		x"2f",	--9081
		x"43",	--9082
		x"3f",	--9083
		x"43",	--9084
		x"43",	--9085
		x"3f",	--9086
		x"93",	--9087
		x"23",	--9088
		x"48",	--9089
		x"49",	--9090
		x"f0",	--9091
		x"00",	--9092
		x"f3",	--9093
		x"93",	--9094
		x"24",	--9095
		x"50",	--9096
		x"00",	--9097
		x"63",	--9098
		x"3f",	--9099
		x"93",	--9100
		x"27",	--9101
		x"3f",	--9102
		x"12",	--9103
		x"12",	--9104
		x"4f",	--9105
		x"4f",	--9106
		x"00",	--9107
		x"f0",	--9108
		x"00",	--9109
		x"4f",	--9110
		x"00",	--9111
		x"c3",	--9112
		x"10",	--9113
		x"c3",	--9114
		x"10",	--9115
		x"c3",	--9116
		x"10",	--9117
		x"c3",	--9118
		x"10",	--9119
		x"c3",	--9120
		x"10",	--9121
		x"c3",	--9122
		x"10",	--9123
		x"c3",	--9124
		x"10",	--9125
		x"4d",	--9126
		x"4f",	--9127
		x"00",	--9128
		x"b0",	--9129
		x"00",	--9130
		x"43",	--9131
		x"6f",	--9132
		x"4f",	--9133
		x"00",	--9134
		x"93",	--9135
		x"20",	--9136
		x"93",	--9137
		x"24",	--9138
		x"40",	--9139
		x"ff",	--9140
		x"00",	--9141
		x"4a",	--9142
		x"4b",	--9143
		x"5c",	--9144
		x"6d",	--9145
		x"5c",	--9146
		x"6d",	--9147
		x"5c",	--9148
		x"6d",	--9149
		x"5c",	--9150
		x"6d",	--9151
		x"5c",	--9152
		x"6d",	--9153
		x"5c",	--9154
		x"6d",	--9155
		x"5c",	--9156
		x"6d",	--9157
		x"40",	--9158
		x"00",	--9159
		x"00",	--9160
		x"90",	--9161
		x"40",	--9162
		x"2c",	--9163
		x"40",	--9164
		x"ff",	--9165
		x"5c",	--9166
		x"6d",	--9167
		x"4f",	--9168
		x"53",	--9169
		x"90",	--9170
		x"40",	--9171
		x"2b",	--9172
		x"4a",	--9173
		x"00",	--9174
		x"4c",	--9175
		x"00",	--9176
		x"4d",	--9177
		x"00",	--9178
		x"41",	--9179
		x"41",	--9180
		x"41",	--9181
		x"90",	--9182
		x"00",	--9183
		x"24",	--9184
		x"50",	--9185
		x"ff",	--9186
		x"4d",	--9187
		x"00",	--9188
		x"40",	--9189
		x"00",	--9190
		x"00",	--9191
		x"4a",	--9192
		x"4b",	--9193
		x"5c",	--9194
		x"6d",	--9195
		x"5c",	--9196
		x"6d",	--9197
		x"5c",	--9198
		x"6d",	--9199
		x"5c",	--9200
		x"6d",	--9201
		x"5c",	--9202
		x"6d",	--9203
		x"5c",	--9204
		x"6d",	--9205
		x"5c",	--9206
		x"6d",	--9207
		x"4c",	--9208
		x"4d",	--9209
		x"d3",	--9210
		x"d0",	--9211
		x"40",	--9212
		x"4a",	--9213
		x"00",	--9214
		x"4b",	--9215
		x"00",	--9216
		x"41",	--9217
		x"41",	--9218
		x"41",	--9219
		x"93",	--9220
		x"23",	--9221
		x"43",	--9222
		x"00",	--9223
		x"41",	--9224
		x"41",	--9225
		x"41",	--9226
		x"93",	--9227
		x"24",	--9228
		x"4a",	--9229
		x"4b",	--9230
		x"f3",	--9231
		x"f0",	--9232
		x"00",	--9233
		x"93",	--9234
		x"20",	--9235
		x"93",	--9236
		x"24",	--9237
		x"43",	--9238
		x"00",	--9239
		x"3f",	--9240
		x"93",	--9241
		x"23",	--9242
		x"42",	--9243
		x"00",	--9244
		x"3f",	--9245
		x"43",	--9246
		x"00",	--9247
		x"3f",	--9248
		x"12",	--9249
		x"4f",	--9250
		x"93",	--9251
		x"28",	--9252
		x"4e",	--9253
		x"93",	--9254
		x"28",	--9255
		x"92",	--9256
		x"24",	--9257
		x"92",	--9258
		x"24",	--9259
		x"93",	--9260
		x"24",	--9261
		x"93",	--9262
		x"24",	--9263
		x"4f",	--9264
		x"00",	--9265
		x"9e",	--9266
		x"00",	--9267
		x"24",	--9268
		x"93",	--9269
		x"20",	--9270
		x"43",	--9271
		x"4e",	--9272
		x"41",	--9273
		x"41",	--9274
		x"93",	--9275
		x"24",	--9276
		x"93",	--9277
		x"00",	--9278
		x"23",	--9279
		x"43",	--9280
		x"4e",	--9281
		x"41",	--9282
		x"41",	--9283
		x"93",	--9284
		x"00",	--9285
		x"27",	--9286
		x"43",	--9287
		x"3f",	--9288
		x"4f",	--9289
		x"00",	--9290
		x"4e",	--9291
		x"00",	--9292
		x"9b",	--9293
		x"3b",	--9294
		x"9c",	--9295
		x"38",	--9296
		x"4f",	--9297
		x"00",	--9298
		x"4f",	--9299
		x"00",	--9300
		x"4e",	--9301
		x"00",	--9302
		x"4e",	--9303
		x"00",	--9304
		x"9f",	--9305
		x"2b",	--9306
		x"9e",	--9307
		x"28",	--9308
		x"9b",	--9309
		x"2b",	--9310
		x"9e",	--9311
		x"28",	--9312
		x"9f",	--9313
		x"28",	--9314
		x"9c",	--9315
		x"28",	--9316
		x"43",	--9317
		x"3f",	--9318
		x"93",	--9319
		x"23",	--9320
		x"43",	--9321
		x"3f",	--9322
		x"92",	--9323
		x"23",	--9324
		x"4e",	--9325
		x"00",	--9326
		x"4f",	--9327
		x"00",	--9328
		x"8f",	--9329
		x"3f",	--9330
		x"42",	--9331
		x"02",	--9332
		x"93",	--9333
		x"38",	--9334
		x"42",	--9335
		x"02",	--9336
		x"4f",	--9337
		x"00",	--9338
		x"53",	--9339
		x"4d",	--9340
		x"02",	--9341
		x"53",	--9342
		x"4e",	--9343
		x"02",	--9344
		x"41",	--9345
		x"43",	--9346
		x"41",	--9347
		x"12",	--9348
		x"12",	--9349
		x"83",	--9350
		x"4e",	--9351
		x"00",	--9352
		x"42",	--9353
		x"02",	--9354
		x"42",	--9355
		x"02",	--9356
		x"4e",	--9357
		x"4f",	--9358
		x"40",	--9359
		x"c8",	--9360
		x"12",	--9361
		x"cb",	--9362
		x"9b",	--9363
		x"38",	--9364
		x"4a",	--9365
		x"5b",	--9366
		x"43",	--9367
		x"ff",	--9368
		x"3c",	--9369
		x"42",	--9370
		x"02",	--9371
		x"43",	--9372
		x"00",	--9373
		x"53",	--9374
		x"41",	--9375
		x"41",	--9376
		x"41",	--9377
		x"41",	--9378
		x"00",	--9379
		x"02",	--9380
		x"40",	--9381
		x"7f",	--9382
		x"02",	--9383
		x"41",	--9384
		x"50",	--9385
		x"00",	--9386
		x"41",	--9387
		x"00",	--9388
		x"12",	--9389
		x"c9",	--9390
		x"41",	--9391
		x"41",	--9392
		x"00",	--9393
		x"02",	--9394
		x"41",	--9395
		x"00",	--9396
		x"02",	--9397
		x"41",	--9398
		x"52",	--9399
		x"41",	--9400
		x"00",	--9401
		x"12",	--9402
		x"c9",	--9403
		x"41",	--9404
		x"4e",	--9405
		x"4f",	--9406
		x"02",	--9407
		x"40",	--9408
		x"7f",	--9409
		x"02",	--9410
		x"4d",	--9411
		x"4c",	--9412
		x"12",	--9413
		x"c9",	--9414
		x"41",	--9415
		x"4f",	--9416
		x"02",	--9417
		x"4e",	--9418
		x"02",	--9419
		x"4c",	--9420
		x"4d",	--9421
		x"12",	--9422
		x"c9",	--9423
		x"41",	--9424
		x"12",	--9425
		x"12",	--9426
		x"12",	--9427
		x"12",	--9428
		x"12",	--9429
		x"12",	--9430
		x"12",	--9431
		x"12",	--9432
		x"82",	--9433
		x"4f",	--9434
		x"4e",	--9435
		x"00",	--9436
		x"4d",	--9437
		x"41",	--9438
		x"00",	--9439
		x"41",	--9440
		x"00",	--9441
		x"4d",	--9442
		x"4d",	--9443
		x"10",	--9444
		x"44",	--9445
		x"4f",	--9446
		x"b0",	--9447
		x"00",	--9448
		x"24",	--9449
		x"40",	--9450
		x"00",	--9451
		x"00",	--9452
		x"4f",	--9453
		x"10",	--9454
		x"f3",	--9455
		x"24",	--9456
		x"40",	--9457
		x"00",	--9458
		x"3c",	--9459
		x"40",	--9460
		x"00",	--9461
		x"4e",	--9462
		x"00",	--9463
		x"41",	--9464
		x"53",	--9465
		x"3c",	--9466
		x"f0",	--9467
		x"00",	--9468
		x"24",	--9469
		x"40",	--9470
		x"00",	--9471
		x"00",	--9472
		x"3c",	--9473
		x"93",	--9474
		x"24",	--9475
		x"4d",	--9476
		x"00",	--9477
		x"41",	--9478
		x"53",	--9479
		x"3c",	--9480
		x"41",	--9481
		x"4c",	--9482
		x"10",	--9483
		x"11",	--9484
		x"10",	--9485
		x"11",	--9486
		x"4c",	--9487
		x"41",	--9488
		x"41",	--9489
		x"10",	--9490
		x"11",	--9491
		x"10",	--9492
		x"11",	--9493
		x"4c",	--9494
		x"86",	--9495
		x"77",	--9496
		x"4f",	--9497
		x"10",	--9498
		x"4e",	--9499
		x"00",	--9500
		x"f2",	--9501
		x"24",	--9502
		x"45",	--9503
		x"3c",	--9504
		x"43",	--9505
		x"4f",	--9506
		x"b0",	--9507
		x"00",	--9508
		x"20",	--9509
		x"41",	--9510
		x"00",	--9511
		x"53",	--9512
		x"53",	--9513
		x"93",	--9514
		x"00",	--9515
		x"23",	--9516
		x"81",	--9517
		x"00",	--9518
		x"9a",	--9519
		x"28",	--9520
		x"8a",	--9521
		x"3c",	--9522
		x"43",	--9523
		x"b3",	--9524
		x"00",	--9525
		x"24",	--9526
		x"95",	--9527
		x"28",	--9528
		x"85",	--9529
		x"3c",	--9530
		x"43",	--9531
		x"4d",	--9532
		x"9d",	--9533
		x"2c",	--9534
		x"47",	--9535
		x"93",	--9536
		x"38",	--9537
		x"40",	--9538
		x"00",	--9539
		x"00",	--9540
		x"43",	--9541
		x"43",	--9542
		x"3c",	--9543
		x"41",	--9544
		x"56",	--9545
		x"4f",	--9546
		x"11",	--9547
		x"53",	--9548
		x"12",	--9549
		x"3c",	--9550
		x"43",	--9551
		x"9a",	--9552
		x"3b",	--9553
		x"4a",	--9554
		x"40",	--9555
		x"00",	--9556
		x"00",	--9557
		x"8b",	--9558
		x"3c",	--9559
		x"41",	--9560
		x"00",	--9561
		x"11",	--9562
		x"12",	--9563
		x"53",	--9564
		x"45",	--9565
		x"5b",	--9566
		x"99",	--9567
		x"2b",	--9568
		x"3c",	--9569
		x"43",	--9570
		x"43",	--9571
		x"3c",	--9572
		x"53",	--9573
		x"41",	--9574
		x"56",	--9575
		x"4f",	--9576
		x"11",	--9577
		x"53",	--9578
		x"12",	--9579
		x"9a",	--9580
		x"3b",	--9581
		x"b3",	--9582
		x"00",	--9583
		x"24",	--9584
		x"44",	--9585
		x"3c",	--9586
		x"41",	--9587
		x"00",	--9588
		x"8b",	--9589
		x"3c",	--9590
		x"40",	--9591
		x"00",	--9592
		x"12",	--9593
		x"53",	--9594
		x"93",	--9595
		x"23",	--9596
		x"44",	--9597
		x"54",	--9598
		x"3f",	--9599
		x"53",	--9600
		x"11",	--9601
		x"12",	--9602
		x"53",	--9603
		x"4a",	--9604
		x"5b",	--9605
		x"4f",	--9606
		x"93",	--9607
		x"24",	--9608
		x"93",	--9609
		x"23",	--9610
		x"3c",	--9611
		x"40",	--9612
		x"00",	--9613
		x"12",	--9614
		x"53",	--9615
		x"99",	--9616
		x"2b",	--9617
		x"4b",	--9618
		x"52",	--9619
		x"41",	--9620
		x"41",	--9621
		x"41",	--9622
		x"41",	--9623
		x"41",	--9624
		x"41",	--9625
		x"41",	--9626
		x"41",	--9627
		x"41",	--9628
		x"12",	--9629
		x"12",	--9630
		x"12",	--9631
		x"12",	--9632
		x"12",	--9633
		x"12",	--9634
		x"12",	--9635
		x"12",	--9636
		x"50",	--9637
		x"ff",	--9638
		x"4f",	--9639
		x"00",	--9640
		x"4e",	--9641
		x"4d",	--9642
		x"4e",	--9643
		x"00",	--9644
		x"43",	--9645
		x"00",	--9646
		x"43",	--9647
		x"00",	--9648
		x"43",	--9649
		x"00",	--9650
		x"43",	--9651
		x"00",	--9652
		x"43",	--9653
		x"00",	--9654
		x"43",	--9655
		x"00",	--9656
		x"43",	--9657
		x"43",	--9658
		x"00",	--9659
		x"41",	--9660
		x"50",	--9661
		x"00",	--9662
		x"4e",	--9663
		x"00",	--9664
		x"40",	--9665
		x"d1",	--9666
		x"46",	--9667
		x"53",	--9668
		x"4f",	--9669
		x"00",	--9670
		x"93",	--9671
		x"20",	--9672
		x"90",	--9673
		x"00",	--9674
		x"20",	--9675
		x"43",	--9676
		x"00",	--9677
		x"43",	--9678
		x"00",	--9679
		x"46",	--9680
		x"00",	--9681
		x"43",	--9682
		x"00",	--9683
		x"43",	--9684
		x"00",	--9685
		x"43",	--9686
		x"00",	--9687
		x"43",	--9688
		x"00",	--9689
		x"43",	--9690
		x"00",	--9691
		x"40",	--9692
		x"d1",	--9693
		x"47",	--9694
		x"11",	--9695
		x"4e",	--9696
		x"12",	--9697
		x"00",	--9698
		x"53",	--9699
		x"00",	--9700
		x"40",	--9701
		x"d1",	--9702
		x"90",	--9703
		x"00",	--9704
		x"24",	--9705
		x"90",	--9706
		x"00",	--9707
		x"34",	--9708
		x"90",	--9709
		x"00",	--9710
		x"24",	--9711
		x"90",	--9712
		x"00",	--9713
		x"34",	--9714
		x"90",	--9715
		x"00",	--9716
		x"24",	--9717
		x"90",	--9718
		x"00",	--9719
		x"34",	--9720
		x"90",	--9721
		x"00",	--9722
		x"24",	--9723
		x"90",	--9724
		x"00",	--9725
		x"27",	--9726
		x"90",	--9727
		x"00",	--9728
		x"20",	--9729
		x"3c",	--9730
		x"90",	--9731
		x"00",	--9732
		x"24",	--9733
		x"90",	--9734
		x"00",	--9735
		x"24",	--9736
		x"90",	--9737
		x"00",	--9738
		x"20",	--9739
		x"3c",	--9740
		x"90",	--9741
		x"00",	--9742
		x"38",	--9743
		x"90",	--9744
		x"00",	--9745
		x"20",	--9746
		x"3c",	--9747
		x"90",	--9748
		x"00",	--9749
		x"24",	--9750
		x"90",	--9751
		x"00",	--9752
		x"34",	--9753
		x"90",	--9754
		x"00",	--9755
		x"24",	--9756
		x"90",	--9757
		x"00",	--9758
		x"24",	--9759
		x"90",	--9760
		x"00",	--9761
		x"20",	--9762
		x"3c",	--9763
		x"90",	--9764
		x"00",	--9765
		x"24",	--9766
		x"90",	--9767
		x"00",	--9768
		x"34",	--9769
		x"90",	--9770
		x"00",	--9771
		x"20",	--9772
		x"3c",	--9773
		x"90",	--9774
		x"00",	--9775
		x"24",	--9776
		x"90",	--9777
		x"00",	--9778
		x"24",	--9779
		x"41",	--9780
		x"00",	--9781
		x"41",	--9782
		x"00",	--9783
		x"89",	--9784
		x"40",	--9785
		x"d1",	--9786
		x"42",	--9787
		x"00",	--9788
		x"3c",	--9789
		x"d2",	--9790
		x"00",	--9791
		x"40",	--9792
		x"d1",	--9793
		x"41",	--9794
		x"f3",	--9795
		x"41",	--9796
		x"24",	--9797
		x"f0",	--9798
		x"ff",	--9799
		x"d3",	--9800
		x"3c",	--9801
		x"d3",	--9802
		x"4e",	--9803
		x"00",	--9804
		x"40",	--9805
		x"d1",	--9806
		x"d0",	--9807
		x"00",	--9808
		x"00",	--9809
		x"40",	--9810
		x"d1",	--9811
		x"40",	--9812
		x"00",	--9813
		x"00",	--9814
		x"40",	--9815
		x"d1",	--9816
		x"90",	--9817
		x"00",	--9818
		x"00",	--9819
		x"20",	--9820
		x"40",	--9821
		x"d1",	--9822
		x"40",	--9823
		x"00",	--9824
		x"00",	--9825
		x"40",	--9826
		x"d1",	--9827
		x"93",	--9828
		x"00",	--9829
		x"24",	--9830
		x"40",	--9831
		x"d1",	--9832
		x"43",	--9833
		x"00",	--9834
		x"40",	--9835
		x"d1",	--9836
		x"45",	--9837
		x"53",	--9838
		x"45",	--9839
		x"93",	--9840
		x"38",	--9841
		x"4a",	--9842
		x"00",	--9843
		x"3c",	--9844
		x"93",	--9845
		x"00",	--9846
		x"24",	--9847
		x"40",	--9848
		x"d1",	--9849
		x"d0",	--9850
		x"00",	--9851
		x"00",	--9852
		x"e3",	--9853
		x"4a",	--9854
		x"00",	--9855
		x"53",	--9856
		x"00",	--9857
		x"4e",	--9858
		x"3c",	--9859
		x"93",	--9860
		x"00",	--9861
		x"20",	--9862
		x"93",	--9863
		x"00",	--9864
		x"20",	--9865
		x"41",	--9866
		x"f0",	--9867
		x"00",	--9868
		x"43",	--9869
		x"24",	--9870
		x"43",	--9871
		x"4e",	--9872
		x"11",	--9873
		x"43",	--9874
		x"10",	--9875
		x"41",	--9876
		x"f0",	--9877
		x"00",	--9878
		x"de",	--9879
		x"4a",	--9880
		x"00",	--9881
		x"40",	--9882
		x"d1",	--9883
		x"41",	--9884
		x"00",	--9885
		x"5a",	--9886
		x"4a",	--9887
		x"5c",	--9888
		x"5c",	--9889
		x"5c",	--9890
		x"4a",	--9891
		x"00",	--9892
		x"50",	--9893
		x"ff",	--9894
		x"00",	--9895
		x"11",	--9896
		x"5e",	--9897
		x"00",	--9898
		x"43",	--9899
		x"00",	--9900
		x"40",	--9901
		x"d1",	--9902
		x"45",	--9903
		x"53",	--9904
		x"45",	--9905
		x"93",	--9906
		x"00",	--9907
		x"20",	--9908
		x"93",	--9909
		x"00",	--9910
		x"27",	--9911
		x"4e",	--9912
		x"00",	--9913
		x"43",	--9914
		x"00",	--9915
		x"41",	--9916
		x"52",	--9917
		x"3c",	--9918
		x"45",	--9919
		x"53",	--9920
		x"45",	--9921
		x"93",	--9922
		x"00",	--9923
		x"24",	--9924
		x"d2",	--9925
		x"00",	--9926
		x"41",	--9927
		x"00",	--9928
		x"4f",	--9929
		x"00",	--9930
		x"3c",	--9931
		x"93",	--9932
		x"00",	--9933
		x"24",	--9934
		x"41",	--9935
		x"00",	--9936
		x"00",	--9937
		x"93",	--9938
		x"20",	--9939
		x"40",	--9940
		x"dc",	--9941
		x"12",	--9942
		x"00",	--9943
		x"12",	--9944
		x"00",	--9945
		x"41",	--9946
		x"00",	--9947
		x"41",	--9948
		x"00",	--9949
		x"12",	--9950
		x"c9",	--9951
		x"52",	--9952
		x"5f",	--9953
		x"00",	--9954
		x"47",	--9955
		x"40",	--9956
		x"d1",	--9957
		x"45",	--9958
		x"53",	--9959
		x"45",	--9960
		x"49",	--9961
		x"00",	--9962
		x"43",	--9963
		x"93",	--9964
		x"20",	--9965
		x"43",	--9966
		x"5e",	--9967
		x"5e",	--9968
		x"5e",	--9969
		x"41",	--9970
		x"f0",	--9971
		x"ff",	--9972
		x"de",	--9973
		x"4a",	--9974
		x"00",	--9975
		x"47",	--9976
		x"40",	--9977
		x"00",	--9978
		x"00",	--9979
		x"3c",	--9980
		x"d3",	--9981
		x"00",	--9982
		x"3c",	--9983
		x"d2",	--9984
		x"00",	--9985
		x"40",	--9986
		x"00",	--9987
		x"00",	--9988
		x"3c",	--9989
		x"40",	--9990
		x"00",	--9991
		x"00",	--9992
		x"41",	--9993
		x"b3",	--9994
		x"24",	--9995
		x"45",	--9996
		x"52",	--9997
		x"45",	--9998
		x"45",	--9999
		x"00",	--10000
		x"45",	--10001
		x"00",	--10002
		x"45",	--10003
		x"00",	--10004
		x"48",	--10005
		x"00",	--10006
		x"47",	--10007
		x"00",	--10008
		x"46",	--10009
		x"00",	--10010
		x"4b",	--10011
		x"00",	--10012
		x"43",	--10013
		x"00",	--10014
		x"93",	--10015
		x"20",	--10016
		x"93",	--10017
		x"20",	--10018
		x"93",	--10019
		x"20",	--10020
		x"93",	--10021
		x"24",	--10022
		x"43",	--10023
		x"00",	--10024
		x"5b",	--10025
		x"43",	--10026
		x"6b",	--10027
		x"4b",	--10028
		x"00",	--10029
		x"4c",	--10030
		x"3c",	--10031
		x"f3",	--10032
		x"45",	--10033
		x"24",	--10034
		x"52",	--10035
		x"45",	--10036
		x"45",	--10037
		x"00",	--10038
		x"48",	--10039
		x"00",	--10040
		x"4b",	--10041
		x"00",	--10042
		x"43",	--10043
		x"00",	--10044
		x"93",	--10045
		x"20",	--10046
		x"3c",	--10047
		x"53",	--10048
		x"45",	--10049
		x"4b",	--10050
		x"00",	--10051
		x"43",	--10052
		x"00",	--10053
		x"93",	--10054
		x"24",	--10055
		x"43",	--10056
		x"00",	--10057
		x"5b",	--10058
		x"43",	--10059
		x"6b",	--10060
		x"4b",	--10061
		x"00",	--10062
		x"47",	--10063
		x"b2",	--10064
		x"00",	--10065
		x"24",	--10066
		x"93",	--10067
		x"00",	--10068
		x"20",	--10069
		x"41",	--10070
		x"90",	--10071
		x"00",	--10072
		x"00",	--10073
		x"20",	--10074
		x"d0",	--10075
		x"00",	--10076
		x"3c",	--10077
		x"92",	--10078
		x"00",	--10079
		x"20",	--10080
		x"d0",	--10081
		x"00",	--10082
		x"48",	--10083
		x"00",	--10084
		x"41",	--10085
		x"b2",	--10086
		x"24",	--10087
		x"93",	--10088
		x"00",	--10089
		x"24",	--10090
		x"40",	--10091
		x"00",	--10092
		x"00",	--10093
		x"b3",	--10094
		x"24",	--10095
		x"e3",	--10096
		x"00",	--10097
		x"e3",	--10098
		x"00",	--10099
		x"e3",	--10100
		x"00",	--10101
		x"e3",	--10102
		x"00",	--10103
		x"53",	--10104
		x"00",	--10105
		x"63",	--10106
		x"00",	--10107
		x"63",	--10108
		x"00",	--10109
		x"63",	--10110
		x"00",	--10111
		x"3c",	--10112
		x"b3",	--10113
		x"24",	--10114
		x"41",	--10115
		x"00",	--10116
		x"41",	--10117
		x"00",	--10118
		x"e3",	--10119
		x"e3",	--10120
		x"4a",	--10121
		x"4b",	--10122
		x"53",	--10123
		x"63",	--10124
		x"4e",	--10125
		x"00",	--10126
		x"4f",	--10127
		x"00",	--10128
		x"3c",	--10129
		x"41",	--10130
		x"00",	--10131
		x"e3",	--10132
		x"53",	--10133
		x"4a",	--10134
		x"00",	--10135
		x"43",	--10136
		x"00",	--10137
		x"b3",	--10138
		x"24",	--10139
		x"41",	--10140
		x"00",	--10141
		x"41",	--10142
		x"00",	--10143
		x"00",	--10144
		x"41",	--10145
		x"00",	--10146
		x"41",	--10147
		x"00",	--10148
		x"41",	--10149
		x"50",	--10150
		x"00",	--10151
		x"46",	--10152
		x"41",	--10153
		x"00",	--10154
		x"00",	--10155
		x"41",	--10156
		x"00",	--10157
		x"10",	--10158
		x"11",	--10159
		x"10",	--10160
		x"11",	--10161
		x"4b",	--10162
		x"00",	--10163
		x"4b",	--10164
		x"00",	--10165
		x"4b",	--10166
		x"00",	--10167
		x"12",	--10168
		x"00",	--10169
		x"12",	--10170
		x"00",	--10171
		x"12",	--10172
		x"00",	--10173
		x"12",	--10174
		x"00",	--10175
		x"49",	--10176
		x"41",	--10177
		x"00",	--10178
		x"48",	--10179
		x"44",	--10180
		x"12",	--10181
		x"d3",	--10182
		x"52",	--10183
		x"4c",	--10184
		x"90",	--10185
		x"00",	--10186
		x"34",	--10187
		x"50",	--10188
		x"00",	--10189
		x"4b",	--10190
		x"00",	--10191
		x"3c",	--10192
		x"4c",	--10193
		x"b3",	--10194
		x"00",	--10195
		x"24",	--10196
		x"40",	--10197
		x"00",	--10198
		x"3c",	--10199
		x"40",	--10200
		x"00",	--10201
		x"5b",	--10202
		x"4a",	--10203
		x"00",	--10204
		x"47",	--10205
		x"53",	--10206
		x"12",	--10207
		x"00",	--10208
		x"12",	--10209
		x"00",	--10210
		x"12",	--10211
		x"00",	--10212
		x"12",	--10213
		x"00",	--10214
		x"49",	--10215
		x"41",	--10216
		x"00",	--10217
		x"48",	--10218
		x"44",	--10219
		x"12",	--10220
		x"d3",	--10221
		x"52",	--10222
		x"4c",	--10223
		x"4d",	--10224
		x"00",	--10225
		x"4e",	--10226
		x"4f",	--10227
		x"53",	--10228
		x"93",	--10229
		x"23",	--10230
		x"93",	--10231
		x"23",	--10232
		x"93",	--10233
		x"23",	--10234
		x"93",	--10235
		x"23",	--10236
		x"43",	--10237
		x"00",	--10238
		x"43",	--10239
		x"00",	--10240
		x"43",	--10241
		x"00",	--10242
		x"43",	--10243
		x"00",	--10244
		x"3c",	--10245
		x"b3",	--10246
		x"24",	--10247
		x"41",	--10248
		x"00",	--10249
		x"41",	--10250
		x"00",	--10251
		x"41",	--10252
		x"50",	--10253
		x"00",	--10254
		x"41",	--10255
		x"00",	--10256
		x"10",	--10257
		x"11",	--10258
		x"10",	--10259
		x"11",	--10260
		x"41",	--10261
		x"00",	--10262
		x"49",	--10263
		x"44",	--10264
		x"47",	--10265
		x"12",	--10266
		x"d2",	--10267
		x"4e",	--10268
		x"90",	--10269
		x"00",	--10270
		x"34",	--10271
		x"50",	--10272
		x"00",	--10273
		x"4b",	--10274
		x"00",	--10275
		x"3c",	--10276
		x"4e",	--10277
		x"b3",	--10278
		x"00",	--10279
		x"24",	--10280
		x"40",	--10281
		x"00",	--10282
		x"3c",	--10283
		x"40",	--10284
		x"00",	--10285
		x"5b",	--10286
		x"4a",	--10287
		x"00",	--10288
		x"48",	--10289
		x"53",	--10290
		x"41",	--10291
		x"00",	--10292
		x"49",	--10293
		x"44",	--10294
		x"47",	--10295
		x"12",	--10296
		x"d2",	--10297
		x"4e",	--10298
		x"4f",	--10299
		x"53",	--10300
		x"93",	--10301
		x"23",	--10302
		x"93",	--10303
		x"23",	--10304
		x"43",	--10305
		x"00",	--10306
		x"43",	--10307
		x"00",	--10308
		x"3c",	--10309
		x"41",	--10310
		x"00",	--10311
		x"41",	--10312
		x"50",	--10313
		x"00",	--10314
		x"41",	--10315
		x"00",	--10316
		x"47",	--10317
		x"12",	--10318
		x"d2",	--10319
		x"4f",	--10320
		x"90",	--10321
		x"00",	--10322
		x"34",	--10323
		x"50",	--10324
		x"00",	--10325
		x"4d",	--10326
		x"00",	--10327
		x"3c",	--10328
		x"4f",	--10329
		x"b3",	--10330
		x"00",	--10331
		x"24",	--10332
		x"40",	--10333
		x"00",	--10334
		x"3c",	--10335
		x"40",	--10336
		x"00",	--10337
		x"5d",	--10338
		x"4c",	--10339
		x"00",	--10340
		x"48",	--10341
		x"53",	--10342
		x"41",	--10343
		x"00",	--10344
		x"47",	--10345
		x"12",	--10346
		x"d2",	--10347
		x"4f",	--10348
		x"53",	--10349
		x"93",	--10350
		x"23",	--10351
		x"43",	--10352
		x"00",	--10353
		x"90",	--10354
		x"00",	--10355
		x"00",	--10356
		x"24",	--10357
		x"43",	--10358
		x"00",	--10359
		x"93",	--10360
		x"00",	--10361
		x"24",	--10362
		x"41",	--10363
		x"50",	--10364
		x"00",	--10365
		x"4f",	--10366
		x"00",	--10367
		x"41",	--10368
		x"00",	--10369
		x"10",	--10370
		x"11",	--10371
		x"10",	--10372
		x"11",	--10373
		x"4a",	--10374
		x"00",	--10375
		x"46",	--10376
		x"00",	--10377
		x"46",	--10378
		x"10",	--10379
		x"11",	--10380
		x"10",	--10381
		x"11",	--10382
		x"4a",	--10383
		x"00",	--10384
		x"41",	--10385
		x"00",	--10386
		x"41",	--10387
		x"00",	--10388
		x"81",	--10389
		x"00",	--10390
		x"71",	--10391
		x"00",	--10392
		x"83",	--10393
		x"91",	--10394
		x"00",	--10395
		x"2c",	--10396
		x"d3",	--10397
		x"00",	--10398
		x"41",	--10399
		x"00",	--10400
		x"8c",	--10401
		x"4e",	--10402
		x"00",	--10403
		x"3c",	--10404
		x"93",	--10405
		x"00",	--10406
		x"24",	--10407
		x"41",	--10408
		x"00",	--10409
		x"00",	--10410
		x"12",	--10411
		x"00",	--10412
		x"12",	--10413
		x"00",	--10414
		x"41",	--10415
		x"00",	--10416
		x"46",	--10417
		x"53",	--10418
		x"41",	--10419
		x"00",	--10420
		x"12",	--10421
		x"c9",	--10422
		x"52",	--10423
		x"5f",	--10424
		x"00",	--10425
		x"3c",	--10426
		x"49",	--10427
		x"11",	--10428
		x"12",	--10429
		x"00",	--10430
		x"49",	--10431
		x"58",	--10432
		x"91",	--10433
		x"00",	--10434
		x"2b",	--10435
		x"49",	--10436
		x"00",	--10437
		x"4e",	--10438
		x"00",	--10439
		x"43",	--10440
		x"3c",	--10441
		x"41",	--10442
		x"00",	--10443
		x"00",	--10444
		x"43",	--10445
		x"00",	--10446
		x"43",	--10447
		x"00",	--10448
		x"3c",	--10449
		x"4e",	--10450
		x"43",	--10451
		x"00",	--10452
		x"43",	--10453
		x"00",	--10454
		x"43",	--10455
		x"41",	--10456
		x"00",	--10457
		x"46",	--10458
		x"93",	--10459
		x"24",	--10460
		x"40",	--10461
		x"cb",	--10462
		x"41",	--10463
		x"00",	--10464
		x"50",	--10465
		x"00",	--10466
		x"41",	--10467
		x"41",	--10468
		x"41",	--10469
		x"41",	--10470
		x"41",	--10471
		x"41",	--10472
		x"41",	--10473
		x"41",	--10474
		x"41",	--10475
		x"43",	--10476
		x"93",	--10477
		x"34",	--10478
		x"40",	--10479
		x"00",	--10480
		x"e3",	--10481
		x"53",	--10482
		x"93",	--10483
		x"34",	--10484
		x"e3",	--10485
		x"e3",	--10486
		x"53",	--10487
		x"12",	--10488
		x"12",	--10489
		x"d2",	--10490
		x"41",	--10491
		x"b3",	--10492
		x"24",	--10493
		x"e3",	--10494
		x"53",	--10495
		x"b3",	--10496
		x"24",	--10497
		x"e3",	--10498
		x"53",	--10499
		x"41",	--10500
		x"12",	--10501
		x"d1",	--10502
		x"4e",	--10503
		x"41",	--10504
		x"12",	--10505
		x"12",	--10506
		x"12",	--10507
		x"40",	--10508
		x"00",	--10509
		x"4c",	--10510
		x"4d",	--10511
		x"43",	--10512
		x"43",	--10513
		x"5e",	--10514
		x"6f",	--10515
		x"6c",	--10516
		x"6d",	--10517
		x"9b",	--10518
		x"28",	--10519
		x"20",	--10520
		x"9a",	--10521
		x"28",	--10522
		x"8a",	--10523
		x"7b",	--10524
		x"d3",	--10525
		x"83",	--10526
		x"23",	--10527
		x"41",	--10528
		x"41",	--10529
		x"41",	--10530
		x"41",	--10531
		x"12",	--10532
		x"d2",	--10533
		x"4c",	--10534
		x"4d",	--10535
		x"41",	--10536
		x"12",	--10537
		x"43",	--10538
		x"93",	--10539
		x"34",	--10540
		x"40",	--10541
		x"00",	--10542
		x"e3",	--10543
		x"e3",	--10544
		x"53",	--10545
		x"63",	--10546
		x"93",	--10547
		x"34",	--10548
		x"e3",	--10549
		x"e3",	--10550
		x"e3",	--10551
		x"53",	--10552
		x"63",	--10553
		x"12",	--10554
		x"d2",	--10555
		x"b3",	--10556
		x"24",	--10557
		x"e3",	--10558
		x"e3",	--10559
		x"53",	--10560
		x"63",	--10561
		x"b3",	--10562
		x"24",	--10563
		x"e3",	--10564
		x"e3",	--10565
		x"53",	--10566
		x"63",	--10567
		x"41",	--10568
		x"41",	--10569
		x"12",	--10570
		x"d2",	--10571
		x"4c",	--10572
		x"4d",	--10573
		x"41",	--10574
		x"40",	--10575
		x"00",	--10576
		x"4e",	--10577
		x"43",	--10578
		x"5f",	--10579
		x"6e",	--10580
		x"9d",	--10581
		x"28",	--10582
		x"8d",	--10583
		x"d3",	--10584
		x"83",	--10585
		x"23",	--10586
		x"41",	--10587
		x"12",	--10588
		x"d2",	--10589
		x"4e",	--10590
		x"41",	--10591
		x"12",	--10592
		x"12",	--10593
		x"12",	--10594
		x"12",	--10595
		x"12",	--10596
		x"00",	--10597
		x"48",	--10598
		x"49",	--10599
		x"4a",	--10600
		x"4b",	--10601
		x"43",	--10602
		x"43",	--10603
		x"43",	--10604
		x"43",	--10605
		x"5c",	--10606
		x"6d",	--10607
		x"6e",	--10608
		x"6f",	--10609
		x"68",	--10610
		x"69",	--10611
		x"6a",	--10612
		x"6b",	--10613
		x"97",	--10614
		x"28",	--10615
		x"20",	--10616
		x"96",	--10617
		x"28",	--10618
		x"20",	--10619
		x"95",	--10620
		x"28",	--10621
		x"20",	--10622
		x"94",	--10623
		x"28",	--10624
		x"84",	--10625
		x"75",	--10626
		x"76",	--10627
		x"77",	--10628
		x"d3",	--10629
		x"83",	--10630
		x"00",	--10631
		x"23",	--10632
		x"53",	--10633
		x"41",	--10634
		x"41",	--10635
		x"41",	--10636
		x"41",	--10637
		x"41",	--10638
		x"12",	--10639
		x"12",	--10640
		x"12",	--10641
		x"12",	--10642
		x"41",	--10643
		x"00",	--10644
		x"41",	--10645
		x"00",	--10646
		x"41",	--10647
		x"00",	--10648
		x"41",	--10649
		x"00",	--10650
		x"12",	--10651
		x"d2",	--10652
		x"41",	--10653
		x"41",	--10654
		x"41",	--10655
		x"41",	--10656
		x"41",	--10657
		x"12",	--10658
		x"12",	--10659
		x"12",	--10660
		x"12",	--10661
		x"41",	--10662
		x"00",	--10663
		x"41",	--10664
		x"00",	--10665
		x"41",	--10666
		x"00",	--10667
		x"41",	--10668
		x"00",	--10669
		x"12",	--10670
		x"d2",	--10671
		x"48",	--10672
		x"49",	--10673
		x"4a",	--10674
		x"4b",	--10675
		x"41",	--10676
		x"41",	--10677
		x"41",	--10678
		x"41",	--10679
		x"41",	--10680
		x"12",	--10681
		x"12",	--10682
		x"12",	--10683
		x"12",	--10684
		x"12",	--10685
		x"41",	--10686
		x"00",	--10687
		x"41",	--10688
		x"00",	--10689
		x"41",	--10690
		x"00",	--10691
		x"41",	--10692
		x"00",	--10693
		x"12",	--10694
		x"d2",	--10695
		x"41",	--10696
		x"00",	--10697
		x"48",	--10698
		x"00",	--10699
		x"49",	--10700
		x"00",	--10701
		x"4a",	--10702
		x"00",	--10703
		x"4b",	--10704
		x"00",	--10705
		x"41",	--10706
		x"41",	--10707
		x"41",	--10708
		x"41",	--10709
		x"41",	--10710
		x"41",	--10711
		x"13",	--10712
		x"d0",	--10713
		x"00",	--10714
		x"3f",	--10715
		x"3d",	--10716
		x"64",	--10717
		x"79",	--10718
		x"25",	--10719
		x"20",	--10720
		x"3d",	--10721
		x"64",	--10722
		x"25",	--10723
		x"0d",	--10724
		x"00",	--10725
		x"64",	--10726
		x"00",	--10727
		x"0a",	--10728
		x"00",	--10729
		x"85",	--10730
		x"85",	--10731
		x"85",	--10732
		x"85",	--10733
		x"85",	--10734
		x"85",	--10735
		x"85",	--10736
		x"85",	--10737
		x"0a",	--10738
		x"3d",	--10739
		x"3d",	--10740
		x"3d",	--10741
		x"4d",	--10742
		x"72",	--10743
		x"65",	--10744
		x"20",	--10745
		x"43",	--10746
		x"20",	--10747
		x"3d",	--10748
		x"3d",	--10749
		x"3d",	--10750
		x"0a",	--10751
		x"69",	--10752
		x"74",	--10753
		x"72",	--10754
		x"63",	--10755
		x"69",	--10756
		x"65",	--10757
		x"6d",	--10758
		x"64",	--10759
		x"00",	--10760
		x"72",	--10761
		x"74",	--10762
		x"00",	--10763
		x"65",	--10764
		x"64",	--10765
		x"62",	--10766
		x"7a",	--10767
		x"65",	--10768
		x"00",	--10769
		x"77",	--10770
		x"00",	--10771
		x"6e",	--10772
		x"6f",	--10773
		x"65",	--10774
		x"00",	--10775
		x"70",	--10776
		x"65",	--10777
		x"20",	--10778
		x"6f",	--10779
		x"74",	--10780
		x"6f",	--10781
		x"6c",	--10782
		x"72",	--10783
		x"6f",	--10784
		x"6f",	--10785
		x"65",	--10786
		x"72",	--10787
		x"00",	--10788
		x"70",	--10789
		x"65",	--10790
		x"20",	--10791
		x"6f",	--10792
		x"66",	--10793
		x"67",	--10794
		x"72",	--10795
		x"74",	--10796
		x"6f",	--10797
		x"00",	--10798
		x"62",	--10799
		x"74",	--10800
		x"63",	--10801
		x"65",	--10802
		x"61",	--10803
		x"6f",	--10804
		x"64",	--10805
		x"6e",	--10806
		x"65",	--10807
		x"72",	--10808
		x"61",	--10809
		x"00",	--10810
		x"6f",	--10811
		x"74",	--10812
		x"6f",	--10813
		x"64",	--10814
		x"72",	--10815
		x"0d",	--10816
		x"00",	--10817
		x"20",	--10818
		x"00",	--10819
		x"63",	--10820
		x"55",	--10821
		x"0d",	--10822
		x"00",	--10823
		x"4f",	--10824
		x"4e",	--10825
		x"0a",	--10826
		x"52",	--10827
		x"47",	--10828
		x"54",	--10829
		x"0a",	--10830
		x"4c",	--10831
		x"46",	--10832
		x"0d",	--10833
		x"00",	--10834
		x"74",	--10835
		x"70",	--10836
		x"0a",	--10837
		x"63",	--10838
		x"72",	--10839
		x"65",	--10840
		x"74",	--10841
		x"75",	--10842
		x"61",	--10843
		x"65",	--10844
		x"0d",	--10845
		x"00",	--10846
		x"25",	--10847
		x"20",	--10848
		x"6f",	--10849
		x"20",	--10850
		x"45",	--10851
		x"54",	--10852
		x"52",	--10853
		x"47",	--10854
		x"54",	--10855
		x"3c",	--10856
		x"49",	--10857
		x"45",	--10858
		x"55",	--10859
		x"3e",	--10860
		x"0a",	--10861
		x"25",	--10862
		x"20",	--10863
		x"64",	--10864
		x"0a",	--10865
		x"4e",	--10866
		x"74",	--10867
		x"69",	--10868
		x"70",	--10869
		x"65",	--10870
		x"65",	--10871
		x"74",	--10872
		x"64",	--10873
		x"59",	--10874
		x"74",	--10875
		x"0a",	--10876
		x"57",	--10877
		x"69",	--10878
		x"69",	--10879
		x"67",	--10880
		x"66",	--10881
		x"72",	--10882
		x"61",	--10883
		x"6e",	--10884
		x"77",	--10885
		x"2e",	--10886
		x"69",	--10887
		x"20",	--10888
		x"69",	--10889
		x"65",	--10890
		x"0a",	--10891
		x"57",	--10892
		x"20",	--10893
		x"68",	--10894
		x"75",	--10895
		x"64",	--10896
		x"6e",	--10897
		x"74",	--10898
		x"73",	--10899
		x"65",	--10900
		x"74",	--10901
		x"61",	--10902
		x"0d",	--10903
		x"00",	--10904
		x"63",	--10905
		x"69",	--10906
		x"20",	--10907
		x"6f",	--10908
		x"20",	--10909
		x"20",	--10910
		x"75",	--10911
		x"62",	--10912
		x"72",	--10913
		x"0a",	--10914
		x"53",	--10915
		x"6f",	--10916
		x"0d",	--10917
		x"00",	--10918
		x"72",	--10919
		x"6f",	--10920
		x"3a",	--10921
		x"6d",	--10922
		x"73",	--10923
		x"69",	--10924
		x"67",	--10925
		x"61",	--10926
		x"67",	--10927
		x"6d",	--10928
		x"6e",	--10929
		x"0d",	--10930
		x"00",	--10931
		x"6f",	--10932
		x"72",	--10933
		x"63",	--10934
		x"20",	--10935
		x"73",	--10936
		x"67",	--10937
		x"3a",	--10938
		x"0a",	--10939
		x"09",	--10940
		x"73",	--10941
		x"4c",	--10942
		x"46",	--10943
		x"20",	--10944
		x"49",	--10945
		x"48",	--10946
		x"20",	--10947
		x"54",	--10948
		x"4d",	--10949
		x"4f",	--10950
		x"54",	--10951
		x"0d",	--10952
		x"00",	--10953
		x"64",	--10954
		x"25",	--10955
		x"0d",	--10956
		x"00",	--10957
		x"6c",	--10958
		x"20",	--10959
		x"6c",	--10960
		x"00",	--10961
		x"73",	--10962
		x"0a",	--10963
		x"25",	--10964
		x"20",	--10965
		x"64",	--10966
		x"0a",	--10967
		x"25",	--10968
		x"20",	--10969
		x"0d",	--10970
		x"00",	--10971
		x"6f",	--10972
		x"62",	--10973
		x"68",	--10974
		x"6e",	--10975
		x"20",	--10976
		x"65",	--10977
		x"62",	--10978
		x"74",	--10979
		x"49",	--10980
		x"64",	--10981
		x"6e",	--10982
		x"74",	--10983
		x"67",	--10984
		x"76",	--10985
		x"20",	--10986
		x"20",	--10987
		x"68",	--10988
		x"74",	--10989
		x"0d",	--10990
		x"00",	--10991
		x"6f",	--10992
		x"69",	--10993
		x"20",	--10994
		x"72",	--10995
		x"6e",	--10996
		x"0d",	--10997
		x"00",	--10998
		x"6f",	--10999
		x"6f",	--11000
		x"20",	--11001
		x"68",	--11002
		x"20",	--11003
		x"69",	--11004
		x"68",	--11005
		x"0d",	--11006
		x"00",	--11007
		x"6f",	--11008
		x"6f",	--11009
		x"20",	--11010
		x"68",	--11011
		x"20",	--11012
		x"65",	--11013
		x"74",	--11014
		x"0a",	--11015
		x"25",	--11016
		x"0d",	--11017
		x"00",	--11018
		x"74",	--11019
		x"70",	--11020
		x"0a",	--11021
		x"66",	--11022
		x"6f",	--11023
		x"74",	--11024
		x"72",	--11025
		x"74",	--11026
		x"74",	--11027
		x"6f",	--11028
		x"0d",	--11029
		x"00",	--11030
		x"65",	--11031
		x"74",	--11032
		x"72",	--11033
		x"74",	--11034
		x"74",	--11035
		x"6f",	--11036
		x"0d",	--11037
		x"00",	--11038
		x"69",	--11039
		x"68",	--11040
		x"3a",	--11041
		x"6f",	--11042
		x"61",	--11043
		x"69",	--11044
		x"6e",	--11045
		x"0a",	--11046
		x"52",	--11047
		x"61",	--11048
		x"69",	--11049
		x"67",	--11050
		x"61",	--11051
		x"74",	--11052
		x"76",	--11053
		x"74",	--11054
		x"64",	--11055
		x"0a",	--11056
		x"52",	--11057
		x"61",	--11058
		x"69",	--11059
		x"67",	--11060
		x"64",	--11061
		x"61",	--11062
		x"74",	--11063
		x"76",	--11064
		x"74",	--11065
		x"64",	--11066
		x"0a",	--11067
		x"77",	--11068
		x"69",	--11069
		x"65",	--11070
		x"0d",	--11071
		x"65",	--11072
		x"72",	--11073
		x"72",	--11074
		x"20",	--11075
		x"69",	--11076
		x"73",	--11077
		x"6e",	--11078
		x"20",	--11079
		x"72",	--11080
		x"75",	--11081
		x"65",	--11082
		x"74",	--11083
		x"0a",	--11084
		x"63",	--11085
		x"72",	--11086
		x"65",	--11087
		x"74",	--11088
		x"75",	--11089
		x"61",	--11090
		x"65",	--11091
		x"0d",	--11092
		x"00",	--11093
		x"25",	--11094
		x"20",	--11095
		x"45",	--11096
		x"49",	--11097
		x"54",	--11098
		x"52",	--11099
		x"56",	--11100
		x"4c",	--11101
		x"45",	--11102
		x"0a",	--11103
		x"72",	--11104
		x"25",	--11105
		x"20",	--11106
		x"3d",	--11107
		x"64",	--11108
		x"0a",	--11109
		x"09",	--11110
		x"73",	--11111
		x"52",	--11112
		x"47",	--11113
		x"53",	--11114
		x"45",	--11115
		x"0d",	--11116
		x"00",	--11117
		x"65",	--11118
		x"64",	--11119
		x"0d",	--11120
		x"25",	--11121
		x"20",	--11122
		x"73",	--11123
		x"0a",	--11124
		x"25",	--11125
		x"3a",	--11126
		x"6e",	--11127
		x"20",	--11128
		x"75",	--11129
		x"68",	--11130
		x"63",	--11131
		x"6d",	--11132
		x"61",	--11133
		x"64",	--11134
		x"0a",	--11135
		x"00",	--11136
		x"9c",	--11137
		x"9b",	--11138
		x"9b",	--11139
		x"9b",	--11140
		x"9b",	--11141
		x"9b",	--11142
		x"9b",	--11143
		x"9b",	--11144
		x"9b",	--11145
		x"9b",	--11146
		x"9b",	--11147
		x"9b",	--11148
		x"9b",	--11149
		x"9b",	--11150
		x"9b",	--11151
		x"9b",	--11152
		x"9b",	--11153
		x"9b",	--11154
		x"9b",	--11155
		x"9b",	--11156
		x"9b",	--11157
		x"9b",	--11158
		x"9b",	--11159
		x"9b",	--11160
		x"9b",	--11161
		x"9b",	--11162
		x"9b",	--11163
		x"9b",	--11164
		x"9b",	--11165
		x"9c",	--11166
		x"9b",	--11167
		x"9b",	--11168
		x"9b",	--11169
		x"9b",	--11170
		x"9b",	--11171
		x"9b",	--11172
		x"9b",	--11173
		x"9b",	--11174
		x"9b",	--11175
		x"9b",	--11176
		x"9b",	--11177
		x"9b",	--11178
		x"9b",	--11179
		x"9b",	--11180
		x"9b",	--11181
		x"9b",	--11182
		x"9b",	--11183
		x"9b",	--11184
		x"9b",	--11185
		x"9b",	--11186
		x"9b",	--11187
		x"9b",	--11188
		x"9b",	--11189
		x"9b",	--11190
		x"9b",	--11191
		x"9b",	--11192
		x"9b",	--11193
		x"9b",	--11194
		x"9b",	--11195
		x"9b",	--11196
		x"9b",	--11197
		x"9c",	--11198
		x"9c",	--11199
		x"9c",	--11200
		x"9b",	--11201
		x"9b",	--11202
		x"9b",	--11203
		x"9b",	--11204
		x"9b",	--11205
		x"9b",	--11206
		x"9b",	--11207
		x"9c",	--11208
		x"9b",	--11209
		x"9c",	--11210
		x"9b",	--11211
		x"9b",	--11212
		x"9b",	--11213
		x"9b",	--11214
		x"9c",	--11215
		x"9b",	--11216
		x"9b",	--11217
		x"9b",	--11218
		x"9b",	--11219
		x"9b",	--11220
		x"31",	--11221
		x"33",	--11222
		x"35",	--11223
		x"37",	--11224
		x"39",	--11225
		x"62",	--11226
		x"64",	--11227
		x"66",	--11228
		x"00",	--11229
		x"63",	--11230
		x"3e",	--11231
		x"0f",	--11232
		x"3f",	--11233
		x"98",	--11234
		x"3f",	--11235
		x"0f",	--11236
		x"3f",	--11237
		x"37",	--11238
		x"31",	--11239
		x"21",	--11240
		x"33",	--11241
		x"0f",	--11242
		x"33",	--11243
		x"21",	--11244
		x"33",	--11245
		x"0f",	--11246
		x"3f",	--11247
		x"0f",	--11248
		x"40",	--11249
		x"cb",	--11250
		x"40",	--11251
		x"0f",	--11252
		x"40",	--11253
		x"53",	--11254
		x"40",	--11255
		x"cb",	--11256
		x"41",	--11257
		x"ed",	--11258
		x"41",	--11259
		x"0f",	--11260
		x"41",	--11261
		x"31",	--11262
		x"41",	--11263
		x"53",	--11264
		x"41",	--11265
		x"3a",	--11266
		x"41",	--11267
		x"cb",	--11268
		x"41",	--11269
		x"5c",	--11270
		x"41",	--11271
		x"ed",	--11272
		x"41",	--11273
		x"7e",	--11274
		x"41",	--11275
		x"0f",	--11276
		x"41",	--11277
		x"a0",	--11278
		x"41",	--11279
		x"31",	--11280
		x"41",	--11281
		x"c2",	--11282
		x"41",	--11283
		x"53",	--11284
		x"41",	--11285
		x"f2",	--11286
		x"42",	--11287
		x"3a",	--11288
		x"42",	--11289
		x"83",	--11290
		x"42",	--11291
		x"cb",	--11292
		x"42",	--11293
		x"14",	--11294
		x"42",	--11295
		x"5c",	--11296
		x"42",	--11297
		x"a5",	--11298
		x"42",	--11299
		x"ed",	--11300
		x"42",	--11301
		x"36",	--11302
		x"42",	--11303
		x"7e",	--11304
		x"42",	--11305
		x"c7",	--11306
		x"42",	--11307
		x"0f",	--11308
		x"42",	--11309
		x"00",	--11310
		x"00",	--11311
		x"00",	--11312
		x"00",	--11313
		x"00",	--11314
		x"00",	--11315
		x"00",	--11316
		x"00",	--11317
		x"00",	--11318
		x"00",	--11319
		x"00",	--11320
		x"00",	--11321
		x"00",	--11322
		x"00",	--11323
		x"00",	--11324
		x"00",	--11325
		x"00",	--11326
		x"00",	--11327
		x"00",	--11328
		x"00",	--11329
		x"00",	--11330
		x"00",	--11331
		x"00",	--11332
		x"00",	--11333
		x"00",	--11334
		x"00",	--11335
		x"00",	--11336
		x"00",	--11337
		x"00",	--11338
		x"00",	--11339
		x"00",	--11340
		x"00",	--11341
		x"00",	--11342
		x"00",	--11343
		x"00",	--11344
		x"00",	--11345
		x"00",	--11346
		x"00",	--11347
		x"00",	--11348
		x"00",	--11349
		x"00",	--11350
		x"00",	--11351
		x"00",	--11352
		x"00",	--11353
		x"00",	--11354
		x"00",	--11355
		x"00",	--11356
		x"00",	--11357
		x"00",	--11358
		x"00",	--11359
		x"00",	--11360
		x"00",	--11361
		x"00",	--11362
		x"00",	--11363
		x"00",	--11364
		x"00",	--11365
		x"00",	--11366
		x"00",	--11367
		x"00",	--11368
		x"00",	--11369
		x"00",	--11370
		x"00",	--11371
		x"00",	--11372
		x"00",	--11373
		x"00",	--11374
		x"00",	--11375
		x"00",	--11376
		x"00",	--11377
		x"00",	--11378
		x"00",	--11379
		x"00",	--11380
		x"00",	--11381
		x"00",	--11382
		x"00",	--11383
		x"00",	--11384
		x"00",	--11385
		x"00",	--11386
		x"00",	--11387
		x"00",	--11388
		x"00",	--11389
		x"00",	--11390
		x"00",	--11391
		x"00",	--11392
		x"00",	--11393
		x"00",	--11394
		x"00",	--11395
		x"00",	--11396
		x"00",	--11397
		x"00",	--11398
		x"00",	--11399
		x"00",	--11400
		x"00",	--11401
		x"00",	--11402
		x"00",	--11403
		x"00",	--11404
		x"00",	--11405
		x"00",	--11406
		x"00",	--11407
		x"00",	--11408
		x"00",	--11409
		x"00",	--11410
		x"00",	--11411
		x"00",	--11412
		x"00",	--11413
		x"00",	--11414
		x"00",	--11415
		x"00",	--11416
		x"00",	--11417
		x"00",	--11418
		x"00",	--11419
		x"00",	--11420
		x"00",	--11421
		x"00",	--11422
		x"00",	--11423
		x"00",	--11424
		x"00",	--11425
		x"00",	--11426
		x"00",	--11427
		x"00",	--11428
		x"00",	--11429
		x"00",	--11430
		x"00",	--11431
		x"00",	--11432
		x"00",	--11433
		x"00",	--11434
		x"00",	--11435
		x"00",	--11436
		x"00",	--11437
		x"00",	--11438
		x"00",	--11439
		x"00",	--11440
		x"00",	--11441
		x"00",	--11442
		x"00",	--11443
		x"00",	--11444
		x"00",	--11445
		x"00",	--11446
		x"00",	--11447
		x"00",	--11448
		x"00",	--11449
		x"00",	--11450
		x"00",	--11451
		x"00",	--11452
		x"00",	--11453
		x"00",	--11454
		x"00",	--11455
		x"00",	--11456
		x"00",	--11457
		x"00",	--11458
		x"00",	--11459
		x"00",	--11460
		x"00",	--11461
		x"00",	--11462
		x"00",	--11463
		x"00",	--11464
		x"00",	--11465
		x"00",	--11466
		x"00",	--11467
		x"00",	--11468
		x"00",	--11469
		x"00",	--11470
		x"00",	--11471
		x"00",	--11472
		x"00",	--11473
		x"00",	--11474
		x"00",	--11475
		x"00",	--11476
		x"00",	--11477
		x"00",	--11478
		x"00",	--11479
		x"00",	--11480
		x"00",	--11481
		x"00",	--11482
		x"00",	--11483
		x"00",	--11484
		x"00",	--11485
		x"00",	--11486
		x"00",	--11487
		x"00",	--11488
		x"00",	--11489
		x"00",	--11490
		x"00",	--11491
		x"00",	--11492
		x"00",	--11493
		x"00",	--11494
		x"00",	--11495
		x"00",	--11496
		x"00",	--11497
		x"00",	--11498
		x"00",	--11499
		x"00",	--11500
		x"00",	--11501
		x"00",	--11502
		x"00",	--11503
		x"00",	--11504
		x"00",	--11505
		x"00",	--11506
		x"00",	--11507
		x"00",	--11508
		x"00",	--11509
		x"00",	--11510
		x"00",	--11511
		x"00",	--11512
		x"00",	--11513
		x"00",	--11514
		x"00",	--11515
		x"00",	--11516
		x"00",	--11517
		x"00",	--11518
		x"00",	--11519
		x"00",	--11520
		x"00",	--11521
		x"00",	--11522
		x"00",	--11523
		x"00",	--11524
		x"00",	--11525
		x"00",	--11526
		x"00",	--11527
		x"00",	--11528
		x"00",	--11529
		x"00",	--11530
		x"00",	--11531
		x"00",	--11532
		x"00",	--11533
		x"00",	--11534
		x"00",	--11535
		x"00",	--11536
		x"00",	--11537
		x"00",	--11538
		x"00",	--11539
		x"00",	--11540
		x"00",	--11541
		x"00",	--11542
		x"00",	--11543
		x"00",	--11544
		x"00",	--11545
		x"00",	--11546
		x"00",	--11547
		x"00",	--11548
		x"00",	--11549
		x"00",	--11550
		x"00",	--11551
		x"00",	--11552
		x"00",	--11553
		x"00",	--11554
		x"00",	--11555
		x"00",	--11556
		x"00",	--11557
		x"00",	--11558
		x"00",	--11559
		x"00",	--11560
		x"00",	--11561
		x"00",	--11562
		x"00",	--11563
		x"00",	--11564
		x"00",	--11565
		x"00",	--11566
		x"00",	--11567
		x"00",	--11568
		x"00",	--11569
		x"00",	--11570
		x"00",	--11571
		x"00",	--11572
		x"00",	--11573
		x"00",	--11574
		x"00",	--11575
		x"00",	--11576
		x"00",	--11577
		x"00",	--11578
		x"00",	--11579
		x"00",	--11580
		x"00",	--11581
		x"00",	--11582
		x"00",	--11583
		x"00",	--11584
		x"00",	--11585
		x"00",	--11586
		x"00",	--11587
		x"00",	--11588
		x"00",	--11589
		x"00",	--11590
		x"00",	--11591
		x"00",	--11592
		x"00",	--11593
		x"00",	--11594
		x"00",	--11595
		x"00",	--11596
		x"00",	--11597
		x"00",	--11598
		x"00",	--11599
		x"00",	--11600
		x"00",	--11601
		x"00",	--11602
		x"00",	--11603
		x"00",	--11604
		x"00",	--11605
		x"00",	--11606
		x"00",	--11607
		x"00",	--11608
		x"00",	--11609
		x"00",	--11610
		x"00",	--11611
		x"00",	--11612
		x"00",	--11613
		x"00",	--11614
		x"00",	--11615
		x"00",	--11616
		x"00",	--11617
		x"00",	--11618
		x"00",	--11619
		x"00",	--11620
		x"00",	--11621
		x"00",	--11622
		x"00",	--11623
		x"00",	--11624
		x"00",	--11625
		x"00",	--11626
		x"00",	--11627
		x"00",	--11628
		x"00",	--11629
		x"00",	--11630
		x"00",	--11631
		x"00",	--11632
		x"00",	--11633
		x"00",	--11634
		x"00",	--11635
		x"00",	--11636
		x"00",	--11637
		x"00",	--11638
		x"00",	--11639
		x"00",	--11640
		x"00",	--11641
		x"00",	--11642
		x"00",	--11643
		x"00",	--11644
		x"00",	--11645
		x"00",	--11646
		x"00",	--11647
		x"00",	--11648
		x"00",	--11649
		x"00",	--11650
		x"00",	--11651
		x"00",	--11652
		x"00",	--11653
		x"00",	--11654
		x"00",	--11655
		x"00",	--11656
		x"00",	--11657
		x"00",	--11658
		x"00",	--11659
		x"00",	--11660
		x"00",	--11661
		x"00",	--11662
		x"00",	--11663
		x"00",	--11664
		x"00",	--11665
		x"00",	--11666
		x"00",	--11667
		x"00",	--11668
		x"00",	--11669
		x"00",	--11670
		x"00",	--11671
		x"00",	--11672
		x"00",	--11673
		x"00",	--11674
		x"00",	--11675
		x"00",	--11676
		x"00",	--11677
		x"00",	--11678
		x"00",	--11679
		x"00",	--11680
		x"00",	--11681
		x"00",	--11682
		x"00",	--11683
		x"00",	--11684
		x"00",	--11685
		x"00",	--11686
		x"00",	--11687
		x"00",	--11688
		x"00",	--11689
		x"00",	--11690
		x"00",	--11691
		x"00",	--11692
		x"00",	--11693
		x"00",	--11694
		x"00",	--11695
		x"00",	--11696
		x"00",	--11697
		x"00",	--11698
		x"00",	--11699
		x"00",	--11700
		x"00",	--11701
		x"00",	--11702
		x"00",	--11703
		x"00",	--11704
		x"00",	--11705
		x"00",	--11706
		x"00",	--11707
		x"00",	--11708
		x"00",	--11709
		x"3f",	--11710
		x"00",	--11711
		x"39",	--11712
		x"00",	--11713
		x"37",	--11714
		x"00",	--11715
		x"33",	--11716
		x"00",	--11717
		x"2e",	--11718
		x"00",	--11719
		x"2b",	--11720
		x"00",	--11721
		x"27",	--11722
		x"00",	--11723
		x"22",	--11724
		x"00",	--11725
		x"1f",	--11726
		x"00",	--11727
		x"1b",	--11728
		x"00",	--11729
		x"17",	--11730
		x"00",	--11731
		x"00",	--11732
		x"00",	--11733
		x"00",	--11734
		x"01",	--11735
		x"02",	--11736
		x"03",	--11737
		x"03",	--11738
		x"04",	--11739
		x"04",	--11740
		x"04",	--11741
		x"04",	--11742
		x"05",	--11743
		x"05",	--11744
		x"05",	--11745
		x"05",	--11746
		x"05",	--11747
		x"05",	--11748
		x"05",	--11749
		x"05",	--11750
		x"06",	--11751
		x"06",	--11752
		x"06",	--11753
		x"06",	--11754
		x"06",	--11755
		x"06",	--11756
		x"06",	--11757
		x"06",	--11758
		x"06",	--11759
		x"06",	--11760
		x"06",	--11761
		x"06",	--11762
		x"06",	--11763
		x"06",	--11764
		x"06",	--11765
		x"06",	--11766
		x"07",	--11767
		x"07",	--11768
		x"07",	--11769
		x"07",	--11770
		x"07",	--11771
		x"07",	--11772
		x"07",	--11773
		x"07",	--11774
		x"07",	--11775
		x"07",	--11776
		x"07",	--11777
		x"07",	--11778
		x"07",	--11779
		x"07",	--11780
		x"07",	--11781
		x"07",	--11782
		x"07",	--11783
		x"07",	--11784
		x"07",	--11785
		x"07",	--11786
		x"07",	--11787
		x"07",	--11788
		x"07",	--11789
		x"07",	--11790
		x"07",	--11791
		x"07",	--11792
		x"07",	--11793
		x"07",	--11794
		x"07",	--11795
		x"07",	--11796
		x"07",	--11797
		x"07",	--11798
		x"08",	--11799
		x"08",	--11800
		x"08",	--11801
		x"08",	--11802
		x"08",	--11803
		x"08",	--11804
		x"08",	--11805
		x"08",	--11806
		x"08",	--11807
		x"08",	--11808
		x"08",	--11809
		x"08",	--11810
		x"08",	--11811
		x"08",	--11812
		x"08",	--11813
		x"08",	--11814
		x"08",	--11815
		x"08",	--11816
		x"08",	--11817
		x"08",	--11818
		x"08",	--11819
		x"08",	--11820
		x"08",	--11821
		x"08",	--11822
		x"08",	--11823
		x"08",	--11824
		x"08",	--11825
		x"08",	--11826
		x"08",	--11827
		x"08",	--11828
		x"08",	--11829
		x"08",	--11830
		x"08",	--11831
		x"08",	--11832
		x"08",	--11833
		x"08",	--11834
		x"08",	--11835
		x"08",	--11836
		x"08",	--11837
		x"08",	--11838
		x"08",	--11839
		x"08",	--11840
		x"08",	--11841
		x"08",	--11842
		x"08",	--11843
		x"08",	--11844
		x"08",	--11845
		x"08",	--11846
		x"08",	--11847
		x"08",	--11848
		x"08",	--11849
		x"08",	--11850
		x"08",	--11851
		x"08",	--11852
		x"08",	--11853
		x"08",	--11854
		x"08",	--11855
		x"08",	--11856
		x"08",	--11857
		x"08",	--11858
		x"08",	--11859
		x"08",	--11860
		x"08",	--11861
		x"08",	--11862
		x"6e",	--11863
		x"6c",	--11864
		x"29",	--11865
		x"00",	--11866
		x"ff",	--11867
		x"ff",	--11868
		x"ff",	--11869
		x"ff",	--11870
		x"01",	--11871
		x"01",	--11872
		x"01",	--11873
		x"01",	--11874
		x"01",	--11875
		x"65",	--11876
		x"70",	--11877
		x"00",	--11878
		x"ff",	--11879
		x"ff",	--11880
		x"ff",	--11881
		x"ff",	--11882
		x"ff",	--11883
		x"ff",	--11884
		x"ff",	--11885
		x"ff",	--11886
		x"ff",	--11887
		x"ff",	--11888
		x"ff",	--11889
		x"ff",	--11890
		x"ff",	--11891
		x"ff",	--11892
		x"ff",	--11893
		x"ff",	--11894
		x"ff",	--11895
		x"ff",	--11896
		x"ff",	--11897
		x"ff",	--11898
		x"ff",	--11899
		x"ff",	--11900
		x"ff",	--11901
		x"ff",	--11902
		x"ff",	--11903
		x"ff",	--11904
		x"ff",	--11905
		x"ff",	--11906
		x"ff",	--11907
		x"ff",	--11908
		x"ff",	--11909
		x"ff",	--11910
		x"ff",	--11911
		x"ff",	--11912
		x"ff",	--11913
		x"ff",	--11914
		x"ff",	--11915
		x"ff",	--11916
		x"ff",	--11917
		x"ff",	--11918
		x"ff",	--11919
		x"ff",	--11920
		x"ff",	--11921
		x"ff",	--11922
		x"ff",	--11923
		x"ff",	--11924
		x"ff",	--11925
		x"ff",	--11926
		x"ff",	--11927
		x"ff",	--11928
		x"ff",	--11929
		x"ff",	--11930
		x"ff",	--11931
		x"ff",	--11932
		x"ff",	--11933
		x"ff",	--11934
		x"ff",	--11935
		x"ff",	--11936
		x"ff",	--11937
		x"ff",	--11938
		x"ff",	--11939
		x"ff",	--11940
		x"ff",	--11941
		x"ff",	--11942
		x"ff",	--11943
		x"ff",	--11944
		x"ff",	--11945
		x"ff",	--11946
		x"ff",	--11947
		x"ff",	--11948
		x"ff",	--11949
		x"ff",	--11950
		x"ff",	--11951
		x"ff",	--11952
		x"ff",	--11953
		x"ff",	--11954
		x"ff",	--11955
		x"ff",	--11956
		x"ff",	--11957
		x"ff",	--11958
		x"ff",	--11959
		x"ff",	--11960
		x"ff",	--11961
		x"ff",	--11962
		x"ff",	--11963
		x"ff",	--11964
		x"ff",	--11965
		x"ff",	--11966
		x"ff",	--11967
		x"ff",	--11968
		x"ff",	--11969
		x"ff",	--11970
		x"ff",	--11971
		x"ff",	--11972
		x"ff",	--11973
		x"ff",	--11974
		x"ff",	--11975
		x"ff",	--11976
		x"ff",	--11977
		x"ff",	--11978
		x"ff",	--11979
		x"ff",	--11980
		x"ff",	--11981
		x"ff",	--11982
		x"ff",	--11983
		x"ff",	--11984
		x"ff",	--11985
		x"ff",	--11986
		x"ff",	--11987
		x"ff",	--11988
		x"ff",	--11989
		x"ff",	--11990
		x"ff",	--11991
		x"ff",	--11992
		x"ff",	--11993
		x"ff",	--11994
		x"ff",	--11995
		x"ff",	--11996
		x"ff",	--11997
		x"ff",	--11998
		x"ff",	--11999
		x"ff",	--12000
		x"ff",	--12001
		x"ff",	--12002
		x"ff",	--12003
		x"ff",	--12004
		x"ff",	--12005
		x"ff",	--12006
		x"ff",	--12007
		x"ff",	--12008
		x"ff",	--12009
		x"ff",	--12010
		x"ff",	--12011
		x"ff",	--12012
		x"ff",	--12013
		x"ff",	--12014
		x"ff",	--12015
		x"ff",	--12016
		x"ff",	--12017
		x"ff",	--12018
		x"ff",	--12019
		x"ff",	--12020
		x"ff",	--12021
		x"ff",	--12022
		x"ff",	--12023
		x"ff",	--12024
		x"ff",	--12025
		x"ff",	--12026
		x"ff",	--12027
		x"ff",	--12028
		x"ff",	--12029
		x"ff",	--12030
		x"ff",	--12031
		x"ff",	--12032
		x"ff",	--12033
		x"ff",	--12034
		x"ff",	--12035
		x"ff",	--12036
		x"ff",	--12037
		x"ff",	--12038
		x"ff",	--12039
		x"ff",	--12040
		x"ff",	--12041
		x"ff",	--12042
		x"ff",	--12043
		x"ff",	--12044
		x"ff",	--12045
		x"ff",	--12046
		x"ff",	--12047
		x"ff",	--12048
		x"ff",	--12049
		x"ff",	--12050
		x"ff",	--12051
		x"ff",	--12052
		x"ff",	--12053
		x"ff",	--12054
		x"ff",	--12055
		x"ff",	--12056
		x"ff",	--12057
		x"ff",	--12058
		x"ff",	--12059
		x"ff",	--12060
		x"ff",	--12061
		x"ff",	--12062
		x"ff",	--12063
		x"ff",	--12064
		x"ff",	--12065
		x"ff",	--12066
		x"ff",	--12067
		x"ff",	--12068
		x"ff",	--12069
		x"ff",	--12070
		x"ff",	--12071
		x"ff",	--12072
		x"ff",	--12073
		x"ff",	--12074
		x"ff",	--12075
		x"ff",	--12076
		x"ff",	--12077
		x"ff",	--12078
		x"ff",	--12079
		x"ff",	--12080
		x"ff",	--12081
		x"ff",	--12082
		x"ff",	--12083
		x"ff",	--12084
		x"ff",	--12085
		x"ff",	--12086
		x"ff",	--12087
		x"ff",	--12088
		x"ff",	--12089
		x"ff",	--12090
		x"ff",	--12091
		x"ff",	--12092
		x"ff",	--12093
		x"ff",	--12094
		x"ff",	--12095
		x"ff",	--12096
		x"ff",	--12097
		x"ff",	--12098
		x"ff",	--12099
		x"ff",	--12100
		x"ff",	--12101
		x"ff",	--12102
		x"ff",	--12103
		x"ff",	--12104
		x"ff",	--12105
		x"ff",	--12106
		x"ff",	--12107
		x"ff",	--12108
		x"ff",	--12109
		x"ff",	--12110
		x"ff",	--12111
		x"ff",	--12112
		x"ff",	--12113
		x"ff",	--12114
		x"ff",	--12115
		x"ff",	--12116
		x"ff",	--12117
		x"ff",	--12118
		x"ff",	--12119
		x"ff",	--12120
		x"ff",	--12121
		x"ff",	--12122
		x"ff",	--12123
		x"ff",	--12124
		x"ff",	--12125
		x"ff",	--12126
		x"ff",	--12127
		x"ff",	--12128
		x"ff",	--12129
		x"ff",	--12130
		x"ff",	--12131
		x"ff",	--12132
		x"ff",	--12133
		x"ff",	--12134
		x"ff",	--12135
		x"ff",	--12136
		x"ff",	--12137
		x"ff",	--12138
		x"ff",	--12139
		x"ff",	--12140
		x"ff",	--12141
		x"ff",	--12142
		x"ff",	--12143
		x"ff",	--12144
		x"ff",	--12145
		x"ff",	--12146
		x"ff",	--12147
		x"ff",	--12148
		x"ff",	--12149
		x"ff",	--12150
		x"ff",	--12151
		x"ff",	--12152
		x"ff",	--12153
		x"ff",	--12154
		x"ff",	--12155
		x"ff",	--12156
		x"ff",	--12157
		x"ff",	--12158
		x"ff",	--12159
		x"ff",	--12160
		x"ff",	--12161
		x"ff",	--12162
		x"ff",	--12163
		x"ff",	--12164
		x"ff",	--12165
		x"ff",	--12166
		x"ff",	--12167
		x"ff",	--12168
		x"ff",	--12169
		x"ff",	--12170
		x"ff",	--12171
		x"ff",	--12172
		x"ff",	--12173
		x"ff",	--12174
		x"ff",	--12175
		x"ff",	--12176
		x"ff",	--12177
		x"ff",	--12178
		x"ff",	--12179
		x"ff",	--12180
		x"ff",	--12181
		x"ff",	--12182
		x"ff",	--12183
		x"ff",	--12184
		x"ff",	--12185
		x"ff",	--12186
		x"ff",	--12187
		x"ff",	--12188
		x"ff",	--12189
		x"ff",	--12190
		x"ff",	--12191
		x"ff",	--12192
		x"ff",	--12193
		x"ff",	--12194
		x"ff",	--12195
		x"ff",	--12196
		x"ff",	--12197
		x"ff",	--12198
		x"ff",	--12199
		x"ff",	--12200
		x"ff",	--12201
		x"ff",	--12202
		x"ff",	--12203
		x"ff",	--12204
		x"ff",	--12205
		x"ff",	--12206
		x"ff",	--12207
		x"ff",	--12208
		x"ff",	--12209
		x"ff",	--12210
		x"ff",	--12211
		x"ff",	--12212
		x"ff",	--12213
		x"ff",	--12214
		x"ff",	--12215
		x"ff",	--12216
		x"ff",	--12217
		x"ff",	--12218
		x"ff",	--12219
		x"ff",	--12220
		x"ff",	--12221
		x"ff",	--12222
		x"ff",	--12223
		x"ff",	--12224
		x"ff",	--12225
		x"ff",	--12226
		x"ff",	--12227
		x"ff",	--12228
		x"ff",	--12229
		x"ff",	--12230
		x"ff",	--12231
		x"ff",	--12232
		x"ff",	--12233
		x"ff",	--12234
		x"ff",	--12235
		x"ff",	--12236
		x"ff",	--12237
		x"ff",	--12238
		x"ff",	--12239
		x"ff",	--12240
		x"ff",	--12241
		x"ff",	--12242
		x"ff",	--12243
		x"ff",	--12244
		x"ff",	--12245
		x"ff",	--12246
		x"ff",	--12247
		x"ff",	--12248
		x"ff",	--12249
		x"ff",	--12250
		x"ff",	--12251
		x"ff",	--12252
		x"ff",	--12253
		x"ff",	--12254
		x"ff",	--12255
		x"ff",	--12256
		x"ff",	--12257
		x"ff",	--12258
		x"ff",	--12259
		x"ff",	--12260
		x"ff",	--12261
		x"ff",	--12262
		x"ff",	--12263
		x"ff",	--12264
		x"ff",	--12265
		x"ff",	--12266
		x"ff",	--12267
		x"ff",	--12268
		x"ff",	--12269
		x"ff",	--12270
		x"ff",	--12271
		x"ff",	--12272
		x"ff",	--12273
		x"ff",	--12274
		x"ff",	--12275
		x"ff",	--12276
		x"ff",	--12277
		x"ff",	--12278
		x"ff",	--12279
		x"ff",	--12280
		x"ff",	--12281
		x"ff",	--12282
		x"ff",	--12283
		x"ff",	--12284
		x"ff",	--12285
		x"ff",	--12286
		x"ff",	--12287
		x"ff",	--12288
		x"ff",	--12289
		x"ff",	--12290
		x"ff",	--12291
		x"ff",	--12292
		x"ff",	--12293
		x"ff",	--12294
		x"ff",	--12295
		x"ff",	--12296
		x"ff",	--12297
		x"ff",	--12298
		x"ff",	--12299
		x"ff",	--12300
		x"ff",	--12301
		x"ff",	--12302
		x"ff",	--12303
		x"ff",	--12304
		x"ff",	--12305
		x"ff",	--12306
		x"ff",	--12307
		x"ff",	--12308
		x"ff",	--12309
		x"ff",	--12310
		x"ff",	--12311
		x"ff",	--12312
		x"ff",	--12313
		x"ff",	--12314
		x"ff",	--12315
		x"ff",	--12316
		x"ff",	--12317
		x"ff",	--12318
		x"ff",	--12319
		x"ff",	--12320
		x"ff",	--12321
		x"ff",	--12322
		x"ff",	--12323
		x"ff",	--12324
		x"ff",	--12325
		x"ff",	--12326
		x"ff",	--12327
		x"ff",	--12328
		x"ff",	--12329
		x"ff",	--12330
		x"ff",	--12331
		x"ff",	--12332
		x"ff",	--12333
		x"ff",	--12334
		x"ff",	--12335
		x"ff",	--12336
		x"ff",	--12337
		x"ff",	--12338
		x"ff",	--12339
		x"ff",	--12340
		x"ff",	--12341
		x"ff",	--12342
		x"ff",	--12343
		x"ff",	--12344
		x"ff",	--12345
		x"ff",	--12346
		x"ff",	--12347
		x"ff",	--12348
		x"ff",	--12349
		x"ff",	--12350
		x"ff",	--12351
		x"ff",	--12352
		x"ff",	--12353
		x"ff",	--12354
		x"ff",	--12355
		x"ff",	--12356
		x"ff",	--12357
		x"ff",	--12358
		x"ff",	--12359
		x"ff",	--12360
		x"ff",	--12361
		x"ff",	--12362
		x"ff",	--12363
		x"ff",	--12364
		x"ff",	--12365
		x"ff",	--12366
		x"ff",	--12367
		x"ff",	--12368
		x"ff",	--12369
		x"ff",	--12370
		x"ff",	--12371
		x"ff",	--12372
		x"ff",	--12373
		x"ff",	--12374
		x"ff",	--12375
		x"ff",	--12376
		x"ff",	--12377
		x"ff",	--12378
		x"ff",	--12379
		x"ff",	--12380
		x"ff",	--12381
		x"ff",	--12382
		x"ff",	--12383
		x"ff",	--12384
		x"ff",	--12385
		x"ff",	--12386
		x"ff",	--12387
		x"ff",	--12388
		x"ff",	--12389
		x"ff",	--12390
		x"ff",	--12391
		x"ff",	--12392
		x"ff",	--12393
		x"ff",	--12394
		x"ff",	--12395
		x"ff",	--12396
		x"ff",	--12397
		x"ff",	--12398
		x"ff",	--12399
		x"ff",	--12400
		x"ff",	--12401
		x"ff",	--12402
		x"ff",	--12403
		x"ff",	--12404
		x"ff",	--12405
		x"ff",	--12406
		x"ff",	--12407
		x"ff",	--12408
		x"ff",	--12409
		x"ff",	--12410
		x"ff",	--12411
		x"ff",	--12412
		x"ff",	--12413
		x"ff",	--12414
		x"ff",	--12415
		x"ff",	--12416
		x"ff",	--12417
		x"ff",	--12418
		x"ff",	--12419
		x"ff",	--12420
		x"ff",	--12421
		x"ff",	--12422
		x"ff",	--12423
		x"ff",	--12424
		x"ff",	--12425
		x"ff",	--12426
		x"ff",	--12427
		x"ff",	--12428
		x"ff",	--12429
		x"ff",	--12430
		x"ff",	--12431
		x"ff",	--12432
		x"ff",	--12433
		x"ff",	--12434
		x"ff",	--12435
		x"ff",	--12436
		x"ff",	--12437
		x"ff",	--12438
		x"ff",	--12439
		x"ff",	--12440
		x"ff",	--12441
		x"ff",	--12442
		x"ff",	--12443
		x"ff",	--12444
		x"ff",	--12445
		x"ff",	--12446
		x"ff",	--12447
		x"ff",	--12448
		x"ff",	--12449
		x"ff",	--12450
		x"ff",	--12451
		x"ff",	--12452
		x"ff",	--12453
		x"ff",	--12454
		x"ff",	--12455
		x"ff",	--12456
		x"ff",	--12457
		x"ff",	--12458
		x"ff",	--12459
		x"ff",	--12460
		x"ff",	--12461
		x"ff",	--12462
		x"ff",	--12463
		x"ff",	--12464
		x"ff",	--12465
		x"ff",	--12466
		x"ff",	--12467
		x"ff",	--12468
		x"ff",	--12469
		x"ff",	--12470
		x"ff",	--12471
		x"ff",	--12472
		x"ff",	--12473
		x"ff",	--12474
		x"ff",	--12475
		x"ff",	--12476
		x"ff",	--12477
		x"ff",	--12478
		x"ff",	--12479
		x"ff",	--12480
		x"ff",	--12481
		x"ff",	--12482
		x"ff",	--12483
		x"ff",	--12484
		x"ff",	--12485
		x"ff",	--12486
		x"ff",	--12487
		x"ff",	--12488
		x"ff",	--12489
		x"ff",	--12490
		x"ff",	--12491
		x"ff",	--12492
		x"ff",	--12493
		x"ff",	--12494
		x"ff",	--12495
		x"ff",	--12496
		x"ff",	--12497
		x"ff",	--12498
		x"ff",	--12499
		x"ff",	--12500
		x"ff",	--12501
		x"ff",	--12502
		x"ff",	--12503
		x"ff",	--12504
		x"ff",	--12505
		x"ff",	--12506
		x"ff",	--12507
		x"ff",	--12508
		x"ff",	--12509
		x"ff",	--12510
		x"ff",	--12511
		x"ff",	--12512
		x"ff",	--12513
		x"ff",	--12514
		x"ff",	--12515
		x"ff",	--12516
		x"ff",	--12517
		x"ff",	--12518
		x"ff",	--12519
		x"ff",	--12520
		x"ff",	--12521
		x"ff",	--12522
		x"ff",	--12523
		x"ff",	--12524
		x"ff",	--12525
		x"ff",	--12526
		x"ff",	--12527
		x"ff",	--12528
		x"ff",	--12529
		x"ff",	--12530
		x"ff",	--12531
		x"ff",	--12532
		x"ff",	--12533
		x"ff",	--12534
		x"ff",	--12535
		x"ff",	--12536
		x"ff",	--12537
		x"ff",	--12538
		x"ff",	--12539
		x"ff",	--12540
		x"ff",	--12541
		x"ff",	--12542
		x"ff",	--12543
		x"ff",	--12544
		x"ff",	--12545
		x"ff",	--12546
		x"ff",	--12547
		x"ff",	--12548
		x"ff",	--12549
		x"ff",	--12550
		x"ff",	--12551
		x"ff",	--12552
		x"ff",	--12553
		x"ff",	--12554
		x"ff",	--12555
		x"ff",	--12556
		x"ff",	--12557
		x"ff",	--12558
		x"ff",	--12559
		x"ff",	--12560
		x"ff",	--12561
		x"ff",	--12562
		x"ff",	--12563
		x"ff",	--12564
		x"ff",	--12565
		x"ff",	--12566
		x"ff",	--12567
		x"ff",	--12568
		x"ff",	--12569
		x"ff",	--12570
		x"ff",	--12571
		x"ff",	--12572
		x"ff",	--12573
		x"ff",	--12574
		x"ff",	--12575
		x"ff",	--12576
		x"ff",	--12577
		x"ff",	--12578
		x"ff",	--12579
		x"ff",	--12580
		x"ff",	--12581
		x"ff",	--12582
		x"ff",	--12583
		x"ff",	--12584
		x"ff",	--12585
		x"ff",	--12586
		x"ff",	--12587
		x"ff",	--12588
		x"ff",	--12589
		x"ff",	--12590
		x"ff",	--12591
		x"ff",	--12592
		x"ff",	--12593
		x"ff",	--12594
		x"ff",	--12595
		x"ff",	--12596
		x"ff",	--12597
		x"ff",	--12598
		x"ff",	--12599
		x"ff",	--12600
		x"ff",	--12601
		x"ff",	--12602
		x"ff",	--12603
		x"ff",	--12604
		x"ff",	--12605
		x"ff",	--12606
		x"ff",	--12607
		x"ff",	--12608
		x"ff",	--12609
		x"ff",	--12610
		x"ff",	--12611
		x"ff",	--12612
		x"ff",	--12613
		x"ff",	--12614
		x"ff",	--12615
		x"ff",	--12616
		x"ff",	--12617
		x"ff",	--12618
		x"ff",	--12619
		x"ff",	--12620
		x"ff",	--12621
		x"ff",	--12622
		x"ff",	--12623
		x"ff",	--12624
		x"ff",	--12625
		x"ff",	--12626
		x"ff",	--12627
		x"ff",	--12628
		x"ff",	--12629
		x"ff",	--12630
		x"ff",	--12631
		x"ff",	--12632
		x"ff",	--12633
		x"ff",	--12634
		x"ff",	--12635
		x"ff",	--12636
		x"ff",	--12637
		x"ff",	--12638
		x"ff",	--12639
		x"ff",	--12640
		x"ff",	--12641
		x"ff",	--12642
		x"ff",	--12643
		x"ff",	--12644
		x"ff",	--12645
		x"ff",	--12646
		x"ff",	--12647
		x"ff",	--12648
		x"ff",	--12649
		x"ff",	--12650
		x"ff",	--12651
		x"ff",	--12652
		x"ff",	--12653
		x"ff",	--12654
		x"ff",	--12655
		x"ff",	--12656
		x"ff",	--12657
		x"ff",	--12658
		x"ff",	--12659
		x"ff",	--12660
		x"ff",	--12661
		x"ff",	--12662
		x"ff",	--12663
		x"ff",	--12664
		x"ff",	--12665
		x"ff",	--12666
		x"ff",	--12667
		x"ff",	--12668
		x"ff",	--12669
		x"ff",	--12670
		x"ff",	--12671
		x"ff",	--12672
		x"ff",	--12673
		x"ff",	--12674
		x"ff",	--12675
		x"ff",	--12676
		x"ff",	--12677
		x"ff",	--12678
		x"ff",	--12679
		x"ff",	--12680
		x"ff",	--12681
		x"ff",	--12682
		x"ff",	--12683
		x"ff",	--12684
		x"ff",	--12685
		x"ff",	--12686
		x"ff",	--12687
		x"ff",	--12688
		x"ff",	--12689
		x"ff",	--12690
		x"ff",	--12691
		x"ff",	--12692
		x"ff",	--12693
		x"ff",	--12694
		x"ff",	--12695
		x"ff",	--12696
		x"ff",	--12697
		x"ff",	--12698
		x"ff",	--12699
		x"ff",	--12700
		x"ff",	--12701
		x"ff",	--12702
		x"ff",	--12703
		x"ff",	--12704
		x"ff",	--12705
		x"ff",	--12706
		x"ff",	--12707
		x"ff",	--12708
		x"ff",	--12709
		x"ff",	--12710
		x"ff",	--12711
		x"ff",	--12712
		x"ff",	--12713
		x"ff",	--12714
		x"ff",	--12715
		x"ff",	--12716
		x"ff",	--12717
		x"ff",	--12718
		x"ff",	--12719
		x"ff",	--12720
		x"ff",	--12721
		x"ff",	--12722
		x"ff",	--12723
		x"ff",	--12724
		x"ff",	--12725
		x"ff",	--12726
		x"ff",	--12727
		x"ff",	--12728
		x"ff",	--12729
		x"ff",	--12730
		x"ff",	--12731
		x"ff",	--12732
		x"ff",	--12733
		x"ff",	--12734
		x"ff",	--12735
		x"ff",	--12736
		x"ff",	--12737
		x"ff",	--12738
		x"ff",	--12739
		x"ff",	--12740
		x"ff",	--12741
		x"ff",	--12742
		x"ff",	--12743
		x"ff",	--12744
		x"ff",	--12745
		x"ff",	--12746
		x"ff",	--12747
		x"ff",	--12748
		x"ff",	--12749
		x"ff",	--12750
		x"ff",	--12751
		x"ff",	--12752
		x"ff",	--12753
		x"ff",	--12754
		x"ff",	--12755
		x"ff",	--12756
		x"ff",	--12757
		x"ff",	--12758
		x"ff",	--12759
		x"ff",	--12760
		x"ff",	--12761
		x"ff",	--12762
		x"ff",	--12763
		x"ff",	--12764
		x"ff",	--12765
		x"ff",	--12766
		x"ff",	--12767
		x"ff",	--12768
		x"ff",	--12769
		x"ff",	--12770
		x"ff",	--12771
		x"ff",	--12772
		x"ff",	--12773
		x"ff",	--12774
		x"ff",	--12775
		x"ff",	--12776
		x"ff",	--12777
		x"ff",	--12778
		x"ff",	--12779
		x"ff",	--12780
		x"ff",	--12781
		x"ff",	--12782
		x"ff",	--12783
		x"ff",	--12784
		x"ff",	--12785
		x"ff",	--12786
		x"ff",	--12787
		x"ff",	--12788
		x"ff",	--12789
		x"ff",	--12790
		x"ff",	--12791
		x"ff",	--12792
		x"ff",	--12793
		x"ff",	--12794
		x"ff",	--12795
		x"ff",	--12796
		x"ff",	--12797
		x"ff",	--12798
		x"ff",	--12799
		x"ff",	--12800
		x"ff",	--12801
		x"ff",	--12802
		x"ff",	--12803
		x"ff",	--12804
		x"ff",	--12805
		x"ff",	--12806
		x"ff",	--12807
		x"ff",	--12808
		x"ff",	--12809
		x"ff",	--12810
		x"ff",	--12811
		x"ff",	--12812
		x"ff",	--12813
		x"ff",	--12814
		x"ff",	--12815
		x"ff",	--12816
		x"ff",	--12817
		x"ff",	--12818
		x"ff",	--12819
		x"ff",	--12820
		x"ff",	--12821
		x"ff",	--12822
		x"ff",	--12823
		x"ff",	--12824
		x"ff",	--12825
		x"ff",	--12826
		x"ff",	--12827
		x"ff",	--12828
		x"ff",	--12829
		x"ff",	--12830
		x"ff",	--12831
		x"ff",	--12832
		x"ff",	--12833
		x"ff",	--12834
		x"ff",	--12835
		x"ff",	--12836
		x"ff",	--12837
		x"ff",	--12838
		x"ff",	--12839
		x"ff",	--12840
		x"ff",	--12841
		x"ff",	--12842
		x"ff",	--12843
		x"ff",	--12844
		x"ff",	--12845
		x"ff",	--12846
		x"ff",	--12847
		x"ff",	--12848
		x"ff",	--12849
		x"ff",	--12850
		x"ff",	--12851
		x"ff",	--12852
		x"ff",	--12853
		x"ff",	--12854
		x"ff",	--12855
		x"ff",	--12856
		x"ff",	--12857
		x"ff",	--12858
		x"ff",	--12859
		x"ff",	--12860
		x"ff",	--12861
		x"ff",	--12862
		x"ff",	--12863
		x"ff",	--12864
		x"ff",	--12865
		x"ff",	--12866
		x"ff",	--12867
		x"ff",	--12868
		x"ff",	--12869
		x"ff",	--12870
		x"ff",	--12871
		x"ff",	--12872
		x"ff",	--12873
		x"ff",	--12874
		x"ff",	--12875
		x"ff",	--12876
		x"ff",	--12877
		x"ff",	--12878
		x"ff",	--12879
		x"ff",	--12880
		x"ff",	--12881
		x"ff",	--12882
		x"ff",	--12883
		x"ff",	--12884
		x"ff",	--12885
		x"ff",	--12886
		x"ff",	--12887
		x"ff",	--12888
		x"ff",	--12889
		x"ff",	--12890
		x"ff",	--12891
		x"ff",	--12892
		x"ff",	--12893
		x"ff",	--12894
		x"ff",	--12895
		x"ff",	--12896
		x"ff",	--12897
		x"ff",	--12898
		x"ff",	--12899
		x"ff",	--12900
		x"ff",	--12901
		x"ff",	--12902
		x"ff",	--12903
		x"ff",	--12904
		x"ff",	--12905
		x"ff",	--12906
		x"ff",	--12907
		x"ff",	--12908
		x"ff",	--12909
		x"ff",	--12910
		x"ff",	--12911
		x"ff",	--12912
		x"ff",	--12913
		x"ff",	--12914
		x"ff",	--12915
		x"ff",	--12916
		x"ff",	--12917
		x"ff",	--12918
		x"ff",	--12919
		x"ff",	--12920
		x"ff",	--12921
		x"ff",	--12922
		x"ff",	--12923
		x"ff",	--12924
		x"ff",	--12925
		x"ff",	--12926
		x"ff",	--12927
		x"ff",	--12928
		x"ff",	--12929
		x"ff",	--12930
		x"ff",	--12931
		x"ff",	--12932
		x"ff",	--12933
		x"ff",	--12934
		x"ff",	--12935
		x"ff",	--12936
		x"ff",	--12937
		x"ff",	--12938
		x"ff",	--12939
		x"ff",	--12940
		x"ff",	--12941
		x"ff",	--12942
		x"ff",	--12943
		x"ff",	--12944
		x"ff",	--12945
		x"ff",	--12946
		x"ff",	--12947
		x"ff",	--12948
		x"ff",	--12949
		x"ff",	--12950
		x"ff",	--12951
		x"ff",	--12952
		x"ff",	--12953
		x"ff",	--12954
		x"ff",	--12955
		x"ff",	--12956
		x"ff",	--12957
		x"ff",	--12958
		x"ff",	--12959
		x"ff",	--12960
		x"ff",	--12961
		x"ff",	--12962
		x"ff",	--12963
		x"ff",	--12964
		x"ff",	--12965
		x"ff",	--12966
		x"ff",	--12967
		x"ff",	--12968
		x"ff",	--12969
		x"ff",	--12970
		x"ff",	--12971
		x"ff",	--12972
		x"ff",	--12973
		x"ff",	--12974
		x"ff",	--12975
		x"ff",	--12976
		x"ff",	--12977
		x"ff",	--12978
		x"ff",	--12979
		x"ff",	--12980
		x"ff",	--12981
		x"ff",	--12982
		x"ff",	--12983
		x"ff",	--12984
		x"ff",	--12985
		x"ff",	--12986
		x"ff",	--12987
		x"ff",	--12988
		x"ff",	--12989
		x"ff",	--12990
		x"ff",	--12991
		x"ff",	--12992
		x"ff",	--12993
		x"ff",	--12994
		x"ff",	--12995
		x"ff",	--12996
		x"ff",	--12997
		x"ff",	--12998
		x"ff",	--12999
		x"ff",	--13000
		x"ff",	--13001
		x"ff",	--13002
		x"ff",	--13003
		x"ff",	--13004
		x"ff",	--13005
		x"ff",	--13006
		x"ff",	--13007
		x"ff",	--13008
		x"ff",	--13009
		x"ff",	--13010
		x"ff",	--13011
		x"ff",	--13012
		x"ff",	--13013
		x"ff",	--13014
		x"ff",	--13015
		x"ff",	--13016
		x"ff",	--13017
		x"ff",	--13018
		x"ff",	--13019
		x"ff",	--13020
		x"ff",	--13021
		x"ff",	--13022
		x"ff",	--13023
		x"ff",	--13024
		x"ff",	--13025
		x"ff",	--13026
		x"ff",	--13027
		x"ff",	--13028
		x"ff",	--13029
		x"ff",	--13030
		x"ff",	--13031
		x"ff",	--13032
		x"ff",	--13033
		x"ff",	--13034
		x"ff",	--13035
		x"ff",	--13036
		x"ff",	--13037
		x"ff",	--13038
		x"ff",	--13039
		x"ff",	--13040
		x"ff",	--13041
		x"ff",	--13042
		x"ff",	--13043
		x"ff",	--13044
		x"ff",	--13045
		x"ff",	--13046
		x"ff",	--13047
		x"ff",	--13048
		x"ff",	--13049
		x"ff",	--13050
		x"ff",	--13051
		x"ff",	--13052
		x"ff",	--13053
		x"ff",	--13054
		x"ff",	--13055
		x"ff",	--13056
		x"ff",	--13057
		x"ff",	--13058
		x"ff",	--13059
		x"ff",	--13060
		x"ff",	--13061
		x"ff",	--13062
		x"ff",	--13063
		x"ff",	--13064
		x"ff",	--13065
		x"ff",	--13066
		x"ff",	--13067
		x"ff",	--13068
		x"ff",	--13069
		x"ff",	--13070
		x"ff",	--13071
		x"ff",	--13072
		x"ff",	--13073
		x"ff",	--13074
		x"ff",	--13075
		x"ff",	--13076
		x"ff",	--13077
		x"ff",	--13078
		x"ff",	--13079
		x"ff",	--13080
		x"ff",	--13081
		x"ff",	--13082
		x"ff",	--13083
		x"ff",	--13084
		x"ff",	--13085
		x"ff",	--13086
		x"ff",	--13087
		x"ff",	--13088
		x"ff",	--13089
		x"ff",	--13090
		x"ff",	--13091
		x"ff",	--13092
		x"ff",	--13093
		x"ff",	--13094
		x"ff",	--13095
		x"ff",	--13096
		x"ff",	--13097
		x"ff",	--13098
		x"ff",	--13099
		x"ff",	--13100
		x"ff",	--13101
		x"ff",	--13102
		x"ff",	--13103
		x"ff",	--13104
		x"ff",	--13105
		x"ff",	--13106
		x"ff",	--13107
		x"ff",	--13108
		x"ff",	--13109
		x"ff",	--13110
		x"ff",	--13111
		x"ff",	--13112
		x"ff",	--13113
		x"ff",	--13114
		x"ff",	--13115
		x"ff",	--13116
		x"ff",	--13117
		x"ff",	--13118
		x"ff",	--13119
		x"ff",	--13120
		x"ff",	--13121
		x"ff",	--13122
		x"ff",	--13123
		x"ff",	--13124
		x"ff",	--13125
		x"ff",	--13126
		x"ff",	--13127
		x"ff",	--13128
		x"ff",	--13129
		x"ff",	--13130
		x"ff",	--13131
		x"ff",	--13132
		x"ff",	--13133
		x"ff",	--13134
		x"ff",	--13135
		x"ff",	--13136
		x"ff",	--13137
		x"ff",	--13138
		x"ff",	--13139
		x"ff",	--13140
		x"ff",	--13141
		x"ff",	--13142
		x"ff",	--13143
		x"ff",	--13144
		x"ff",	--13145
		x"ff",	--13146
		x"ff",	--13147
		x"ff",	--13148
		x"ff",	--13149
		x"ff",	--13150
		x"ff",	--13151
		x"ff",	--13152
		x"ff",	--13153
		x"ff",	--13154
		x"ff",	--13155
		x"ff",	--13156
		x"ff",	--13157
		x"ff",	--13158
		x"ff",	--13159
		x"ff",	--13160
		x"ff",	--13161
		x"ff",	--13162
		x"ff",	--13163
		x"ff",	--13164
		x"ff",	--13165
		x"ff",	--13166
		x"ff",	--13167
		x"ff",	--13168
		x"ff",	--13169
		x"ff",	--13170
		x"ff",	--13171
		x"ff",	--13172
		x"ff",	--13173
		x"ff",	--13174
		x"ff",	--13175
		x"ff",	--13176
		x"ff",	--13177
		x"ff",	--13178
		x"ff",	--13179
		x"ff",	--13180
		x"ff",	--13181
		x"ff",	--13182
		x"ff",	--13183
		x"ff",	--13184
		x"ff",	--13185
		x"ff",	--13186
		x"ff",	--13187
		x"ff",	--13188
		x"ff",	--13189
		x"ff",	--13190
		x"ff",	--13191
		x"ff",	--13192
		x"ff",	--13193
		x"ff",	--13194
		x"ff",	--13195
		x"ff",	--13196
		x"ff",	--13197
		x"ff",	--13198
		x"ff",	--13199
		x"ff",	--13200
		x"ff",	--13201
		x"ff",	--13202
		x"ff",	--13203
		x"ff",	--13204
		x"ff",	--13205
		x"ff",	--13206
		x"ff",	--13207
		x"ff",	--13208
		x"ff",	--13209
		x"ff",	--13210
		x"ff",	--13211
		x"ff",	--13212
		x"ff",	--13213
		x"ff",	--13214
		x"ff",	--13215
		x"ff",	--13216
		x"ff",	--13217
		x"ff",	--13218
		x"ff",	--13219
		x"ff",	--13220
		x"ff",	--13221
		x"ff",	--13222
		x"ff",	--13223
		x"ff",	--13224
		x"ff",	--13225
		x"ff",	--13226
		x"ff",	--13227
		x"ff",	--13228
		x"ff",	--13229
		x"ff",	--13230
		x"ff",	--13231
		x"ff",	--13232
		x"ff",	--13233
		x"ff",	--13234
		x"ff",	--13235
		x"ff",	--13236
		x"ff",	--13237
		x"ff",	--13238
		x"ff",	--13239
		x"ff",	--13240
		x"ff",	--13241
		x"ff",	--13242
		x"ff",	--13243
		x"ff",	--13244
		x"ff",	--13245
		x"ff",	--13246
		x"ff",	--13247
		x"ff",	--13248
		x"ff",	--13249
		x"ff",	--13250
		x"ff",	--13251
		x"ff",	--13252
		x"ff",	--13253
		x"ff",	--13254
		x"ff",	--13255
		x"ff",	--13256
		x"ff",	--13257
		x"ff",	--13258
		x"ff",	--13259
		x"ff",	--13260
		x"ff",	--13261
		x"ff",	--13262
		x"ff",	--13263
		x"ff",	--13264
		x"ff",	--13265
		x"ff",	--13266
		x"ff",	--13267
		x"ff",	--13268
		x"ff",	--13269
		x"ff",	--13270
		x"ff",	--13271
		x"ff",	--13272
		x"ff",	--13273
		x"ff",	--13274
		x"ff",	--13275
		x"ff",	--13276
		x"ff",	--13277
		x"ff",	--13278
		x"ff",	--13279
		x"ff",	--13280
		x"ff",	--13281
		x"ff",	--13282
		x"ff",	--13283
		x"ff",	--13284
		x"ff",	--13285
		x"ff",	--13286
		x"ff",	--13287
		x"ff",	--13288
		x"ff",	--13289
		x"ff",	--13290
		x"ff",	--13291
		x"ff",	--13292
		x"ff",	--13293
		x"ff",	--13294
		x"ff",	--13295
		x"ff",	--13296
		x"ff",	--13297
		x"ff",	--13298
		x"ff",	--13299
		x"ff",	--13300
		x"ff",	--13301
		x"ff",	--13302
		x"ff",	--13303
		x"ff",	--13304
		x"ff",	--13305
		x"ff",	--13306
		x"ff",	--13307
		x"ff",	--13308
		x"ff",	--13309
		x"ff",	--13310
		x"ff",	--13311
		x"ff",	--13312
		x"ff",	--13313
		x"ff",	--13314
		x"ff",	--13315
		x"ff",	--13316
		x"ff",	--13317
		x"ff",	--13318
		x"ff",	--13319
		x"ff",	--13320
		x"ff",	--13321
		x"ff",	--13322
		x"ff",	--13323
		x"ff",	--13324
		x"ff",	--13325
		x"ff",	--13326
		x"ff",	--13327
		x"ff",	--13328
		x"ff",	--13329
		x"ff",	--13330
		x"ff",	--13331
		x"ff",	--13332
		x"ff",	--13333
		x"ff",	--13334
		x"ff",	--13335
		x"ff",	--13336
		x"ff",	--13337
		x"ff",	--13338
		x"ff",	--13339
		x"ff",	--13340
		x"ff",	--13341
		x"ff",	--13342
		x"ff",	--13343
		x"ff",	--13344
		x"ff",	--13345
		x"ff",	--13346
		x"ff",	--13347
		x"ff",	--13348
		x"ff",	--13349
		x"ff",	--13350
		x"ff",	--13351
		x"ff",	--13352
		x"ff",	--13353
		x"ff",	--13354
		x"ff",	--13355
		x"ff",	--13356
		x"ff",	--13357
		x"ff",	--13358
		x"ff",	--13359
		x"ff",	--13360
		x"ff",	--13361
		x"ff",	--13362
		x"ff",	--13363
		x"ff",	--13364
		x"ff",	--13365
		x"ff",	--13366
		x"ff",	--13367
		x"ff",	--13368
		x"ff",	--13369
		x"ff",	--13370
		x"ff",	--13371
		x"ff",	--13372
		x"ff",	--13373
		x"ff",	--13374
		x"ff",	--13375
		x"ff",	--13376
		x"ff",	--13377
		x"ff",	--13378
		x"ff",	--13379
		x"ff",	--13380
		x"ff",	--13381
		x"ff",	--13382
		x"ff",	--13383
		x"ff",	--13384
		x"ff",	--13385
		x"ff",	--13386
		x"ff",	--13387
		x"ff",	--13388
		x"ff",	--13389
		x"ff",	--13390
		x"ff",	--13391
		x"ff",	--13392
		x"ff",	--13393
		x"ff",	--13394
		x"ff",	--13395
		x"ff",	--13396
		x"ff",	--13397
		x"ff",	--13398
		x"ff",	--13399
		x"ff",	--13400
		x"ff",	--13401
		x"ff",	--13402
		x"ff",	--13403
		x"ff",	--13404
		x"ff",	--13405
		x"ff",	--13406
		x"ff",	--13407
		x"ff",	--13408
		x"ff",	--13409
		x"ff",	--13410
		x"ff",	--13411
		x"ff",	--13412
		x"ff",	--13413
		x"ff",	--13414
		x"ff",	--13415
		x"ff",	--13416
		x"ff",	--13417
		x"ff",	--13418
		x"ff",	--13419
		x"ff",	--13420
		x"ff",	--13421
		x"ff",	--13422
		x"ff",	--13423
		x"ff",	--13424
		x"ff",	--13425
		x"ff",	--13426
		x"ff",	--13427
		x"ff",	--13428
		x"ff",	--13429
		x"ff",	--13430
		x"ff",	--13431
		x"ff",	--13432
		x"ff",	--13433
		x"ff",	--13434
		x"ff",	--13435
		x"ff",	--13436
		x"ff",	--13437
		x"ff",	--13438
		x"ff",	--13439
		x"ff",	--13440
		x"ff",	--13441
		x"ff",	--13442
		x"ff",	--13443
		x"ff",	--13444
		x"ff",	--13445
		x"ff",	--13446
		x"ff",	--13447
		x"ff",	--13448
		x"ff",	--13449
		x"ff",	--13450
		x"ff",	--13451
		x"ff",	--13452
		x"ff",	--13453
		x"ff",	--13454
		x"ff",	--13455
		x"ff",	--13456
		x"ff",	--13457
		x"ff",	--13458
		x"ff",	--13459
		x"ff",	--13460
		x"ff",	--13461
		x"ff",	--13462
		x"ff",	--13463
		x"ff",	--13464
		x"ff",	--13465
		x"ff",	--13466
		x"ff",	--13467
		x"ff",	--13468
		x"ff",	--13469
		x"ff",	--13470
		x"ff",	--13471
		x"ff",	--13472
		x"ff",	--13473
		x"ff",	--13474
		x"ff",	--13475
		x"ff",	--13476
		x"ff",	--13477
		x"ff",	--13478
		x"ff",	--13479
		x"ff",	--13480
		x"ff",	--13481
		x"ff",	--13482
		x"ff",	--13483
		x"ff",	--13484
		x"ff",	--13485
		x"ff",	--13486
		x"ff",	--13487
		x"ff",	--13488
		x"ff",	--13489
		x"ff",	--13490
		x"ff",	--13491
		x"ff",	--13492
		x"ff",	--13493
		x"ff",	--13494
		x"ff",	--13495
		x"ff",	--13496
		x"ff",	--13497
		x"ff",	--13498
		x"ff",	--13499
		x"ff",	--13500
		x"ff",	--13501
		x"ff",	--13502
		x"ff",	--13503
		x"ff",	--13504
		x"ff",	--13505
		x"ff",	--13506
		x"ff",	--13507
		x"ff",	--13508
		x"ff",	--13509
		x"ff",	--13510
		x"ff",	--13511
		x"ff",	--13512
		x"ff",	--13513
		x"ff",	--13514
		x"ff",	--13515
		x"ff",	--13516
		x"ff",	--13517
		x"ff",	--13518
		x"ff",	--13519
		x"ff",	--13520
		x"ff",	--13521
		x"ff",	--13522
		x"ff",	--13523
		x"ff",	--13524
		x"ff",	--13525
		x"ff",	--13526
		x"ff",	--13527
		x"ff",	--13528
		x"ff",	--13529
		x"ff",	--13530
		x"ff",	--13531
		x"ff",	--13532
		x"ff",	--13533
		x"ff",	--13534
		x"ff",	--13535
		x"ff",	--13536
		x"ff",	--13537
		x"ff",	--13538
		x"ff",	--13539
		x"ff",	--13540
		x"ff",	--13541
		x"ff",	--13542
		x"ff",	--13543
		x"ff",	--13544
		x"ff",	--13545
		x"ff",	--13546
		x"ff",	--13547
		x"ff",	--13548
		x"ff",	--13549
		x"ff",	--13550
		x"ff",	--13551
		x"ff",	--13552
		x"ff",	--13553
		x"ff",	--13554
		x"ff",	--13555
		x"ff",	--13556
		x"ff",	--13557
		x"ff",	--13558
		x"ff",	--13559
		x"ff",	--13560
		x"ff",	--13561
		x"ff",	--13562
		x"ff",	--13563
		x"ff",	--13564
		x"ff",	--13565
		x"ff",	--13566
		x"ff",	--13567
		x"ff",	--13568
		x"ff",	--13569
		x"ff",	--13570
		x"ff",	--13571
		x"ff",	--13572
		x"ff",	--13573
		x"ff",	--13574
		x"ff",	--13575
		x"ff",	--13576
		x"ff",	--13577
		x"ff",	--13578
		x"ff",	--13579
		x"ff",	--13580
		x"ff",	--13581
		x"ff",	--13582
		x"ff",	--13583
		x"ff",	--13584
		x"ff",	--13585
		x"ff",	--13586
		x"ff",	--13587
		x"ff",	--13588
		x"ff",	--13589
		x"ff",	--13590
		x"ff",	--13591
		x"ff",	--13592
		x"ff",	--13593
		x"ff",	--13594
		x"ff",	--13595
		x"ff",	--13596
		x"ff",	--13597
		x"ff",	--13598
		x"ff",	--13599
		x"ff",	--13600
		x"ff",	--13601
		x"ff",	--13602
		x"ff",	--13603
		x"ff",	--13604
		x"ff",	--13605
		x"ff",	--13606
		x"ff",	--13607
		x"ff",	--13608
		x"ff",	--13609
		x"ff",	--13610
		x"ff",	--13611
		x"ff",	--13612
		x"ff",	--13613
		x"ff",	--13614
		x"ff",	--13615
		x"ff",	--13616
		x"ff",	--13617
		x"ff",	--13618
		x"ff",	--13619
		x"ff",	--13620
		x"ff",	--13621
		x"ff",	--13622
		x"ff",	--13623
		x"ff",	--13624
		x"ff",	--13625
		x"ff",	--13626
		x"ff",	--13627
		x"ff",	--13628
		x"ff",	--13629
		x"ff",	--13630
		x"ff",	--13631
		x"ff",	--13632
		x"ff",	--13633
		x"ff",	--13634
		x"ff",	--13635
		x"ff",	--13636
		x"ff",	--13637
		x"ff",	--13638
		x"ff",	--13639
		x"ff",	--13640
		x"ff",	--13641
		x"ff",	--13642
		x"ff",	--13643
		x"ff",	--13644
		x"ff",	--13645
		x"ff",	--13646
		x"ff",	--13647
		x"ff",	--13648
		x"ff",	--13649
		x"ff",	--13650
		x"ff",	--13651
		x"ff",	--13652
		x"ff",	--13653
		x"ff",	--13654
		x"ff",	--13655
		x"ff",	--13656
		x"ff",	--13657
		x"ff",	--13658
		x"ff",	--13659
		x"ff",	--13660
		x"ff",	--13661
		x"ff",	--13662
		x"ff",	--13663
		x"ff",	--13664
		x"ff",	--13665
		x"ff",	--13666
		x"ff",	--13667
		x"ff",	--13668
		x"ff",	--13669
		x"ff",	--13670
		x"ff",	--13671
		x"ff",	--13672
		x"ff",	--13673
		x"ff",	--13674
		x"ff",	--13675
		x"ff",	--13676
		x"ff",	--13677
		x"ff",	--13678
		x"ff",	--13679
		x"ff",	--13680
		x"ff",	--13681
		x"ff",	--13682
		x"ff",	--13683
		x"ff",	--13684
		x"ff",	--13685
		x"ff",	--13686
		x"ff",	--13687
		x"ff",	--13688
		x"ff",	--13689
		x"ff",	--13690
		x"ff",	--13691
		x"ff",	--13692
		x"ff",	--13693
		x"ff",	--13694
		x"ff",	--13695
		x"ff",	--13696
		x"ff",	--13697
		x"ff",	--13698
		x"ff",	--13699
		x"ff",	--13700
		x"ff",	--13701
		x"ff",	--13702
		x"ff",	--13703
		x"ff",	--13704
		x"ff",	--13705
		x"ff",	--13706
		x"ff",	--13707
		x"ff",	--13708
		x"ff",	--13709
		x"ff",	--13710
		x"ff",	--13711
		x"ff",	--13712
		x"ff",	--13713
		x"ff",	--13714
		x"ff",	--13715
		x"ff",	--13716
		x"ff",	--13717
		x"ff",	--13718
		x"ff",	--13719
		x"ff",	--13720
		x"ff",	--13721
		x"ff",	--13722
		x"ff",	--13723
		x"ff",	--13724
		x"ff",	--13725
		x"ff",	--13726
		x"ff",	--13727
		x"ff",	--13728
		x"ff",	--13729
		x"ff",	--13730
		x"ff",	--13731
		x"ff",	--13732
		x"ff",	--13733
		x"ff",	--13734
		x"ff",	--13735
		x"ff",	--13736
		x"ff",	--13737
		x"ff",	--13738
		x"ff",	--13739
		x"ff",	--13740
		x"ff",	--13741
		x"ff",	--13742
		x"ff",	--13743
		x"ff",	--13744
		x"ff",	--13745
		x"ff",	--13746
		x"ff",	--13747
		x"ff",	--13748
		x"ff",	--13749
		x"ff",	--13750
		x"ff",	--13751
		x"ff",	--13752
		x"ff",	--13753
		x"ff",	--13754
		x"ff",	--13755
		x"ff",	--13756
		x"ff",	--13757
		x"ff",	--13758
		x"ff",	--13759
		x"ff",	--13760
		x"ff",	--13761
		x"ff",	--13762
		x"ff",	--13763
		x"ff",	--13764
		x"ff",	--13765
		x"ff",	--13766
		x"ff",	--13767
		x"ff",	--13768
		x"ff",	--13769
		x"ff",	--13770
		x"ff",	--13771
		x"ff",	--13772
		x"ff",	--13773
		x"ff",	--13774
		x"ff",	--13775
		x"ff",	--13776
		x"ff",	--13777
		x"ff",	--13778
		x"ff",	--13779
		x"ff",	--13780
		x"ff",	--13781
		x"ff",	--13782
		x"ff",	--13783
		x"ff",	--13784
		x"ff",	--13785
		x"ff",	--13786
		x"ff",	--13787
		x"ff",	--13788
		x"ff",	--13789
		x"ff",	--13790
		x"ff",	--13791
		x"ff",	--13792
		x"ff",	--13793
		x"ff",	--13794
		x"ff",	--13795
		x"ff",	--13796
		x"ff",	--13797
		x"ff",	--13798
		x"ff",	--13799
		x"ff",	--13800
		x"ff",	--13801
		x"ff",	--13802
		x"ff",	--13803
		x"ff",	--13804
		x"ff",	--13805
		x"ff",	--13806
		x"ff",	--13807
		x"ff",	--13808
		x"ff",	--13809
		x"ff",	--13810
		x"ff",	--13811
		x"ff",	--13812
		x"ff",	--13813
		x"ff",	--13814
		x"ff",	--13815
		x"ff",	--13816
		x"ff",	--13817
		x"ff",	--13818
		x"ff",	--13819
		x"ff",	--13820
		x"ff",	--13821
		x"ff",	--13822
		x"ff",	--13823
		x"ff",	--13824
		x"ff",	--13825
		x"ff",	--13826
		x"ff",	--13827
		x"ff",	--13828
		x"ff",	--13829
		x"ff",	--13830
		x"ff",	--13831
		x"ff",	--13832
		x"ff",	--13833
		x"ff",	--13834
		x"ff",	--13835
		x"ff",	--13836
		x"ff",	--13837
		x"ff",	--13838
		x"ff",	--13839
		x"ff",	--13840
		x"ff",	--13841
		x"ff",	--13842
		x"ff",	--13843
		x"ff",	--13844
		x"ff",	--13845
		x"ff",	--13846
		x"ff",	--13847
		x"ff",	--13848
		x"ff",	--13849
		x"ff",	--13850
		x"ff",	--13851
		x"ff",	--13852
		x"ff",	--13853
		x"ff",	--13854
		x"ff",	--13855
		x"ff",	--13856
		x"ff",	--13857
		x"ff",	--13858
		x"ff",	--13859
		x"ff",	--13860
		x"ff",	--13861
		x"ff",	--13862
		x"ff",	--13863
		x"ff",	--13864
		x"ff",	--13865
		x"ff",	--13866
		x"ff",	--13867
		x"ff",	--13868
		x"ff",	--13869
		x"ff",	--13870
		x"ff",	--13871
		x"ff",	--13872
		x"ff",	--13873
		x"ff",	--13874
		x"ff",	--13875
		x"ff",	--13876
		x"ff",	--13877
		x"ff",	--13878
		x"ff",	--13879
		x"ff",	--13880
		x"ff",	--13881
		x"ff",	--13882
		x"ff",	--13883
		x"ff",	--13884
		x"ff",	--13885
		x"ff",	--13886
		x"ff",	--13887
		x"ff",	--13888
		x"ff",	--13889
		x"ff",	--13890
		x"ff",	--13891
		x"ff",	--13892
		x"ff",	--13893
		x"ff",	--13894
		x"ff",	--13895
		x"ff",	--13896
		x"ff",	--13897
		x"ff",	--13898
		x"ff",	--13899
		x"ff",	--13900
		x"ff",	--13901
		x"ff",	--13902
		x"ff",	--13903
		x"ff",	--13904
		x"ff",	--13905
		x"ff",	--13906
		x"ff",	--13907
		x"ff",	--13908
		x"ff",	--13909
		x"ff",	--13910
		x"ff",	--13911
		x"ff",	--13912
		x"ff",	--13913
		x"ff",	--13914
		x"ff",	--13915
		x"ff",	--13916
		x"ff",	--13917
		x"ff",	--13918
		x"ff",	--13919
		x"ff",	--13920
		x"ff",	--13921
		x"ff",	--13922
		x"ff",	--13923
		x"ff",	--13924
		x"ff",	--13925
		x"ff",	--13926
		x"ff",	--13927
		x"ff",	--13928
		x"ff",	--13929
		x"ff",	--13930
		x"ff",	--13931
		x"ff",	--13932
		x"ff",	--13933
		x"ff",	--13934
		x"ff",	--13935
		x"ff",	--13936
		x"ff",	--13937
		x"ff",	--13938
		x"ff",	--13939
		x"ff",	--13940
		x"ff",	--13941
		x"ff",	--13942
		x"ff",	--13943
		x"ff",	--13944
		x"ff",	--13945
		x"ff",	--13946
		x"ff",	--13947
		x"ff",	--13948
		x"ff",	--13949
		x"ff",	--13950
		x"ff",	--13951
		x"ff",	--13952
		x"ff",	--13953
		x"ff",	--13954
		x"ff",	--13955
		x"ff",	--13956
		x"ff",	--13957
		x"ff",	--13958
		x"ff",	--13959
		x"ff",	--13960
		x"ff",	--13961
		x"ff",	--13962
		x"ff",	--13963
		x"ff",	--13964
		x"ff",	--13965
		x"ff",	--13966
		x"ff",	--13967
		x"ff",	--13968
		x"ff",	--13969
		x"ff",	--13970
		x"ff",	--13971
		x"ff",	--13972
		x"ff",	--13973
		x"ff",	--13974
		x"ff",	--13975
		x"ff",	--13976
		x"ff",	--13977
		x"ff",	--13978
		x"ff",	--13979
		x"ff",	--13980
		x"ff",	--13981
		x"ff",	--13982
		x"ff",	--13983
		x"ff",	--13984
		x"ff",	--13985
		x"ff",	--13986
		x"ff",	--13987
		x"ff",	--13988
		x"ff",	--13989
		x"ff",	--13990
		x"ff",	--13991
		x"ff",	--13992
		x"ff",	--13993
		x"ff",	--13994
		x"ff",	--13995
		x"ff",	--13996
		x"ff",	--13997
		x"ff",	--13998
		x"ff",	--13999
		x"ff",	--14000
		x"ff",	--14001
		x"ff",	--14002
		x"ff",	--14003
		x"ff",	--14004
		x"ff",	--14005
		x"ff",	--14006
		x"ff",	--14007
		x"ff",	--14008
		x"ff",	--14009
		x"ff",	--14010
		x"ff",	--14011
		x"ff",	--14012
		x"ff",	--14013
		x"ff",	--14014
		x"ff",	--14015
		x"ff",	--14016
		x"ff",	--14017
		x"ff",	--14018
		x"ff",	--14019
		x"ff",	--14020
		x"ff",	--14021
		x"ff",	--14022
		x"ff",	--14023
		x"ff",	--14024
		x"ff",	--14025
		x"ff",	--14026
		x"ff",	--14027
		x"ff",	--14028
		x"ff",	--14029
		x"ff",	--14030
		x"ff",	--14031
		x"ff",	--14032
		x"ff",	--14033
		x"ff",	--14034
		x"ff",	--14035
		x"ff",	--14036
		x"ff",	--14037
		x"ff",	--14038
		x"ff",	--14039
		x"ff",	--14040
		x"ff",	--14041
		x"ff",	--14042
		x"ff",	--14043
		x"ff",	--14044
		x"ff",	--14045
		x"ff",	--14046
		x"ff",	--14047
		x"ff",	--14048
		x"ff",	--14049
		x"ff",	--14050
		x"ff",	--14051
		x"ff",	--14052
		x"ff",	--14053
		x"ff",	--14054
		x"ff",	--14055
		x"ff",	--14056
		x"ff",	--14057
		x"ff",	--14058
		x"ff",	--14059
		x"ff",	--14060
		x"ff",	--14061
		x"ff",	--14062
		x"ff",	--14063
		x"ff",	--14064
		x"ff",	--14065
		x"ff",	--14066
		x"ff",	--14067
		x"ff",	--14068
		x"ff",	--14069
		x"ff",	--14070
		x"ff",	--14071
		x"ff",	--14072
		x"ff",	--14073
		x"ff",	--14074
		x"ff",	--14075
		x"ff",	--14076
		x"ff",	--14077
		x"ff",	--14078
		x"ff",	--14079
		x"ff",	--14080
		x"ff",	--14081
		x"ff",	--14082
		x"ff",	--14083
		x"ff",	--14084
		x"ff",	--14085
		x"ff",	--14086
		x"ff",	--14087
		x"ff",	--14088
		x"ff",	--14089
		x"ff",	--14090
		x"ff",	--14091
		x"ff",	--14092
		x"ff",	--14093
		x"ff",	--14094
		x"ff",	--14095
		x"ff",	--14096
		x"ff",	--14097
		x"ff",	--14098
		x"ff",	--14099
		x"ff",	--14100
		x"ff",	--14101
		x"ff",	--14102
		x"ff",	--14103
		x"ff",	--14104
		x"ff",	--14105
		x"ff",	--14106
		x"ff",	--14107
		x"ff",	--14108
		x"ff",	--14109
		x"ff",	--14110
		x"ff",	--14111
		x"ff",	--14112
		x"ff",	--14113
		x"ff",	--14114
		x"ff",	--14115
		x"ff",	--14116
		x"ff",	--14117
		x"ff",	--14118
		x"ff",	--14119
		x"ff",	--14120
		x"ff",	--14121
		x"ff",	--14122
		x"ff",	--14123
		x"ff",	--14124
		x"ff",	--14125
		x"ff",	--14126
		x"ff",	--14127
		x"ff",	--14128
		x"ff",	--14129
		x"ff",	--14130
		x"ff",	--14131
		x"ff",	--14132
		x"ff",	--14133
		x"ff",	--14134
		x"ff",	--14135
		x"ff",	--14136
		x"ff",	--14137
		x"ff",	--14138
		x"ff",	--14139
		x"ff",	--14140
		x"ff",	--14141
		x"ff",	--14142
		x"ff",	--14143
		x"ff",	--14144
		x"ff",	--14145
		x"ff",	--14146
		x"ff",	--14147
		x"ff",	--14148
		x"ff",	--14149
		x"ff",	--14150
		x"ff",	--14151
		x"ff",	--14152
		x"ff",	--14153
		x"ff",	--14154
		x"ff",	--14155
		x"ff",	--14156
		x"ff",	--14157
		x"ff",	--14158
		x"ff",	--14159
		x"ff",	--14160
		x"ff",	--14161
		x"ff",	--14162
		x"ff",	--14163
		x"ff",	--14164
		x"ff",	--14165
		x"ff",	--14166
		x"ff",	--14167
		x"ff",	--14168
		x"ff",	--14169
		x"ff",	--14170
		x"ff",	--14171
		x"ff",	--14172
		x"ff",	--14173
		x"ff",	--14174
		x"ff",	--14175
		x"ff",	--14176
		x"ff",	--14177
		x"ff",	--14178
		x"ff",	--14179
		x"ff",	--14180
		x"ff",	--14181
		x"ff",	--14182
		x"ff",	--14183
		x"ff",	--14184
		x"ff",	--14185
		x"ff",	--14186
		x"ff",	--14187
		x"ff",	--14188
		x"ff",	--14189
		x"ff",	--14190
		x"ff",	--14191
		x"ff",	--14192
		x"ff",	--14193
		x"ff",	--14194
		x"ff",	--14195
		x"ff",	--14196
		x"ff",	--14197
		x"ff",	--14198
		x"ff",	--14199
		x"ff",	--14200
		x"ff",	--14201
		x"ff",	--14202
		x"ff",	--14203
		x"ff",	--14204
		x"ff",	--14205
		x"ff",	--14206
		x"ff",	--14207
		x"ff",	--14208
		x"ff",	--14209
		x"ff",	--14210
		x"ff",	--14211
		x"ff",	--14212
		x"ff",	--14213
		x"ff",	--14214
		x"ff",	--14215
		x"ff",	--14216
		x"ff",	--14217
		x"ff",	--14218
		x"ff",	--14219
		x"ff",	--14220
		x"ff",	--14221
		x"ff",	--14222
		x"ff",	--14223
		x"ff",	--14224
		x"ff",	--14225
		x"ff",	--14226
		x"ff",	--14227
		x"ff",	--14228
		x"ff",	--14229
		x"ff",	--14230
		x"ff",	--14231
		x"ff",	--14232
		x"ff",	--14233
		x"ff",	--14234
		x"ff",	--14235
		x"ff",	--14236
		x"ff",	--14237
		x"ff",	--14238
		x"ff",	--14239
		x"ff",	--14240
		x"ff",	--14241
		x"ff",	--14242
		x"ff",	--14243
		x"ff",	--14244
		x"ff",	--14245
		x"ff",	--14246
		x"ff",	--14247
		x"ff",	--14248
		x"ff",	--14249
		x"ff",	--14250
		x"ff",	--14251
		x"ff",	--14252
		x"ff",	--14253
		x"ff",	--14254
		x"ff",	--14255
		x"ff",	--14256
		x"ff",	--14257
		x"ff",	--14258
		x"ff",	--14259
		x"ff",	--14260
		x"ff",	--14261
		x"ff",	--14262
		x"ff",	--14263
		x"ff",	--14264
		x"ff",	--14265
		x"ff",	--14266
		x"ff",	--14267
		x"ff",	--14268
		x"ff",	--14269
		x"ff",	--14270
		x"ff",	--14271
		x"ff",	--14272
		x"ff",	--14273
		x"ff",	--14274
		x"ff",	--14275
		x"ff",	--14276
		x"ff",	--14277
		x"ff",	--14278
		x"ff",	--14279
		x"ff",	--14280
		x"ff",	--14281
		x"ff",	--14282
		x"ff",	--14283
		x"ff",	--14284
		x"ff",	--14285
		x"ff",	--14286
		x"ff",	--14287
		x"ff",	--14288
		x"ff",	--14289
		x"ff",	--14290
		x"ff",	--14291
		x"ff",	--14292
		x"ff",	--14293
		x"ff",	--14294
		x"ff",	--14295
		x"ff",	--14296
		x"ff",	--14297
		x"ff",	--14298
		x"ff",	--14299
		x"ff",	--14300
		x"ff",	--14301
		x"ff",	--14302
		x"ff",	--14303
		x"ff",	--14304
		x"ff",	--14305
		x"ff",	--14306
		x"ff",	--14307
		x"ff",	--14308
		x"ff",	--14309
		x"ff",	--14310
		x"ff",	--14311
		x"ff",	--14312
		x"ff",	--14313
		x"ff",	--14314
		x"ff",	--14315
		x"ff",	--14316
		x"ff",	--14317
		x"ff",	--14318
		x"ff",	--14319
		x"ff",	--14320
		x"ff",	--14321
		x"ff",	--14322
		x"ff",	--14323
		x"ff",	--14324
		x"ff",	--14325
		x"ff",	--14326
		x"ff",	--14327
		x"ff",	--14328
		x"ff",	--14329
		x"ff",	--14330
		x"ff",	--14331
		x"ff",	--14332
		x"ff",	--14333
		x"ff",	--14334
		x"ff",	--14335
		x"ff",	--14336
		x"ff",	--14337
		x"ff",	--14338
		x"ff",	--14339
		x"ff",	--14340
		x"ff",	--14341
		x"ff",	--14342
		x"ff",	--14343
		x"ff",	--14344
		x"ff",	--14345
		x"ff",	--14346
		x"ff",	--14347
		x"ff",	--14348
		x"ff",	--14349
		x"ff",	--14350
		x"ff",	--14351
		x"ff",	--14352
		x"ff",	--14353
		x"ff",	--14354
		x"ff",	--14355
		x"ff",	--14356
		x"ff",	--14357
		x"ff",	--14358
		x"ff",	--14359
		x"ff",	--14360
		x"ff",	--14361
		x"ff",	--14362
		x"ff",	--14363
		x"ff",	--14364
		x"ff",	--14365
		x"ff",	--14366
		x"ff",	--14367
		x"ff",	--14368
		x"ff",	--14369
		x"ff",	--14370
		x"ff",	--14371
		x"ff",	--14372
		x"ff",	--14373
		x"ff",	--14374
		x"ff",	--14375
		x"ff",	--14376
		x"ff",	--14377
		x"ff",	--14378
		x"ff",	--14379
		x"ff",	--14380
		x"ff",	--14381
		x"ff",	--14382
		x"ff",	--14383
		x"ff",	--14384
		x"ff",	--14385
		x"ff",	--14386
		x"ff",	--14387
		x"ff",	--14388
		x"ff",	--14389
		x"ff",	--14390
		x"ff",	--14391
		x"ff",	--14392
		x"ff",	--14393
		x"ff",	--14394
		x"ff",	--14395
		x"ff",	--14396
		x"ff",	--14397
		x"ff",	--14398
		x"ff",	--14399
		x"ff",	--14400
		x"ff",	--14401
		x"ff",	--14402
		x"ff",	--14403
		x"ff",	--14404
		x"ff",	--14405
		x"ff",	--14406
		x"ff",	--14407
		x"ff",	--14408
		x"ff",	--14409
		x"ff",	--14410
		x"ff",	--14411
		x"ff",	--14412
		x"ff",	--14413
		x"ff",	--14414
		x"ff",	--14415
		x"ff",	--14416
		x"ff",	--14417
		x"ff",	--14418
		x"ff",	--14419
		x"ff",	--14420
		x"ff",	--14421
		x"ff",	--14422
		x"ff",	--14423
		x"ff",	--14424
		x"ff",	--14425
		x"ff",	--14426
		x"ff",	--14427
		x"ff",	--14428
		x"ff",	--14429
		x"ff",	--14430
		x"ff",	--14431
		x"ff",	--14432
		x"ff",	--14433
		x"ff",	--14434
		x"ff",	--14435
		x"ff",	--14436
		x"ff",	--14437
		x"ff",	--14438
		x"ff",	--14439
		x"ff",	--14440
		x"ff",	--14441
		x"ff",	--14442
		x"ff",	--14443
		x"ff",	--14444
		x"ff",	--14445
		x"ff",	--14446
		x"ff",	--14447
		x"ff",	--14448
		x"ff",	--14449
		x"ff",	--14450
		x"ff",	--14451
		x"ff",	--14452
		x"ff",	--14453
		x"ff",	--14454
		x"ff",	--14455
		x"ff",	--14456
		x"ff",	--14457
		x"ff",	--14458
		x"ff",	--14459
		x"ff",	--14460
		x"ff",	--14461
		x"ff",	--14462
		x"ff",	--14463
		x"ff",	--14464
		x"ff",	--14465
		x"ff",	--14466
		x"ff",	--14467
		x"ff",	--14468
		x"ff",	--14469
		x"ff",	--14470
		x"ff",	--14471
		x"ff",	--14472
		x"ff",	--14473
		x"ff",	--14474
		x"ff",	--14475
		x"ff",	--14476
		x"ff",	--14477
		x"ff",	--14478
		x"ff",	--14479
		x"ff",	--14480
		x"ff",	--14481
		x"ff",	--14482
		x"ff",	--14483
		x"ff",	--14484
		x"ff",	--14485
		x"ff",	--14486
		x"ff",	--14487
		x"ff",	--14488
		x"ff",	--14489
		x"ff",	--14490
		x"ff",	--14491
		x"ff",	--14492
		x"ff",	--14493
		x"ff",	--14494
		x"ff",	--14495
		x"ff",	--14496
		x"ff",	--14497
		x"ff",	--14498
		x"ff",	--14499
		x"ff",	--14500
		x"ff",	--14501
		x"ff",	--14502
		x"ff",	--14503
		x"ff",	--14504
		x"ff",	--14505
		x"ff",	--14506
		x"ff",	--14507
		x"ff",	--14508
		x"ff",	--14509
		x"ff",	--14510
		x"ff",	--14511
		x"ff",	--14512
		x"ff",	--14513
		x"ff",	--14514
		x"ff",	--14515
		x"ff",	--14516
		x"ff",	--14517
		x"ff",	--14518
		x"ff",	--14519
		x"ff",	--14520
		x"ff",	--14521
		x"ff",	--14522
		x"ff",	--14523
		x"ff",	--14524
		x"ff",	--14525
		x"ff",	--14526
		x"ff",	--14527
		x"ff",	--14528
		x"ff",	--14529
		x"ff",	--14530
		x"ff",	--14531
		x"ff",	--14532
		x"ff",	--14533
		x"ff",	--14534
		x"ff",	--14535
		x"ff",	--14536
		x"ff",	--14537
		x"ff",	--14538
		x"ff",	--14539
		x"ff",	--14540
		x"ff",	--14541
		x"ff",	--14542
		x"ff",	--14543
		x"ff",	--14544
		x"ff",	--14545
		x"ff",	--14546
		x"ff",	--14547
		x"ff",	--14548
		x"ff",	--14549
		x"ff",	--14550
		x"ff",	--14551
		x"ff",	--14552
		x"ff",	--14553
		x"ff",	--14554
		x"ff",	--14555
		x"ff",	--14556
		x"ff",	--14557
		x"ff",	--14558
		x"ff",	--14559
		x"ff",	--14560
		x"ff",	--14561
		x"ff",	--14562
		x"ff",	--14563
		x"ff",	--14564
		x"ff",	--14565
		x"ff",	--14566
		x"ff",	--14567
		x"ff",	--14568
		x"ff",	--14569
		x"ff",	--14570
		x"ff",	--14571
		x"ff",	--14572
		x"ff",	--14573
		x"ff",	--14574
		x"ff",	--14575
		x"ff",	--14576
		x"ff",	--14577
		x"ff",	--14578
		x"ff",	--14579
		x"ff",	--14580
		x"ff",	--14581
		x"ff",	--14582
		x"ff",	--14583
		x"ff",	--14584
		x"ff",	--14585
		x"ff",	--14586
		x"ff",	--14587
		x"ff",	--14588
		x"ff",	--14589
		x"ff",	--14590
		x"ff",	--14591
		x"ff",	--14592
		x"ff",	--14593
		x"ff",	--14594
		x"ff",	--14595
		x"ff",	--14596
		x"ff",	--14597
		x"ff",	--14598
		x"ff",	--14599
		x"ff",	--14600
		x"ff",	--14601
		x"ff",	--14602
		x"ff",	--14603
		x"ff",	--14604
		x"ff",	--14605
		x"ff",	--14606
		x"ff",	--14607
		x"ff",	--14608
		x"ff",	--14609
		x"ff",	--14610
		x"ff",	--14611
		x"ff",	--14612
		x"ff",	--14613
		x"ff",	--14614
		x"ff",	--14615
		x"ff",	--14616
		x"ff",	--14617
		x"ff",	--14618
		x"ff",	--14619
		x"ff",	--14620
		x"ff",	--14621
		x"ff",	--14622
		x"ff",	--14623
		x"ff",	--14624
		x"ff",	--14625
		x"ff",	--14626
		x"ff",	--14627
		x"ff",	--14628
		x"ff",	--14629
		x"ff",	--14630
		x"ff",	--14631
		x"ff",	--14632
		x"ff",	--14633
		x"ff",	--14634
		x"ff",	--14635
		x"ff",	--14636
		x"ff",	--14637
		x"ff",	--14638
		x"ff",	--14639
		x"ff",	--14640
		x"ff",	--14641
		x"ff",	--14642
		x"ff",	--14643
		x"ff",	--14644
		x"ff",	--14645
		x"ff",	--14646
		x"ff",	--14647
		x"ff",	--14648
		x"ff",	--14649
		x"ff",	--14650
		x"ff",	--14651
		x"ff",	--14652
		x"ff",	--14653
		x"ff",	--14654
		x"ff",	--14655
		x"ff",	--14656
		x"ff",	--14657
		x"ff",	--14658
		x"ff",	--14659
		x"ff",	--14660
		x"ff",	--14661
		x"ff",	--14662
		x"ff",	--14663
		x"ff",	--14664
		x"ff",	--14665
		x"ff",	--14666
		x"ff",	--14667
		x"ff",	--14668
		x"ff",	--14669
		x"ff",	--14670
		x"ff",	--14671
		x"ff",	--14672
		x"ff",	--14673
		x"ff",	--14674
		x"ff",	--14675
		x"ff",	--14676
		x"ff",	--14677
		x"ff",	--14678
		x"ff",	--14679
		x"ff",	--14680
		x"ff",	--14681
		x"ff",	--14682
		x"ff",	--14683
		x"ff",	--14684
		x"ff",	--14685
		x"ff",	--14686
		x"ff",	--14687
		x"ff",	--14688
		x"ff",	--14689
		x"ff",	--14690
		x"ff",	--14691
		x"ff",	--14692
		x"ff",	--14693
		x"ff",	--14694
		x"ff",	--14695
		x"ff",	--14696
		x"ff",	--14697
		x"ff",	--14698
		x"ff",	--14699
		x"ff",	--14700
		x"ff",	--14701
		x"ff",	--14702
		x"ff",	--14703
		x"ff",	--14704
		x"ff",	--14705
		x"ff",	--14706
		x"ff",	--14707
		x"ff",	--14708
		x"ff",	--14709
		x"ff",	--14710
		x"ff",	--14711
		x"ff",	--14712
		x"ff",	--14713
		x"ff",	--14714
		x"ff",	--14715
		x"ff",	--14716
		x"ff",	--14717
		x"ff",	--14718
		x"ff",	--14719
		x"ff",	--14720
		x"ff",	--14721
		x"ff",	--14722
		x"ff",	--14723
		x"ff",	--14724
		x"ff",	--14725
		x"ff",	--14726
		x"ff",	--14727
		x"ff",	--14728
		x"ff",	--14729
		x"ff",	--14730
		x"ff",	--14731
		x"ff",	--14732
		x"ff",	--14733
		x"ff",	--14734
		x"ff",	--14735
		x"ff",	--14736
		x"ff",	--14737
		x"ff",	--14738
		x"ff",	--14739
		x"ff",	--14740
		x"ff",	--14741
		x"ff",	--14742
		x"ff",	--14743
		x"ff",	--14744
		x"ff",	--14745
		x"ff",	--14746
		x"ff",	--14747
		x"ff",	--14748
		x"ff",	--14749
		x"ff",	--14750
		x"ff",	--14751
		x"ff",	--14752
		x"ff",	--14753
		x"ff",	--14754
		x"ff",	--14755
		x"ff",	--14756
		x"ff",	--14757
		x"ff",	--14758
		x"ff",	--14759
		x"ff",	--14760
		x"ff",	--14761
		x"ff",	--14762
		x"ff",	--14763
		x"ff",	--14764
		x"ff",	--14765
		x"ff",	--14766
		x"ff",	--14767
		x"ff",	--14768
		x"ff",	--14769
		x"ff",	--14770
		x"ff",	--14771
		x"ff",	--14772
		x"ff",	--14773
		x"ff",	--14774
		x"ff",	--14775
		x"ff",	--14776
		x"ff",	--14777
		x"ff",	--14778
		x"ff",	--14779
		x"ff",	--14780
		x"ff",	--14781
		x"ff",	--14782
		x"ff",	--14783
		x"ff",	--14784
		x"ff",	--14785
		x"ff",	--14786
		x"ff",	--14787
		x"ff",	--14788
		x"ff",	--14789
		x"ff",	--14790
		x"ff",	--14791
		x"ff",	--14792
		x"ff",	--14793
		x"ff",	--14794
		x"ff",	--14795
		x"ff",	--14796
		x"ff",	--14797
		x"ff",	--14798
		x"ff",	--14799
		x"ff",	--14800
		x"ff",	--14801
		x"ff",	--14802
		x"ff",	--14803
		x"ff",	--14804
		x"ff",	--14805
		x"ff",	--14806
		x"ff",	--14807
		x"ff",	--14808
		x"ff",	--14809
		x"ff",	--14810
		x"ff",	--14811
		x"ff",	--14812
		x"ff",	--14813
		x"ff",	--14814
		x"ff",	--14815
		x"ff",	--14816
		x"ff",	--14817
		x"ff",	--14818
		x"ff",	--14819
		x"ff",	--14820
		x"ff",	--14821
		x"ff",	--14822
		x"ff",	--14823
		x"ff",	--14824
		x"ff",	--14825
		x"ff",	--14826
		x"ff",	--14827
		x"ff",	--14828
		x"ff",	--14829
		x"ff",	--14830
		x"ff",	--14831
		x"ff",	--14832
		x"ff",	--14833
		x"ff",	--14834
		x"ff",	--14835
		x"ff",	--14836
		x"ff",	--14837
		x"ff",	--14838
		x"ff",	--14839
		x"ff",	--14840
		x"ff",	--14841
		x"ff",	--14842
		x"ff",	--14843
		x"ff",	--14844
		x"ff",	--14845
		x"ff",	--14846
		x"ff",	--14847
		x"ff",	--14848
		x"ff",	--14849
		x"ff",	--14850
		x"ff",	--14851
		x"ff",	--14852
		x"ff",	--14853
		x"ff",	--14854
		x"ff",	--14855
		x"ff",	--14856
		x"ff",	--14857
		x"ff",	--14858
		x"ff",	--14859
		x"ff",	--14860
		x"ff",	--14861
		x"ff",	--14862
		x"ff",	--14863
		x"ff",	--14864
		x"ff",	--14865
		x"ff",	--14866
		x"ff",	--14867
		x"ff",	--14868
		x"ff",	--14869
		x"ff",	--14870
		x"ff",	--14871
		x"ff",	--14872
		x"ff",	--14873
		x"ff",	--14874
		x"ff",	--14875
		x"ff",	--14876
		x"ff",	--14877
		x"ff",	--14878
		x"ff",	--14879
		x"ff",	--14880
		x"ff",	--14881
		x"ff",	--14882
		x"ff",	--14883
		x"ff",	--14884
		x"ff",	--14885
		x"ff",	--14886
		x"ff",	--14887
		x"ff",	--14888
		x"ff",	--14889
		x"ff",	--14890
		x"ff",	--14891
		x"ff",	--14892
		x"ff",	--14893
		x"ff",	--14894
		x"ff",	--14895
		x"ff",	--14896
		x"ff",	--14897
		x"ff",	--14898
		x"ff",	--14899
		x"ff",	--14900
		x"ff",	--14901
		x"ff",	--14902
		x"ff",	--14903
		x"ff",	--14904
		x"ff",	--14905
		x"ff",	--14906
		x"ff",	--14907
		x"ff",	--14908
		x"ff",	--14909
		x"ff",	--14910
		x"ff",	--14911
		x"ff",	--14912
		x"ff",	--14913
		x"ff",	--14914
		x"ff",	--14915
		x"ff",	--14916
		x"ff",	--14917
		x"ff",	--14918
		x"ff",	--14919
		x"ff",	--14920
		x"ff",	--14921
		x"ff",	--14922
		x"ff",	--14923
		x"ff",	--14924
		x"ff",	--14925
		x"ff",	--14926
		x"ff",	--14927
		x"ff",	--14928
		x"ff",	--14929
		x"ff",	--14930
		x"ff",	--14931
		x"ff",	--14932
		x"ff",	--14933
		x"ff",	--14934
		x"ff",	--14935
		x"ff",	--14936
		x"ff",	--14937
		x"ff",	--14938
		x"ff",	--14939
		x"ff",	--14940
		x"ff",	--14941
		x"ff",	--14942
		x"ff",	--14943
		x"ff",	--14944
		x"ff",	--14945
		x"ff",	--14946
		x"ff",	--14947
		x"ff",	--14948
		x"ff",	--14949
		x"ff",	--14950
		x"ff",	--14951
		x"ff",	--14952
		x"ff",	--14953
		x"ff",	--14954
		x"ff",	--14955
		x"ff",	--14956
		x"ff",	--14957
		x"ff",	--14958
		x"ff",	--14959
		x"ff",	--14960
		x"ff",	--14961
		x"ff",	--14962
		x"ff",	--14963
		x"ff",	--14964
		x"ff",	--14965
		x"ff",	--14966
		x"ff",	--14967
		x"ff",	--14968
		x"ff",	--14969
		x"ff",	--14970
		x"ff",	--14971
		x"ff",	--14972
		x"ff",	--14973
		x"ff",	--14974
		x"ff",	--14975
		x"ff",	--14976
		x"ff",	--14977
		x"ff",	--14978
		x"ff",	--14979
		x"ff",	--14980
		x"ff",	--14981
		x"ff",	--14982
		x"ff",	--14983
		x"ff",	--14984
		x"ff",	--14985
		x"ff",	--14986
		x"ff",	--14987
		x"ff",	--14988
		x"ff",	--14989
		x"ff",	--14990
		x"ff",	--14991
		x"ff",	--14992
		x"ff",	--14993
		x"ff",	--14994
		x"ff",	--14995
		x"ff",	--14996
		x"ff",	--14997
		x"ff",	--14998
		x"ff",	--14999
		x"ff",	--15000
		x"ff",	--15001
		x"ff",	--15002
		x"ff",	--15003
		x"ff",	--15004
		x"ff",	--15005
		x"ff",	--15006
		x"ff",	--15007
		x"ff",	--15008
		x"ff",	--15009
		x"ff",	--15010
		x"ff",	--15011
		x"ff",	--15012
		x"ff",	--15013
		x"ff",	--15014
		x"ff",	--15015
		x"ff",	--15016
		x"ff",	--15017
		x"ff",	--15018
		x"ff",	--15019
		x"ff",	--15020
		x"ff",	--15021
		x"ff",	--15022
		x"ff",	--15023
		x"ff",	--15024
		x"ff",	--15025
		x"ff",	--15026
		x"ff",	--15027
		x"ff",	--15028
		x"ff",	--15029
		x"ff",	--15030
		x"ff",	--15031
		x"ff",	--15032
		x"ff",	--15033
		x"ff",	--15034
		x"ff",	--15035
		x"ff",	--15036
		x"ff",	--15037
		x"ff",	--15038
		x"ff",	--15039
		x"ff",	--15040
		x"ff",	--15041
		x"ff",	--15042
		x"ff",	--15043
		x"ff",	--15044
		x"ff",	--15045
		x"ff",	--15046
		x"ff",	--15047
		x"ff",	--15048
		x"ff",	--15049
		x"ff",	--15050
		x"ff",	--15051
		x"ff",	--15052
		x"ff",	--15053
		x"ff",	--15054
		x"ff",	--15055
		x"ff",	--15056
		x"ff",	--15057
		x"ff",	--15058
		x"ff",	--15059
		x"ff",	--15060
		x"ff",	--15061
		x"ff",	--15062
		x"ff",	--15063
		x"ff",	--15064
		x"ff",	--15065
		x"ff",	--15066
		x"ff",	--15067
		x"ff",	--15068
		x"ff",	--15069
		x"ff",	--15070
		x"ff",	--15071
		x"ff",	--15072
		x"ff",	--15073
		x"ff",	--15074
		x"ff",	--15075
		x"ff",	--15076
		x"ff",	--15077
		x"ff",	--15078
		x"ff",	--15079
		x"ff",	--15080
		x"ff",	--15081
		x"ff",	--15082
		x"ff",	--15083
		x"ff",	--15084
		x"ff",	--15085
		x"ff",	--15086
		x"ff",	--15087
		x"ff",	--15088
		x"ff",	--15089
		x"ff",	--15090
		x"ff",	--15091
		x"ff",	--15092
		x"ff",	--15093
		x"ff",	--15094
		x"ff",	--15095
		x"ff",	--15096
		x"ff",	--15097
		x"ff",	--15098
		x"ff",	--15099
		x"ff",	--15100
		x"ff",	--15101
		x"ff",	--15102
		x"ff",	--15103
		x"ff",	--15104
		x"ff",	--15105
		x"ff",	--15106
		x"ff",	--15107
		x"ff",	--15108
		x"ff",	--15109
		x"ff",	--15110
		x"ff",	--15111
		x"ff",	--15112
		x"ff",	--15113
		x"ff",	--15114
		x"ff",	--15115
		x"ff",	--15116
		x"ff",	--15117
		x"ff",	--15118
		x"ff",	--15119
		x"ff",	--15120
		x"ff",	--15121
		x"ff",	--15122
		x"ff",	--15123
		x"ff",	--15124
		x"ff",	--15125
		x"ff",	--15126
		x"ff",	--15127
		x"ff",	--15128
		x"ff",	--15129
		x"ff",	--15130
		x"ff",	--15131
		x"ff",	--15132
		x"ff",	--15133
		x"ff",	--15134
		x"ff",	--15135
		x"ff",	--15136
		x"ff",	--15137
		x"ff",	--15138
		x"ff",	--15139
		x"ff",	--15140
		x"ff",	--15141
		x"ff",	--15142
		x"ff",	--15143
		x"ff",	--15144
		x"ff",	--15145
		x"ff",	--15146
		x"ff",	--15147
		x"ff",	--15148
		x"ff",	--15149
		x"ff",	--15150
		x"ff",	--15151
		x"ff",	--15152
		x"ff",	--15153
		x"ff",	--15154
		x"ff",	--15155
		x"ff",	--15156
		x"ff",	--15157
		x"ff",	--15158
		x"ff",	--15159
		x"ff",	--15160
		x"ff",	--15161
		x"ff",	--15162
		x"ff",	--15163
		x"ff",	--15164
		x"ff",	--15165
		x"ff",	--15166
		x"ff",	--15167
		x"ff",	--15168
		x"ff",	--15169
		x"ff",	--15170
		x"ff",	--15171
		x"ff",	--15172
		x"ff",	--15173
		x"ff",	--15174
		x"ff",	--15175
		x"ff",	--15176
		x"ff",	--15177
		x"ff",	--15178
		x"ff",	--15179
		x"ff",	--15180
		x"ff",	--15181
		x"ff",	--15182
		x"ff",	--15183
		x"ff",	--15184
		x"ff",	--15185
		x"ff",	--15186
		x"ff",	--15187
		x"ff",	--15188
		x"ff",	--15189
		x"ff",	--15190
		x"ff",	--15191
		x"ff",	--15192
		x"ff",	--15193
		x"ff",	--15194
		x"ff",	--15195
		x"ff",	--15196
		x"ff",	--15197
		x"ff",	--15198
		x"ff",	--15199
		x"ff",	--15200
		x"ff",	--15201
		x"ff",	--15202
		x"ff",	--15203
		x"ff",	--15204
		x"ff",	--15205
		x"ff",	--15206
		x"ff",	--15207
		x"ff",	--15208
		x"ff",	--15209
		x"ff",	--15210
		x"ff",	--15211
		x"ff",	--15212
		x"ff",	--15213
		x"ff",	--15214
		x"ff",	--15215
		x"ff",	--15216
		x"ff",	--15217
		x"ff",	--15218
		x"ff",	--15219
		x"ff",	--15220
		x"ff",	--15221
		x"ff",	--15222
		x"ff",	--15223
		x"ff",	--15224
		x"ff",	--15225
		x"ff",	--15226
		x"ff",	--15227
		x"ff",	--15228
		x"ff",	--15229
		x"ff",	--15230
		x"ff",	--15231
		x"ff",	--15232
		x"ff",	--15233
		x"ff",	--15234
		x"ff",	--15235
		x"ff",	--15236
		x"ff",	--15237
		x"ff",	--15238
		x"ff",	--15239
		x"ff",	--15240
		x"ff",	--15241
		x"ff",	--15242
		x"ff",	--15243
		x"ff",	--15244
		x"ff",	--15245
		x"ff",	--15246
		x"ff",	--15247
		x"ff",	--15248
		x"ff",	--15249
		x"ff",	--15250
		x"ff",	--15251
		x"ff",	--15252
		x"ff",	--15253
		x"ff",	--15254
		x"ff",	--15255
		x"ff",	--15256
		x"ff",	--15257
		x"ff",	--15258
		x"ff",	--15259
		x"ff",	--15260
		x"ff",	--15261
		x"ff",	--15262
		x"ff",	--15263
		x"ff",	--15264
		x"ff",	--15265
		x"ff",	--15266
		x"ff",	--15267
		x"ff",	--15268
		x"ff",	--15269
		x"ff",	--15270
		x"ff",	--15271
		x"ff",	--15272
		x"ff",	--15273
		x"ff",	--15274
		x"ff",	--15275
		x"ff",	--15276
		x"ff",	--15277
		x"ff",	--15278
		x"ff",	--15279
		x"ff",	--15280
		x"ff",	--15281
		x"ff",	--15282
		x"ff",	--15283
		x"ff",	--15284
		x"ff",	--15285
		x"ff",	--15286
		x"ff",	--15287
		x"ff",	--15288
		x"ff",	--15289
		x"ff",	--15290
		x"ff",	--15291
		x"ff",	--15292
		x"ff",	--15293
		x"ff",	--15294
		x"ff",	--15295
		x"ff",	--15296
		x"ff",	--15297
		x"ff",	--15298
		x"ff",	--15299
		x"ff",	--15300
		x"ff",	--15301
		x"ff",	--15302
		x"ff",	--15303
		x"ff",	--15304
		x"ff",	--15305
		x"ff",	--15306
		x"ff",	--15307
		x"ff",	--15308
		x"ff",	--15309
		x"ff",	--15310
		x"ff",	--15311
		x"ff",	--15312
		x"ff",	--15313
		x"ff",	--15314
		x"ff",	--15315
		x"ff",	--15316
		x"ff",	--15317
		x"ff",	--15318
		x"ff",	--15319
		x"ff",	--15320
		x"ff",	--15321
		x"ff",	--15322
		x"ff",	--15323
		x"ff",	--15324
		x"ff",	--15325
		x"ff",	--15326
		x"ff",	--15327
		x"ff",	--15328
		x"ff",	--15329
		x"ff",	--15330
		x"ff",	--15331
		x"ff",	--15332
		x"ff",	--15333
		x"ff",	--15334
		x"ff",	--15335
		x"ff",	--15336
		x"ff",	--15337
		x"ff",	--15338
		x"ff",	--15339
		x"ff",	--15340
		x"ff",	--15341
		x"ff",	--15342
		x"ff",	--15343
		x"ff",	--15344
		x"ff",	--15345
		x"ff",	--15346
		x"ff",	--15347
		x"ff",	--15348
		x"ff",	--15349
		x"ff",	--15350
		x"ff",	--15351
		x"ff",	--15352
		x"ff",	--15353
		x"ff",	--15354
		x"ff",	--15355
		x"ff",	--15356
		x"ff",	--15357
		x"ff",	--15358
		x"ff",	--15359
		x"ff",	--15360
		x"ff",	--15361
		x"ff",	--15362
		x"ff",	--15363
		x"ff",	--15364
		x"ff",	--15365
		x"ff",	--15366
		x"ff",	--15367
		x"ff",	--15368
		x"ff",	--15369
		x"ff",	--15370
		x"ff",	--15371
		x"ff",	--15372
		x"ff",	--15373
		x"ff",	--15374
		x"ff",	--15375
		x"ff",	--15376
		x"ff",	--15377
		x"ff",	--15378
		x"ff",	--15379
		x"ff",	--15380
		x"ff",	--15381
		x"ff",	--15382
		x"ff",	--15383
		x"ff",	--15384
		x"ff",	--15385
		x"ff",	--15386
		x"ff",	--15387
		x"ff",	--15388
		x"ff",	--15389
		x"ff",	--15390
		x"ff",	--15391
		x"ff",	--15392
		x"ff",	--15393
		x"ff",	--15394
		x"ff",	--15395
		x"ff",	--15396
		x"ff",	--15397
		x"ff",	--15398
		x"ff",	--15399
		x"ff",	--15400
		x"ff",	--15401
		x"ff",	--15402
		x"ff",	--15403
		x"ff",	--15404
		x"ff",	--15405
		x"ff",	--15406
		x"ff",	--15407
		x"ff",	--15408
		x"ff",	--15409
		x"ff",	--15410
		x"ff",	--15411
		x"ff",	--15412
		x"ff",	--15413
		x"ff",	--15414
		x"ff",	--15415
		x"ff",	--15416
		x"ff",	--15417
		x"ff",	--15418
		x"ff",	--15419
		x"ff",	--15420
		x"ff",	--15421
		x"ff",	--15422
		x"ff",	--15423
		x"ff",	--15424
		x"ff",	--15425
		x"ff",	--15426
		x"ff",	--15427
		x"ff",	--15428
		x"ff",	--15429
		x"ff",	--15430
		x"ff",	--15431
		x"ff",	--15432
		x"ff",	--15433
		x"ff",	--15434
		x"ff",	--15435
		x"ff",	--15436
		x"ff",	--15437
		x"ff",	--15438
		x"ff",	--15439
		x"ff",	--15440
		x"ff",	--15441
		x"ff",	--15442
		x"ff",	--15443
		x"ff",	--15444
		x"ff",	--15445
		x"ff",	--15446
		x"ff",	--15447
		x"ff",	--15448
		x"ff",	--15449
		x"ff",	--15450
		x"ff",	--15451
		x"ff",	--15452
		x"ff",	--15453
		x"ff",	--15454
		x"ff",	--15455
		x"ff",	--15456
		x"ff",	--15457
		x"ff",	--15458
		x"ff",	--15459
		x"ff",	--15460
		x"ff",	--15461
		x"ff",	--15462
		x"ff",	--15463
		x"ff",	--15464
		x"ff",	--15465
		x"ff",	--15466
		x"ff",	--15467
		x"ff",	--15468
		x"ff",	--15469
		x"ff",	--15470
		x"ff",	--15471
		x"ff",	--15472
		x"ff",	--15473
		x"ff",	--15474
		x"ff",	--15475
		x"ff",	--15476
		x"ff",	--15477
		x"ff",	--15478
		x"ff",	--15479
		x"ff",	--15480
		x"ff",	--15481
		x"ff",	--15482
		x"ff",	--15483
		x"ff",	--15484
		x"ff",	--15485
		x"ff",	--15486
		x"ff",	--15487
		x"ff",	--15488
		x"ff",	--15489
		x"ff",	--15490
		x"ff",	--15491
		x"ff",	--15492
		x"ff",	--15493
		x"ff",	--15494
		x"ff",	--15495
		x"ff",	--15496
		x"ff",	--15497
		x"ff",	--15498
		x"ff",	--15499
		x"ff",	--15500
		x"ff",	--15501
		x"ff",	--15502
		x"ff",	--15503
		x"ff",	--15504
		x"ff",	--15505
		x"ff",	--15506
		x"ff",	--15507
		x"ff",	--15508
		x"ff",	--15509
		x"ff",	--15510
		x"ff",	--15511
		x"ff",	--15512
		x"ff",	--15513
		x"ff",	--15514
		x"ff",	--15515
		x"ff",	--15516
		x"ff",	--15517
		x"ff",	--15518
		x"ff",	--15519
		x"ff",	--15520
		x"ff",	--15521
		x"ff",	--15522
		x"ff",	--15523
		x"ff",	--15524
		x"ff",	--15525
		x"ff",	--15526
		x"ff",	--15527
		x"ff",	--15528
		x"ff",	--15529
		x"ff",	--15530
		x"ff",	--15531
		x"ff",	--15532
		x"ff",	--15533
		x"ff",	--15534
		x"ff",	--15535
		x"ff",	--15536
		x"ff",	--15537
		x"ff",	--15538
		x"ff",	--15539
		x"ff",	--15540
		x"ff",	--15541
		x"ff",	--15542
		x"ff",	--15543
		x"ff",	--15544
		x"ff",	--15545
		x"ff",	--15546
		x"ff",	--15547
		x"ff",	--15548
		x"ff",	--15549
		x"ff",	--15550
		x"ff",	--15551
		x"ff",	--15552
		x"ff",	--15553
		x"ff",	--15554
		x"ff",	--15555
		x"ff",	--15556
		x"ff",	--15557
		x"ff",	--15558
		x"ff",	--15559
		x"ff",	--15560
		x"ff",	--15561
		x"ff",	--15562
		x"ff",	--15563
		x"ff",	--15564
		x"ff",	--15565
		x"ff",	--15566
		x"ff",	--15567
		x"ff",	--15568
		x"ff",	--15569
		x"ff",	--15570
		x"ff",	--15571
		x"ff",	--15572
		x"ff",	--15573
		x"ff",	--15574
		x"ff",	--15575
		x"ff",	--15576
		x"ff",	--15577
		x"ff",	--15578
		x"ff",	--15579
		x"ff",	--15580
		x"ff",	--15581
		x"ff",	--15582
		x"ff",	--15583
		x"ff",	--15584
		x"ff",	--15585
		x"ff",	--15586
		x"ff",	--15587
		x"ff",	--15588
		x"ff",	--15589
		x"ff",	--15590
		x"ff",	--15591
		x"ff",	--15592
		x"ff",	--15593
		x"ff",	--15594
		x"ff",	--15595
		x"ff",	--15596
		x"ff",	--15597
		x"ff",	--15598
		x"ff",	--15599
		x"ff",	--15600
		x"ff",	--15601
		x"ff",	--15602
		x"ff",	--15603
		x"ff",	--15604
		x"ff",	--15605
		x"ff",	--15606
		x"ff",	--15607
		x"ff",	--15608
		x"ff",	--15609
		x"ff",	--15610
		x"ff",	--15611
		x"ff",	--15612
		x"ff",	--15613
		x"ff",	--15614
		x"ff",	--15615
		x"ff",	--15616
		x"ff",	--15617
		x"ff",	--15618
		x"ff",	--15619
		x"ff",	--15620
		x"ff",	--15621
		x"ff",	--15622
		x"ff",	--15623
		x"ff",	--15624
		x"ff",	--15625
		x"ff",	--15626
		x"ff",	--15627
		x"ff",	--15628
		x"ff",	--15629
		x"ff",	--15630
		x"ff",	--15631
		x"ff",	--15632
		x"ff",	--15633
		x"ff",	--15634
		x"ff",	--15635
		x"ff",	--15636
		x"ff",	--15637
		x"ff",	--15638
		x"ff",	--15639
		x"ff",	--15640
		x"ff",	--15641
		x"ff",	--15642
		x"ff",	--15643
		x"ff",	--15644
		x"ff",	--15645
		x"ff",	--15646
		x"ff",	--15647
		x"ff",	--15648
		x"ff",	--15649
		x"ff",	--15650
		x"ff",	--15651
		x"ff",	--15652
		x"ff",	--15653
		x"ff",	--15654
		x"ff",	--15655
		x"ff",	--15656
		x"ff",	--15657
		x"ff",	--15658
		x"ff",	--15659
		x"ff",	--15660
		x"ff",	--15661
		x"ff",	--15662
		x"ff",	--15663
		x"ff",	--15664
		x"ff",	--15665
		x"ff",	--15666
		x"ff",	--15667
		x"ff",	--15668
		x"ff",	--15669
		x"ff",	--15670
		x"ff",	--15671
		x"ff",	--15672
		x"ff",	--15673
		x"ff",	--15674
		x"ff",	--15675
		x"ff",	--15676
		x"ff",	--15677
		x"ff",	--15678
		x"ff",	--15679
		x"ff",	--15680
		x"ff",	--15681
		x"ff",	--15682
		x"ff",	--15683
		x"ff",	--15684
		x"ff",	--15685
		x"ff",	--15686
		x"ff",	--15687
		x"ff",	--15688
		x"ff",	--15689
		x"ff",	--15690
		x"ff",	--15691
		x"ff",	--15692
		x"ff",	--15693
		x"ff",	--15694
		x"ff",	--15695
		x"ff",	--15696
		x"ff",	--15697
		x"ff",	--15698
		x"ff",	--15699
		x"ff",	--15700
		x"ff",	--15701
		x"ff",	--15702
		x"ff",	--15703
		x"ff",	--15704
		x"ff",	--15705
		x"ff",	--15706
		x"ff",	--15707
		x"ff",	--15708
		x"ff",	--15709
		x"ff",	--15710
		x"ff",	--15711
		x"ff",	--15712
		x"ff",	--15713
		x"ff",	--15714
		x"ff",	--15715
		x"ff",	--15716
		x"ff",	--15717
		x"ff",	--15718
		x"ff",	--15719
		x"ff",	--15720
		x"ff",	--15721
		x"ff",	--15722
		x"ff",	--15723
		x"ff",	--15724
		x"ff",	--15725
		x"ff",	--15726
		x"ff",	--15727
		x"ff",	--15728
		x"ff",	--15729
		x"ff",	--15730
		x"ff",	--15731
		x"ff",	--15732
		x"ff",	--15733
		x"ff",	--15734
		x"ff",	--15735
		x"ff",	--15736
		x"ff",	--15737
		x"ff",	--15738
		x"ff",	--15739
		x"ff",	--15740
		x"ff",	--15741
		x"ff",	--15742
		x"ff",	--15743
		x"ff",	--15744
		x"ff",	--15745
		x"ff",	--15746
		x"ff",	--15747
		x"ff",	--15748
		x"ff",	--15749
		x"ff",	--15750
		x"ff",	--15751
		x"ff",	--15752
		x"ff",	--15753
		x"ff",	--15754
		x"ff",	--15755
		x"ff",	--15756
		x"ff",	--15757
		x"ff",	--15758
		x"ff",	--15759
		x"ff",	--15760
		x"ff",	--15761
		x"ff",	--15762
		x"ff",	--15763
		x"ff",	--15764
		x"ff",	--15765
		x"ff",	--15766
		x"ff",	--15767
		x"ff",	--15768
		x"ff",	--15769
		x"ff",	--15770
		x"ff",	--15771
		x"ff",	--15772
		x"ff",	--15773
		x"ff",	--15774
		x"ff",	--15775
		x"ff",	--15776
		x"ff",	--15777
		x"ff",	--15778
		x"ff",	--15779
		x"ff",	--15780
		x"ff",	--15781
		x"ff",	--15782
		x"ff",	--15783
		x"ff",	--15784
		x"ff",	--15785
		x"ff",	--15786
		x"ff",	--15787
		x"ff",	--15788
		x"ff",	--15789
		x"ff",	--15790
		x"ff",	--15791
		x"ff",	--15792
		x"ff",	--15793
		x"ff",	--15794
		x"ff",	--15795
		x"ff",	--15796
		x"ff",	--15797
		x"ff",	--15798
		x"ff",	--15799
		x"ff",	--15800
		x"ff",	--15801
		x"ff",	--15802
		x"ff",	--15803
		x"ff",	--15804
		x"ff",	--15805
		x"ff",	--15806
		x"ff",	--15807
		x"ff",	--15808
		x"ff",	--15809
		x"ff",	--15810
		x"ff",	--15811
		x"ff",	--15812
		x"ff",	--15813
		x"ff",	--15814
		x"ff",	--15815
		x"ff",	--15816
		x"ff",	--15817
		x"ff",	--15818
		x"ff",	--15819
		x"ff",	--15820
		x"ff",	--15821
		x"ff",	--15822
		x"ff",	--15823
		x"ff",	--15824
		x"ff",	--15825
		x"ff",	--15826
		x"ff",	--15827
		x"ff",	--15828
		x"ff",	--15829
		x"ff",	--15830
		x"ff",	--15831
		x"ff",	--15832
		x"ff",	--15833
		x"ff",	--15834
		x"ff",	--15835
		x"ff",	--15836
		x"ff",	--15837
		x"ff",	--15838
		x"ff",	--15839
		x"ff",	--15840
		x"ff",	--15841
		x"ff",	--15842
		x"ff",	--15843
		x"ff",	--15844
		x"ff",	--15845
		x"ff",	--15846
		x"ff",	--15847
		x"ff",	--15848
		x"ff",	--15849
		x"ff",	--15850
		x"ff",	--15851
		x"ff",	--15852
		x"ff",	--15853
		x"ff",	--15854
		x"ff",	--15855
		x"ff",	--15856
		x"ff",	--15857
		x"ff",	--15858
		x"ff",	--15859
		x"ff",	--15860
		x"ff",	--15861
		x"ff",	--15862
		x"ff",	--15863
		x"ff",	--15864
		x"ff",	--15865
		x"ff",	--15866
		x"ff",	--15867
		x"ff",	--15868
		x"ff",	--15869
		x"ff",	--15870
		x"ff",	--15871
		x"ff",	--15872
		x"ff",	--15873
		x"ff",	--15874
		x"ff",	--15875
		x"ff",	--15876
		x"ff",	--15877
		x"ff",	--15878
		x"ff",	--15879
		x"ff",	--15880
		x"ff",	--15881
		x"ff",	--15882
		x"ff",	--15883
		x"ff",	--15884
		x"ff",	--15885
		x"ff",	--15886
		x"ff",	--15887
		x"ff",	--15888
		x"ff",	--15889
		x"ff",	--15890
		x"ff",	--15891
		x"ff",	--15892
		x"ff",	--15893
		x"ff",	--15894
		x"ff",	--15895
		x"ff",	--15896
		x"ff",	--15897
		x"ff",	--15898
		x"ff",	--15899
		x"ff",	--15900
		x"ff",	--15901
		x"ff",	--15902
		x"ff",	--15903
		x"ff",	--15904
		x"ff",	--15905
		x"ff",	--15906
		x"ff",	--15907
		x"ff",	--15908
		x"ff",	--15909
		x"ff",	--15910
		x"ff",	--15911
		x"ff",	--15912
		x"ff",	--15913
		x"ff",	--15914
		x"ff",	--15915
		x"ff",	--15916
		x"ff",	--15917
		x"ff",	--15918
		x"ff",	--15919
		x"ff",	--15920
		x"ff",	--15921
		x"ff",	--15922
		x"ff",	--15923
		x"ff",	--15924
		x"ff",	--15925
		x"ff",	--15926
		x"ff",	--15927
		x"ff",	--15928
		x"ff",	--15929
		x"ff",	--15930
		x"ff",	--15931
		x"ff",	--15932
		x"ff",	--15933
		x"ff",	--15934
		x"ff",	--15935
		x"ff",	--15936
		x"ff",	--15937
		x"ff",	--15938
		x"ff",	--15939
		x"ff",	--15940
		x"ff",	--15941
		x"ff",	--15942
		x"ff",	--15943
		x"ff",	--15944
		x"ff",	--15945
		x"ff",	--15946
		x"ff",	--15947
		x"ff",	--15948
		x"ff",	--15949
		x"ff",	--15950
		x"ff",	--15951
		x"ff",	--15952
		x"ff",	--15953
		x"ff",	--15954
		x"ff",	--15955
		x"ff",	--15956
		x"ff",	--15957
		x"ff",	--15958
		x"ff",	--15959
		x"ff",	--15960
		x"ff",	--15961
		x"ff",	--15962
		x"ff",	--15963
		x"ff",	--15964
		x"ff",	--15965
		x"ff",	--15966
		x"ff",	--15967
		x"ff",	--15968
		x"ff",	--15969
		x"ff",	--15970
		x"ff",	--15971
		x"ff",	--15972
		x"ff",	--15973
		x"ff",	--15974
		x"ff",	--15975
		x"ff",	--15976
		x"ff",	--15977
		x"ff",	--15978
		x"ff",	--15979
		x"ff",	--15980
		x"ff",	--15981
		x"ff",	--15982
		x"ff",	--15983
		x"ff",	--15984
		x"ff",	--15985
		x"ff",	--15986
		x"ff",	--15987
		x"ff",	--15988
		x"ff",	--15989
		x"ff",	--15990
		x"ff",	--15991
		x"ff",	--15992
		x"ff",	--15993
		x"ff",	--15994
		x"ff",	--15995
		x"ff",	--15996
		x"ff",	--15997
		x"ff",	--15998
		x"ff",	--15999
		x"ff",	--16000
		x"ff",	--16001
		x"ff",	--16002
		x"ff",	--16003
		x"ff",	--16004
		x"ff",	--16005
		x"ff",	--16006
		x"ff",	--16007
		x"ff",	--16008
		x"ff",	--16009
		x"ff",	--16010
		x"ff",	--16011
		x"ff",	--16012
		x"ff",	--16013
		x"ff",	--16014
		x"ff",	--16015
		x"ff",	--16016
		x"ff",	--16017
		x"ff",	--16018
		x"ff",	--16019
		x"ff",	--16020
		x"ff",	--16021
		x"ff",	--16022
		x"ff",	--16023
		x"ff",	--16024
		x"ff",	--16025
		x"ff",	--16026
		x"ff",	--16027
		x"ff",	--16028
		x"ff",	--16029
		x"ff",	--16030
		x"ff",	--16031
		x"ff",	--16032
		x"ff",	--16033
		x"ff",	--16034
		x"ff",	--16035
		x"ff",	--16036
		x"ff",	--16037
		x"ff",	--16038
		x"ff",	--16039
		x"ff",	--16040
		x"ff",	--16041
		x"ff",	--16042
		x"ff",	--16043
		x"ff",	--16044
		x"ff",	--16045
		x"ff",	--16046
		x"ff",	--16047
		x"ff",	--16048
		x"ff",	--16049
		x"ff",	--16050
		x"ff",	--16051
		x"ff",	--16052
		x"ff",	--16053
		x"ff",	--16054
		x"ff",	--16055
		x"ff",	--16056
		x"ff",	--16057
		x"ff",	--16058
		x"ff",	--16059
		x"ff",	--16060
		x"ff",	--16061
		x"ff",	--16062
		x"ff",	--16063
		x"ff",	--16064
		x"ff",	--16065
		x"ff",	--16066
		x"ff",	--16067
		x"ff",	--16068
		x"ff",	--16069
		x"ff",	--16070
		x"ff",	--16071
		x"ff",	--16072
		x"ff",	--16073
		x"ff",	--16074
		x"ff",	--16075
		x"ff",	--16076
		x"ff",	--16077
		x"ff",	--16078
		x"ff",	--16079
		x"ff",	--16080
		x"ff",	--16081
		x"ff",	--16082
		x"ff",	--16083
		x"ff",	--16084
		x"ff",	--16085
		x"ff",	--16086
		x"ff",	--16087
		x"ff",	--16088
		x"ff",	--16089
		x"ff",	--16090
		x"ff",	--16091
		x"ff",	--16092
		x"ff",	--16093
		x"ff",	--16094
		x"ff",	--16095
		x"ff",	--16096
		x"ff",	--16097
		x"ff",	--16098
		x"ff",	--16099
		x"ff",	--16100
		x"ff",	--16101
		x"ff",	--16102
		x"ff",	--16103
		x"ff",	--16104
		x"ff",	--16105
		x"ff",	--16106
		x"ff",	--16107
		x"ff",	--16108
		x"ff",	--16109
		x"ff",	--16110
		x"ff",	--16111
		x"ff",	--16112
		x"ff",	--16113
		x"ff",	--16114
		x"ff",	--16115
		x"ff",	--16116
		x"ff",	--16117
		x"ff",	--16118
		x"ff",	--16119
		x"ff",	--16120
		x"ff",	--16121
		x"ff",	--16122
		x"ff",	--16123
		x"ff",	--16124
		x"ff",	--16125
		x"ff",	--16126
		x"ff",	--16127
		x"ff",	--16128
		x"ff",	--16129
		x"ff",	--16130
		x"ff",	--16131
		x"ff",	--16132
		x"ff",	--16133
		x"ff",	--16134
		x"ff",	--16135
		x"ff",	--16136
		x"ff",	--16137
		x"ff",	--16138
		x"ff",	--16139
		x"ff",	--16140
		x"ff",	--16141
		x"ff",	--16142
		x"ff",	--16143
		x"ff",	--16144
		x"ff",	--16145
		x"ff",	--16146
		x"ff",	--16147
		x"ff",	--16148
		x"ff",	--16149
		x"ff",	--16150
		x"ff",	--16151
		x"ff",	--16152
		x"ff",	--16153
		x"ff",	--16154
		x"ff",	--16155
		x"ff",	--16156
		x"ff",	--16157
		x"ff",	--16158
		x"ff",	--16159
		x"ff",	--16160
		x"ff",	--16161
		x"ff",	--16162
		x"ff",	--16163
		x"ff",	--16164
		x"ff",	--16165
		x"ff",	--16166
		x"ff",	--16167
		x"ff",	--16168
		x"ff",	--16169
		x"ff",	--16170
		x"ff",	--16171
		x"ff",	--16172
		x"ff",	--16173
		x"ff",	--16174
		x"ff",	--16175
		x"ff",	--16176
		x"ff",	--16177
		x"ff",	--16178
		x"ff",	--16179
		x"ff",	--16180
		x"ff",	--16181
		x"ff",	--16182
		x"ff",	--16183
		x"ff",	--16184
		x"ff",	--16185
		x"ff",	--16186
		x"ff",	--16187
		x"ff",	--16188
		x"ff",	--16189
		x"ff",	--16190
		x"ff",	--16191
		x"ff",	--16192
		x"ff",	--16193
		x"ff",	--16194
		x"ff",	--16195
		x"ff",	--16196
		x"ff",	--16197
		x"ff",	--16198
		x"ff",	--16199
		x"ff",	--16200
		x"ff",	--16201
		x"ff",	--16202
		x"ff",	--16203
		x"ff",	--16204
		x"ff",	--16205
		x"ff",	--16206
		x"ff",	--16207
		x"ff",	--16208
		x"ff",	--16209
		x"ff",	--16210
		x"ff",	--16211
		x"ff",	--16212
		x"ff",	--16213
		x"ff",	--16214
		x"ff",	--16215
		x"ff",	--16216
		x"ff",	--16217
		x"ff",	--16218
		x"ff",	--16219
		x"ff",	--16220
		x"ff",	--16221
		x"ff",	--16222
		x"ff",	--16223
		x"ff",	--16224
		x"ff",	--16225
		x"ff",	--16226
		x"ff",	--16227
		x"ff",	--16228
		x"ff",	--16229
		x"ff",	--16230
		x"ff",	--16231
		x"ff",	--16232
		x"ff",	--16233
		x"ff",	--16234
		x"ff",	--16235
		x"ff",	--16236
		x"ff",	--16237
		x"ff",	--16238
		x"ff",	--16239
		x"ff",	--16240
		x"ff",	--16241
		x"ff",	--16242
		x"ff",	--16243
		x"ff",	--16244
		x"ff",	--16245
		x"ff",	--16246
		x"ff",	--16247
		x"ff",	--16248
		x"ff",	--16249
		x"ff",	--16250
		x"ff",	--16251
		x"ff",	--16252
		x"ff",	--16253
		x"ff",	--16254
		x"ff",	--16255
		x"ff",	--16256
		x"ff",	--16257
		x"ff",	--16258
		x"ff",	--16259
		x"ff",	--16260
		x"ff",	--16261
		x"ff",	--16262
		x"ff",	--16263
		x"ff",	--16264
		x"ff",	--16265
		x"ff",	--16266
		x"ff",	--16267
		x"ff",	--16268
		x"ff",	--16269
		x"ff",	--16270
		x"ff",	--16271
		x"ff",	--16272
		x"ff",	--16273
		x"ff",	--16274
		x"ff",	--16275
		x"ff",	--16276
		x"ff",	--16277
		x"ff",	--16278
		x"ff",	--16279
		x"ff",	--16280
		x"ff",	--16281
		x"ff",	--16282
		x"ff",	--16283
		x"ff",	--16284
		x"ff",	--16285
		x"ff",	--16286
		x"ff",	--16287
		x"ff",	--16288
		x"ff",	--16289
		x"ff",	--16290
		x"ff",	--16291
		x"ff",	--16292
		x"ff",	--16293
		x"ff",	--16294
		x"ff",	--16295
		x"ff",	--16296
		x"ff",	--16297
		x"ff",	--16298
		x"ff",	--16299
		x"ff",	--16300
		x"ff",	--16301
		x"ff",	--16302
		x"ff",	--16303
		x"ff",	--16304
		x"ff",	--16305
		x"ff",	--16306
		x"ff",	--16307
		x"ff",	--16308
		x"ff",	--16309
		x"ff",	--16310
		x"ff",	--16311
		x"ff",	--16312
		x"ff",	--16313
		x"ff",	--16314
		x"ff",	--16315
		x"ff",	--16316
		x"ff",	--16317
		x"ff",	--16318
		x"ff",	--16319
		x"ff",	--16320
		x"ff",	--16321
		x"ff",	--16322
		x"ff",	--16323
		x"ff",	--16324
		x"ff",	--16325
		x"ff",	--16326
		x"ff",	--16327
		x"ff",	--16328
		x"ff",	--16329
		x"ff",	--16330
		x"ff",	--16331
		x"ff",	--16332
		x"ff",	--16333
		x"ff",	--16334
		x"ff",	--16335
		x"ff",	--16336
		x"ff",	--16337
		x"ff",	--16338
		x"ff",	--16339
		x"ff",	--16340
		x"ff",	--16341
		x"ff",	--16342
		x"ff",	--16343
		x"ff",	--16344
		x"ff",	--16345
		x"ff",	--16346
		x"ff",	--16347
		x"ff",	--16348
		x"ff",	--16349
		x"ff",	--16350
		x"ff",	--16351
		x"ff",	--16352
		x"ff",	--16353
		x"ff",	--16354
		x"ff",	--16355
		x"ff",	--16356
		x"ff",	--16357
		x"ff",	--16358
		x"ff",	--16359
		x"ff",	--16360
		x"ff",	--16361
		x"ff",	--16362
		x"ff",	--16363
		x"ff",	--16364
		x"ff",	--16365
		x"ff",	--16366
		x"ff",	--16367
		x"83",	--16368
		x"83",	--16369
		x"83",	--16370
		x"83",	--16371
		x"83",	--16372
		x"83",	--16373
		x"83",	--16374
		x"9c",	--16375
		x"98",	--16376
		x"83",	--16377
		x"83",	--16378
		x"83",	--16379
		x"83",	--16380
		x"83",	--16381
		x"83",	--16382
		x"80");	--16383

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
