library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"4a",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"00",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"4a",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"5e",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"4a",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"4a",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"00",	--29
		x"f9",	--30
		x"31",	--31
		x"c2",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"f2",	--38
		x"19",	--39
		x"c2",	--40
		x"22",	--41
		x"3e",	--42
		x"00",	--43
		x"1f",	--44
		x"b0",	--45
		x"3e",	--46
		x"b0",	--47
		x"a6",	--48
		x"c2",	--49
		x"19",	--50
		x"30",	--51
		x"92",	--52
		x"b0",	--53
		x"fc",	--54
		x"b1",	--55
		x"b9",	--56
		x"00",	--57
		x"b0",	--58
		x"fc",	--59
		x"21",	--60
		x"03",	--61
		x"30",	--62
		x"cf",	--63
		x"30",	--64
		x"d6",	--65
		x"b0",	--66
		x"fc",	--67
		x"31",	--68
		x"06",	--69
		x"30",	--70
		x"78",	--71
		x"30",	--72
		x"e2",	--73
		x"b0",	--74
		x"fc",	--75
		x"21",	--76
		x"3e",	--77
		x"7e",	--78
		x"7f",	--79
		x"77",	--80
		x"b0",	--81
		x"a8",	--82
		x"3e",	--83
		x"1e",	--84
		x"7f",	--85
		x"72",	--86
		x"b0",	--87
		x"a8",	--88
		x"3e",	--89
		x"cc",	--90
		x"7f",	--91
		x"70",	--92
		x"b0",	--93
		x"a8",	--94
		x"0c",	--95
		x"3d",	--96
		x"20",	--97
		x"3e",	--98
		x"80",	--99
		x"0f",	--100
		x"3f",	--101
		x"0a",	--102
		x"b0",	--103
		x"b6",	--104
		x"0f",	--105
		x"3f",	--106
		x"0a",	--107
		x"b0",	--108
		x"fe",	--109
		x"0c",	--110
		x"3d",	--111
		x"20",	--112
		x"3e",	--113
		x"88",	--114
		x"0f",	--115
		x"b0",	--116
		x"b6",	--117
		x"0f",	--118
		x"b0",	--119
		x"fe",	--120
		x"0e",	--121
		x"0f",	--122
		x"3f",	--123
		x"0a",	--124
		x"b0",	--125
		x"c2",	--126
		x"32",	--127
		x"0b",	--128
		x"30",	--129
		x"ee",	--130
		x"b0",	--131
		x"fc",	--132
		x"21",	--133
		x"0a",	--134
		x"32",	--135
		x"10",	--136
		x"1b",	--137
		x"3b",	--138
		x"09",	--139
		x"0a",	--140
		x"1f",	--141
		x"4e",	--142
		x"7e",	--143
		x"0f",	--144
		x"03",	--145
		x"0f",	--146
		x"7e",	--147
		x"fd",	--148
		x"4f",	--149
		x"02",	--150
		x"5f",	--151
		x"0b",	--152
		x"c2",	--153
		x"19",	--154
		x"b0",	--155
		x"4c",	--156
		x"0f",	--157
		x"e8",	--158
		x"b0",	--159
		x"74",	--160
		x"7f",	--161
		x"1c",	--162
		x"7f",	--163
		x"0d",	--164
		x"22",	--165
		x"30",	--166
		x"f1",	--167
		x"b0",	--168
		x"fc",	--169
		x"21",	--170
		x"3f",	--171
		x"14",	--172
		x"0f",	--173
		x"0a",	--174
		x"ca",	--175
		x"00",	--176
		x"0f",	--177
		x"30",	--178
		x"f4",	--179
		x"b0",	--180
		x"fc",	--181
		x"21",	--182
		x"0e",	--183
		x"3e",	--184
		x"14",	--185
		x"5f",	--186
		x"14",	--187
		x"b0",	--188
		x"d2",	--189
		x"c2",	--190
		x"0a",	--191
		x"c6",	--192
		x"3a",	--193
		x"30",	--194
		x"fa",	--195
		x"b0",	--196
		x"fc",	--197
		x"21",	--198
		x"bf",	--199
		x"3a",	--200
		x"28",	--201
		x"bc",	--202
		x"4e",	--203
		x"8e",	--204
		x"0e",	--205
		x"30",	--206
		x"fe",	--207
		x"81",	--208
		x"40",	--209
		x"b0",	--210
		x"fc",	--211
		x"21",	--212
		x"3e",	--213
		x"14",	--214
		x"0e",	--215
		x"0e",	--216
		x"1f",	--217
		x"3c",	--218
		x"ce",	--219
		x"00",	--220
		x"1a",	--221
		x"a8",	--222
		x"30",	--223
		x"48",	--224
		x"82",	--225
		x"08",	--226
		x"82",	--227
		x"06",	--228
		x"30",	--229
		x"31",	--230
		x"ff",	--231
		x"20",	--232
		x"01",	--233
		x"39",	--234
		x"cf",	--235
		x"02",	--236
		x"36",	--237
		x"0d",	--238
		x"0e",	--239
		x"2e",	--240
		x"0f",	--241
		x"2f",	--242
		x"b0",	--243
		x"9c",	--244
		x"81",	--245
		x"00",	--246
		x"40",	--247
		x"0d",	--248
		x"0e",	--249
		x"0f",	--250
		x"2f",	--251
		x"b0",	--252
		x"9c",	--253
		x"81",	--254
		x"00",	--255
		x"37",	--256
		x"1e",	--257
		x"04",	--258
		x"0f",	--259
		x"b0",	--260
		x"66",	--261
		x"0c",	--262
		x"3d",	--263
		x"c8",	--264
		x"b0",	--265
		x"36",	--266
		x"0d",	--267
		x"0e",	--268
		x"1f",	--269
		x"08",	--270
		x"b0",	--271
		x"52",	--272
		x"1e",	--273
		x"02",	--274
		x"0f",	--275
		x"b0",	--276
		x"66",	--277
		x"0c",	--278
		x"3d",	--279
		x"c8",	--280
		x"b0",	--281
		x"36",	--282
		x"0d",	--283
		x"0e",	--284
		x"1f",	--285
		x"06",	--286
		x"b0",	--287
		x"52",	--288
		x"0f",	--289
		x"31",	--290
		x"30",	--291
		x"30",	--292
		x"50",	--293
		x"81",	--294
		x"08",	--295
		x"b0",	--296
		x"fc",	--297
		x"1f",	--298
		x"08",	--299
		x"6f",	--300
		x"8f",	--301
		x"81",	--302
		x"00",	--303
		x"30",	--304
		x"61",	--305
		x"b0",	--306
		x"fc",	--307
		x"21",	--308
		x"3f",	--309
		x"31",	--310
		x"30",	--311
		x"30",	--312
		x"72",	--313
		x"b0",	--314
		x"fc",	--315
		x"21",	--316
		x"3f",	--317
		x"e3",	--318
		x"0b",	--319
		x"31",	--320
		x"fa",	--321
		x"0b",	--322
		x"30",	--323
		x"01",	--324
		x"b0",	--325
		x"fc",	--326
		x"21",	--327
		x"fb",	--328
		x"20",	--329
		x"01",	--330
		x"2a",	--331
		x"cb",	--332
		x"02",	--333
		x"27",	--334
		x"0d",	--335
		x"0e",	--336
		x"2e",	--337
		x"0f",	--338
		x"2f",	--339
		x"b0",	--340
		x"9c",	--341
		x"81",	--342
		x"00",	--343
		x"2f",	--344
		x"0d",	--345
		x"0e",	--346
		x"0f",	--347
		x"2f",	--348
		x"b0",	--349
		x"9c",	--350
		x"81",	--351
		x"00",	--352
		x"26",	--353
		x"11",	--354
		x"04",	--355
		x"11",	--356
		x"08",	--357
		x"30",	--358
		x"4f",	--359
		x"b0",	--360
		x"fc",	--361
		x"31",	--362
		x"06",	--363
		x"1f",	--364
		x"04",	--365
		x"9f",	--366
		x"02",	--367
		x"00",	--368
		x"0f",	--369
		x"31",	--370
		x"06",	--371
		x"3b",	--372
		x"30",	--373
		x"30",	--374
		x"09",	--375
		x"b0",	--376
		x"fc",	--377
		x"6f",	--378
		x"8f",	--379
		x"81",	--380
		x"00",	--381
		x"30",	--382
		x"1a",	--383
		x"b0",	--384
		x"fc",	--385
		x"21",	--386
		x"3f",	--387
		x"31",	--388
		x"06",	--389
		x"3b",	--390
		x"30",	--391
		x"30",	--392
		x"2f",	--393
		x"b0",	--394
		x"fc",	--395
		x"21",	--396
		x"3f",	--397
		x"e3",	--398
		x"0b",	--399
		x"21",	--400
		x"0b",	--401
		x"30",	--402
		x"5b",	--403
		x"b0",	--404
		x"fc",	--405
		x"21",	--406
		x"fb",	--407
		x"20",	--408
		x"01",	--409
		x"1b",	--410
		x"cb",	--411
		x"02",	--412
		x"18",	--413
		x"0d",	--414
		x"0e",	--415
		x"2e",	--416
		x"0f",	--417
		x"2f",	--418
		x"b0",	--419
		x"9c",	--420
		x"81",	--421
		x"00",	--422
		x"1f",	--423
		x"1f",	--424
		x"02",	--425
		x"2f",	--426
		x"0f",	--427
		x"30",	--428
		x"4f",	--429
		x"b0",	--430
		x"fc",	--431
		x"31",	--432
		x"06",	--433
		x"0f",	--434
		x"21",	--435
		x"3b",	--436
		x"30",	--437
		x"30",	--438
		x"09",	--439
		x"b0",	--440
		x"fc",	--441
		x"6f",	--442
		x"8f",	--443
		x"81",	--444
		x"00",	--445
		x"30",	--446
		x"62",	--447
		x"b0",	--448
		x"fc",	--449
		x"21",	--450
		x"3f",	--451
		x"21",	--452
		x"3b",	--453
		x"30",	--454
		x"30",	--455
		x"2f",	--456
		x"b0",	--457
		x"fc",	--458
		x"21",	--459
		x"3f",	--460
		x"e5",	--461
		x"0b",	--462
		x"0a",	--463
		x"09",	--464
		x"08",	--465
		x"07",	--466
		x"8f",	--467
		x"00",	--468
		x"8d",	--469
		x"00",	--470
		x"6c",	--471
		x"4c",	--472
		x"5f",	--473
		x"0b",	--474
		x"1b",	--475
		x"08",	--476
		x"0a",	--477
		x"07",	--478
		x"09",	--479
		x"18",	--480
		x"7a",	--481
		x"0a",	--482
		x"35",	--483
		x"2c",	--484
		x"0c",	--485
		x"0c",	--486
		x"0c",	--487
		x"0c",	--488
		x"8f",	--489
		x"00",	--490
		x"3c",	--491
		x"d0",	--492
		x"6a",	--493
		x"8a",	--494
		x"0c",	--495
		x"8f",	--496
		x"00",	--497
		x"17",	--498
		x"19",	--499
		x"0a",	--500
		x"08",	--501
		x"7c",	--502
		x"4c",	--503
		x"40",	--504
		x"7c",	--505
		x"78",	--506
		x"1b",	--507
		x"7c",	--508
		x"20",	--509
		x"43",	--510
		x"4a",	--511
		x"7a",	--512
		x"d0",	--513
		x"07",	--514
		x"dd",	--515
		x"7a",	--516
		x"0a",	--517
		x"46",	--518
		x"2a",	--519
		x"0a",	--520
		x"0c",	--521
		x"0c",	--522
		x"0c",	--523
		x"0c",	--524
		x"8f",	--525
		x"00",	--526
		x"3c",	--527
		x"d0",	--528
		x"68",	--529
		x"88",	--530
		x"0c",	--531
		x"8f",	--532
		x"00",	--533
		x"dc",	--534
		x"17",	--535
		x"da",	--536
		x"4a",	--537
		x"7a",	--538
		x"9f",	--539
		x"7a",	--540
		x"06",	--541
		x"0a",	--542
		x"2c",	--543
		x"0c",	--544
		x"0c",	--545
		x"0c",	--546
		x"0c",	--547
		x"8f",	--548
		x"00",	--549
		x"3c",	--550
		x"a9",	--551
		x"c4",	--552
		x"4a",	--553
		x"7a",	--554
		x"bf",	--555
		x"7a",	--556
		x"06",	--557
		x"1e",	--558
		x"2c",	--559
		x"0c",	--560
		x"0c",	--561
		x"0c",	--562
		x"0c",	--563
		x"8f",	--564
		x"00",	--565
		x"3c",	--566
		x"c9",	--567
		x"b4",	--568
		x"9d",	--569
		x"00",	--570
		x"0f",	--571
		x"37",	--572
		x"38",	--573
		x"39",	--574
		x"3a",	--575
		x"3b",	--576
		x"30",	--577
		x"9d",	--578
		x"00",	--579
		x"0f",	--580
		x"1f",	--581
		x"0f",	--582
		x"37",	--583
		x"38",	--584
		x"39",	--585
		x"3a",	--586
		x"3b",	--587
		x"30",	--588
		x"8c",	--589
		x"0c",	--590
		x"30",	--591
		x"71",	--592
		x"b0",	--593
		x"fc",	--594
		x"21",	--595
		x"0f",	--596
		x"37",	--597
		x"38",	--598
		x"39",	--599
		x"3a",	--600
		x"3b",	--601
		x"30",	--602
		x"0b",	--603
		x"0a",	--604
		x"0b",	--605
		x"0a",	--606
		x"8f",	--607
		x"00",	--608
		x"8f",	--609
		x"02",	--610
		x"8f",	--611
		x"04",	--612
		x"0c",	--613
		x"0d",	--614
		x"3e",	--615
		x"00",	--616
		x"3f",	--617
		x"6e",	--618
		x"b0",	--619
		x"9a",	--620
		x"8b",	--621
		x"02",	--622
		x"02",	--623
		x"32",	--624
		x"03",	--625
		x"82",	--626
		x"32",	--627
		x"b2",	--628
		x"18",	--629
		x"38",	--630
		x"9b",	--631
		x"3a",	--632
		x"06",	--633
		x"32",	--634
		x"0f",	--635
		x"3a",	--636
		x"3b",	--637
		x"30",	--638
		x"0b",	--639
		x"09",	--640
		x"08",	--641
		x"8f",	--642
		x"06",	--643
		x"bf",	--644
		x"00",	--645
		x"08",	--646
		x"2b",	--647
		x"1e",	--648
		x"02",	--649
		x"0f",	--650
		x"b0",	--651
		x"66",	--652
		x"0c",	--653
		x"3d",	--654
		x"00",	--655
		x"b0",	--656
		x"12",	--657
		x"08",	--658
		x"09",	--659
		x"1e",	--660
		x"06",	--661
		x"0f",	--662
		x"b0",	--663
		x"66",	--664
		x"0c",	--665
		x"0d",	--666
		x"0e",	--667
		x"0f",	--668
		x"b0",	--669
		x"c2",	--670
		x"b0",	--671
		x"a2",	--672
		x"8b",	--673
		x"04",	--674
		x"9b",	--675
		x"00",	--676
		x"38",	--677
		x"39",	--678
		x"3b",	--679
		x"30",	--680
		x"0b",	--681
		x"0a",	--682
		x"09",	--683
		x"0a",	--684
		x"0b",	--685
		x"8f",	--686
		x"06",	--687
		x"8f",	--688
		x"08",	--689
		x"29",	--690
		x"1e",	--691
		x"02",	--692
		x"0f",	--693
		x"b0",	--694
		x"66",	--695
		x"0c",	--696
		x"0d",	--697
		x"0e",	--698
		x"0f",	--699
		x"b0",	--700
		x"12",	--701
		x"0a",	--702
		x"0b",	--703
		x"1e",	--704
		x"06",	--705
		x"0f",	--706
		x"b0",	--707
		x"66",	--708
		x"0c",	--709
		x"0d",	--710
		x"0e",	--711
		x"0f",	--712
		x"b0",	--713
		x"c2",	--714
		x"b0",	--715
		x"a2",	--716
		x"89",	--717
		x"04",	--718
		x"39",	--719
		x"3a",	--720
		x"3b",	--721
		x"30",	--722
		x"30",	--723
		x"1c",	--724
		x"00",	--725
		x"3c",	--726
		x"40",	--727
		x"0e",	--728
		x"0d",	--729
		x"0d",	--730
		x"0d",	--731
		x"3d",	--732
		x"0a",	--733
		x"cd",	--734
		x"00",	--735
		x"8d",	--736
		x"02",	--737
		x"1c",	--738
		x"82",	--739
		x"00",	--740
		x"0f",	--741
		x"30",	--742
		x"3f",	--743
		x"30",	--744
		x"0b",	--745
		x"1b",	--746
		x"00",	--747
		x"1b",	--748
		x"0e",	--749
		x"5f",	--750
		x"0a",	--751
		x"13",	--752
		x"3d",	--753
		x"0e",	--754
		x"0c",	--755
		x"04",	--756
		x"2d",	--757
		x"cd",	--758
		x"fc",	--759
		x"0c",	--760
		x"1c",	--761
		x"0c",	--762
		x"f9",	--763
		x"30",	--764
		x"86",	--765
		x"b0",	--766
		x"fc",	--767
		x"21",	--768
		x"3f",	--769
		x"3b",	--770
		x"30",	--771
		x"0c",	--772
		x"0c",	--773
		x"0c",	--774
		x"3c",	--775
		x"0a",	--776
		x"0f",	--777
		x"9c",	--778
		x"02",	--779
		x"3b",	--780
		x"30",	--781
		x"5e",	--782
		x"81",	--783
		x"3e",	--784
		x"fc",	--785
		x"c2",	--786
		x"19",	--787
		x"c2",	--788
		x"84",	--789
		x"0f",	--790
		x"30",	--791
		x"3f",	--792
		x"0f",	--793
		x"5f",	--794
		x"44",	--795
		x"8f",	--796
		x"b0",	--797
		x"1c",	--798
		x"30",	--799
		x"0b",	--800
		x"0b",	--801
		x"0e",	--802
		x"0e",	--803
		x"0e",	--804
		x"0e",	--805
		x"0e",	--806
		x"0f",	--807
		x"b0",	--808
		x"30",	--809
		x"0f",	--810
		x"b0",	--811
		x"30",	--812
		x"3b",	--813
		x"30",	--814
		x"0b",	--815
		x"0a",	--816
		x"0a",	--817
		x"3b",	--818
		x"07",	--819
		x"0e",	--820
		x"4d",	--821
		x"7d",	--822
		x"0f",	--823
		x"03",	--824
		x"0e",	--825
		x"7d",	--826
		x"fd",	--827
		x"1e",	--828
		x"0a",	--829
		x"3f",	--830
		x"31",	--831
		x"b0",	--832
		x"1c",	--833
		x"3b",	--834
		x"3b",	--835
		x"ef",	--836
		x"3a",	--837
		x"3b",	--838
		x"30",	--839
		x"3f",	--840
		x"30",	--841
		x"f5",	--842
		x"0b",	--843
		x"0b",	--844
		x"0e",	--845
		x"8e",	--846
		x"8e",	--847
		x"0f",	--848
		x"b0",	--849
		x"40",	--850
		x"0f",	--851
		x"b0",	--852
		x"40",	--853
		x"3b",	--854
		x"30",	--855
		x"0b",	--856
		x"0a",	--857
		x"0a",	--858
		x"0b",	--859
		x"0d",	--860
		x"8d",	--861
		x"8d",	--862
		x"0f",	--863
		x"b0",	--864
		x"40",	--865
		x"0f",	--866
		x"b0",	--867
		x"40",	--868
		x"0c",	--869
		x"0d",	--870
		x"8d",	--871
		x"8c",	--872
		x"4d",	--873
		x"0d",	--874
		x"0f",	--875
		x"b0",	--876
		x"40",	--877
		x"0f",	--878
		x"b0",	--879
		x"40",	--880
		x"3a",	--881
		x"3b",	--882
		x"30",	--883
		x"0b",	--884
		x"0a",	--885
		x"09",	--886
		x"0a",	--887
		x"0e",	--888
		x"19",	--889
		x"09",	--890
		x"39",	--891
		x"0b",	--892
		x"0d",	--893
		x"0d",	--894
		x"6f",	--895
		x"8f",	--896
		x"b0",	--897
		x"40",	--898
		x"0b",	--899
		x"0e",	--900
		x"1b",	--901
		x"3b",	--902
		x"07",	--903
		x"05",	--904
		x"3f",	--905
		x"20",	--906
		x"b0",	--907
		x"1c",	--908
		x"ef",	--909
		x"3f",	--910
		x"3a",	--911
		x"b0",	--912
		x"1c",	--913
		x"ea",	--914
		x"39",	--915
		x"3a",	--916
		x"3b",	--917
		x"30",	--918
		x"0b",	--919
		x"0a",	--920
		x"09",	--921
		x"0a",	--922
		x"0e",	--923
		x"17",	--924
		x"09",	--925
		x"39",	--926
		x"0b",	--927
		x"6f",	--928
		x"8f",	--929
		x"b0",	--930
		x"30",	--931
		x"0b",	--932
		x"0e",	--933
		x"1b",	--934
		x"3b",	--935
		x"07",	--936
		x"f6",	--937
		x"3f",	--938
		x"20",	--939
		x"b0",	--940
		x"1c",	--941
		x"6f",	--942
		x"8f",	--943
		x"b0",	--944
		x"30",	--945
		x"0b",	--946
		x"f2",	--947
		x"39",	--948
		x"3a",	--949
		x"3b",	--950
		x"30",	--951
		x"0b",	--952
		x"0a",	--953
		x"09",	--954
		x"31",	--955
		x"ec",	--956
		x"0b",	--957
		x"0f",	--958
		x"34",	--959
		x"3b",	--960
		x"0a",	--961
		x"38",	--962
		x"09",	--963
		x"0a",	--964
		x"0a",	--965
		x"3e",	--966
		x"0a",	--967
		x"0f",	--968
		x"b0",	--969
		x"92",	--970
		x"7f",	--971
		x"30",	--972
		x"ca",	--973
		x"00",	--974
		x"19",	--975
		x"3e",	--976
		x"0a",	--977
		x"0f",	--978
		x"b0",	--979
		x"60",	--980
		x"0b",	--981
		x"3f",	--982
		x"0a",	--983
		x"eb",	--984
		x"0a",	--985
		x"1a",	--986
		x"09",	--987
		x"3e",	--988
		x"0a",	--989
		x"0f",	--990
		x"b0",	--991
		x"92",	--992
		x"7f",	--993
		x"30",	--994
		x"c9",	--995
		x"00",	--996
		x"3a",	--997
		x"0f",	--998
		x"0f",	--999
		x"6f",	--1000
		x"8f",	--1001
		x"b0",	--1002
		x"1c",	--1003
		x"0a",	--1004
		x"f7",	--1005
		x"31",	--1006
		x"14",	--1007
		x"39",	--1008
		x"3a",	--1009
		x"3b",	--1010
		x"30",	--1011
		x"3f",	--1012
		x"2d",	--1013
		x"b0",	--1014
		x"1c",	--1015
		x"3b",	--1016
		x"1b",	--1017
		x"c5",	--1018
		x"1a",	--1019
		x"09",	--1020
		x"dd",	--1021
		x"0b",	--1022
		x"0a",	--1023
		x"09",	--1024
		x"0b",	--1025
		x"3b",	--1026
		x"39",	--1027
		x"6f",	--1028
		x"4f",	--1029
		x"0b",	--1030
		x"1a",	--1031
		x"8f",	--1032
		x"b0",	--1033
		x"1c",	--1034
		x"0a",	--1035
		x"09",	--1036
		x"19",	--1037
		x"5f",	--1038
		x"01",	--1039
		x"4f",	--1040
		x"10",	--1041
		x"7f",	--1042
		x"25",	--1043
		x"f3",	--1044
		x"0a",	--1045
		x"1a",	--1046
		x"5f",	--1047
		x"01",	--1048
		x"7f",	--1049
		x"db",	--1050
		x"7f",	--1051
		x"54",	--1052
		x"ee",	--1053
		x"4f",	--1054
		x"0f",	--1055
		x"10",	--1056
		x"9c",	--1057
		x"39",	--1058
		x"3a",	--1059
		x"3b",	--1060
		x"30",	--1061
		x"09",	--1062
		x"29",	--1063
		x"1e",	--1064
		x"02",	--1065
		x"2f",	--1066
		x"b0",	--1067
		x"e8",	--1068
		x"0b",	--1069
		x"dd",	--1070
		x"09",	--1071
		x"29",	--1072
		x"2f",	--1073
		x"b0",	--1074
		x"96",	--1075
		x"0b",	--1076
		x"d6",	--1077
		x"0f",	--1078
		x"2b",	--1079
		x"29",	--1080
		x"6f",	--1081
		x"4f",	--1082
		x"d0",	--1083
		x"19",	--1084
		x"8f",	--1085
		x"b0",	--1086
		x"1c",	--1087
		x"7f",	--1088
		x"4f",	--1089
		x"fa",	--1090
		x"c8",	--1091
		x"09",	--1092
		x"29",	--1093
		x"1e",	--1094
		x"02",	--1095
		x"2f",	--1096
		x"b0",	--1097
		x"2e",	--1098
		x"0b",	--1099
		x"bf",	--1100
		x"09",	--1101
		x"29",	--1102
		x"2e",	--1103
		x"0f",	--1104
		x"8f",	--1105
		x"8f",	--1106
		x"8f",	--1107
		x"8f",	--1108
		x"b0",	--1109
		x"b0",	--1110
		x"0b",	--1111
		x"b3",	--1112
		x"09",	--1113
		x"29",	--1114
		x"2f",	--1115
		x"b0",	--1116
		x"70",	--1117
		x"0b",	--1118
		x"ac",	--1119
		x"09",	--1120
		x"29",	--1121
		x"2f",	--1122
		x"b0",	--1123
		x"1c",	--1124
		x"0b",	--1125
		x"a5",	--1126
		x"09",	--1127
		x"29",	--1128
		x"2f",	--1129
		x"b0",	--1130
		x"40",	--1131
		x"0b",	--1132
		x"9e",	--1133
		x"09",	--1134
		x"29",	--1135
		x"2f",	--1136
		x"b0",	--1137
		x"5e",	--1138
		x"0b",	--1139
		x"97",	--1140
		x"3f",	--1141
		x"25",	--1142
		x"b0",	--1143
		x"1c",	--1144
		x"92",	--1145
		x"0f",	--1146
		x"0e",	--1147
		x"1f",	--1148
		x"02",	--1149
		x"df",	--1150
		x"85",	--1151
		x"0a",	--1152
		x"1f",	--1153
		x"02",	--1154
		x"3f",	--1155
		x"3f",	--1156
		x"16",	--1157
		x"92",	--1158
		x"02",	--1159
		x"1e",	--1160
		x"02",	--1161
		x"1f",	--1162
		x"04",	--1163
		x"0e",	--1164
		x"02",	--1165
		x"92",	--1166
		x"04",	--1167
		x"f2",	--1168
		x"10",	--1169
		x"81",	--1170
		x"b1",	--1171
		x"10",	--1172
		x"04",	--1173
		x"3e",	--1174
		x"3f",	--1175
		x"b1",	--1176
		x"f0",	--1177
		x"00",	--1178
		x"00",	--1179
		x"82",	--1180
		x"02",	--1181
		x"e9",	--1182
		x"b2",	--1183
		x"c3",	--1184
		x"82",	--1185
		x"f2",	--1186
		x"11",	--1187
		x"80",	--1188
		x"30",	--1189
		x"1e",	--1190
		x"02",	--1191
		x"1f",	--1192
		x"04",	--1193
		x"0e",	--1194
		x"05",	--1195
		x"1f",	--1196
		x"02",	--1197
		x"1f",	--1198
		x"04",	--1199
		x"30",	--1200
		x"1d",	--1201
		x"02",	--1202
		x"1e",	--1203
		x"04",	--1204
		x"3f",	--1205
		x"40",	--1206
		x"0f",	--1207
		x"0f",	--1208
		x"30",	--1209
		x"1f",	--1210
		x"04",	--1211
		x"5f",	--1212
		x"0a",	--1213
		x"1d",	--1214
		x"04",	--1215
		x"1e",	--1216
		x"02",	--1217
		x"0d",	--1218
		x"0b",	--1219
		x"1e",	--1220
		x"04",	--1221
		x"3e",	--1222
		x"3f",	--1223
		x"03",	--1224
		x"82",	--1225
		x"04",	--1226
		x"30",	--1227
		x"92",	--1228
		x"04",	--1229
		x"30",	--1230
		x"4f",	--1231
		x"30",	--1232
		x"0b",	--1233
		x"0a",	--1234
		x"0a",	--1235
		x"0b",	--1236
		x"0c",	--1237
		x"3d",	--1238
		x"00",	--1239
		x"b0",	--1240
		x"86",	--1241
		x"0f",	--1242
		x"07",	--1243
		x"0e",	--1244
		x"0f",	--1245
		x"b0",	--1246
		x"d6",	--1247
		x"3a",	--1248
		x"3b",	--1249
		x"30",	--1250
		x"0c",	--1251
		x"3d",	--1252
		x"00",	--1253
		x"0e",	--1254
		x"0f",	--1255
		x"b0",	--1256
		x"c2",	--1257
		x"b0",	--1258
		x"d6",	--1259
		x"0e",	--1260
		x"3f",	--1261
		x"00",	--1262
		x"3a",	--1263
		x"3b",	--1264
		x"30",	--1265
		x"0b",	--1266
		x"0a",	--1267
		x"09",	--1268
		x"08",	--1269
		x"07",	--1270
		x"06",	--1271
		x"05",	--1272
		x"04",	--1273
		x"31",	--1274
		x"fa",	--1275
		x"08",	--1276
		x"6b",	--1277
		x"6b",	--1278
		x"67",	--1279
		x"6c",	--1280
		x"6c",	--1281
		x"e9",	--1282
		x"6b",	--1283
		x"02",	--1284
		x"30",	--1285
		x"64",	--1286
		x"6c",	--1287
		x"e3",	--1288
		x"6c",	--1289
		x"bb",	--1290
		x"6b",	--1291
		x"df",	--1292
		x"91",	--1293
		x"02",	--1294
		x"00",	--1295
		x"1b",	--1296
		x"02",	--1297
		x"14",	--1298
		x"04",	--1299
		x"15",	--1300
		x"06",	--1301
		x"16",	--1302
		x"04",	--1303
		x"17",	--1304
		x"06",	--1305
		x"2c",	--1306
		x"0c",	--1307
		x"09",	--1308
		x"0c",	--1309
		x"bf",	--1310
		x"39",	--1311
		x"20",	--1312
		x"50",	--1313
		x"1c",	--1314
		x"d7",	--1315
		x"81",	--1316
		x"02",	--1317
		x"81",	--1318
		x"04",	--1319
		x"4c",	--1320
		x"7c",	--1321
		x"1f",	--1322
		x"0b",	--1323
		x"0a",	--1324
		x"0b",	--1325
		x"12",	--1326
		x"0b",	--1327
		x"0a",	--1328
		x"7c",	--1329
		x"fb",	--1330
		x"81",	--1331
		x"02",	--1332
		x"81",	--1333
		x"04",	--1334
		x"1c",	--1335
		x"0d",	--1336
		x"79",	--1337
		x"1f",	--1338
		x"04",	--1339
		x"0c",	--1340
		x"0d",	--1341
		x"79",	--1342
		x"fc",	--1343
		x"3c",	--1344
		x"3d",	--1345
		x"0c",	--1346
		x"0d",	--1347
		x"1a",	--1348
		x"0b",	--1349
		x"0c",	--1350
		x"02",	--1351
		x"0d",	--1352
		x"e5",	--1353
		x"16",	--1354
		x"02",	--1355
		x"17",	--1356
		x"04",	--1357
		x"06",	--1358
		x"07",	--1359
		x"5f",	--1360
		x"01",	--1361
		x"5f",	--1362
		x"01",	--1363
		x"28",	--1364
		x"c8",	--1365
		x"01",	--1366
		x"a8",	--1367
		x"02",	--1368
		x"0e",	--1369
		x"0f",	--1370
		x"0e",	--1371
		x"0f",	--1372
		x"88",	--1373
		x"04",	--1374
		x"88",	--1375
		x"06",	--1376
		x"f8",	--1377
		x"03",	--1378
		x"00",	--1379
		x"0f",	--1380
		x"4d",	--1381
		x"0f",	--1382
		x"31",	--1383
		x"06",	--1384
		x"34",	--1385
		x"35",	--1386
		x"36",	--1387
		x"37",	--1388
		x"38",	--1389
		x"39",	--1390
		x"3a",	--1391
		x"3b",	--1392
		x"30",	--1393
		x"2b",	--1394
		x"67",	--1395
		x"81",	--1396
		x"00",	--1397
		x"04",	--1398
		x"05",	--1399
		x"5f",	--1400
		x"01",	--1401
		x"5f",	--1402
		x"01",	--1403
		x"d8",	--1404
		x"4f",	--1405
		x"68",	--1406
		x"0e",	--1407
		x"0f",	--1408
		x"0e",	--1409
		x"0f",	--1410
		x"0f",	--1411
		x"69",	--1412
		x"c8",	--1413
		x"01",	--1414
		x"a8",	--1415
		x"02",	--1416
		x"88",	--1417
		x"04",	--1418
		x"88",	--1419
		x"06",	--1420
		x"0c",	--1421
		x"0d",	--1422
		x"3c",	--1423
		x"3d",	--1424
		x"3d",	--1425
		x"ff",	--1426
		x"05",	--1427
		x"3d",	--1428
		x"00",	--1429
		x"17",	--1430
		x"3c",	--1431
		x"15",	--1432
		x"1b",	--1433
		x"02",	--1434
		x"3b",	--1435
		x"0e",	--1436
		x"0f",	--1437
		x"0a",	--1438
		x"3b",	--1439
		x"0c",	--1440
		x"0d",	--1441
		x"3c",	--1442
		x"3d",	--1443
		x"3d",	--1444
		x"ff",	--1445
		x"f5",	--1446
		x"3c",	--1447
		x"88",	--1448
		x"04",	--1449
		x"88",	--1450
		x"06",	--1451
		x"88",	--1452
		x"02",	--1453
		x"f8",	--1454
		x"03",	--1455
		x"00",	--1456
		x"0f",	--1457
		x"b3",	--1458
		x"0c",	--1459
		x"0d",	--1460
		x"1c",	--1461
		x"0d",	--1462
		x"12",	--1463
		x"0f",	--1464
		x"0e",	--1465
		x"0a",	--1466
		x"0b",	--1467
		x"0a",	--1468
		x"0b",	--1469
		x"88",	--1470
		x"04",	--1471
		x"88",	--1472
		x"06",	--1473
		x"98",	--1474
		x"02",	--1475
		x"0f",	--1476
		x"a1",	--1477
		x"6b",	--1478
		x"9f",	--1479
		x"ad",	--1480
		x"00",	--1481
		x"9d",	--1482
		x"02",	--1483
		x"02",	--1484
		x"9d",	--1485
		x"04",	--1486
		x"04",	--1487
		x"9d",	--1488
		x"06",	--1489
		x"06",	--1490
		x"5e",	--1491
		x"01",	--1492
		x"5e",	--1493
		x"01",	--1494
		x"cd",	--1495
		x"01",	--1496
		x"0f",	--1497
		x"8c",	--1498
		x"06",	--1499
		x"07",	--1500
		x"9a",	--1501
		x"39",	--1502
		x"19",	--1503
		x"39",	--1504
		x"20",	--1505
		x"8f",	--1506
		x"3e",	--1507
		x"3c",	--1508
		x"b6",	--1509
		x"c1",	--1510
		x"0e",	--1511
		x"0f",	--1512
		x"0e",	--1513
		x"0f",	--1514
		x"97",	--1515
		x"0f",	--1516
		x"79",	--1517
		x"d8",	--1518
		x"01",	--1519
		x"a8",	--1520
		x"02",	--1521
		x"3e",	--1522
		x"3f",	--1523
		x"1e",	--1524
		x"0f",	--1525
		x"88",	--1526
		x"04",	--1527
		x"88",	--1528
		x"06",	--1529
		x"92",	--1530
		x"0c",	--1531
		x"7b",	--1532
		x"81",	--1533
		x"00",	--1534
		x"81",	--1535
		x"02",	--1536
		x"81",	--1537
		x"04",	--1538
		x"4d",	--1539
		x"7d",	--1540
		x"1f",	--1541
		x"0c",	--1542
		x"4b",	--1543
		x"0c",	--1544
		x"0d",	--1545
		x"12",	--1546
		x"0d",	--1547
		x"0c",	--1548
		x"7b",	--1549
		x"fb",	--1550
		x"81",	--1551
		x"02",	--1552
		x"81",	--1553
		x"04",	--1554
		x"1c",	--1555
		x"0d",	--1556
		x"79",	--1557
		x"1f",	--1558
		x"04",	--1559
		x"0c",	--1560
		x"0d",	--1561
		x"79",	--1562
		x"fc",	--1563
		x"3c",	--1564
		x"3d",	--1565
		x"0c",	--1566
		x"0d",	--1567
		x"1a",	--1568
		x"0b",	--1569
		x"0c",	--1570
		x"04",	--1571
		x"0d",	--1572
		x"02",	--1573
		x"0a",	--1574
		x"0b",	--1575
		x"14",	--1576
		x"02",	--1577
		x"15",	--1578
		x"04",	--1579
		x"04",	--1580
		x"05",	--1581
		x"49",	--1582
		x"0a",	--1583
		x"0b",	--1584
		x"18",	--1585
		x"6c",	--1586
		x"33",	--1587
		x"df",	--1588
		x"01",	--1589
		x"01",	--1590
		x"2f",	--1591
		x"3f",	--1592
		x"56",	--1593
		x"2c",	--1594
		x"31",	--1595
		x"e0",	--1596
		x"81",	--1597
		x"04",	--1598
		x"81",	--1599
		x"06",	--1600
		x"81",	--1601
		x"00",	--1602
		x"81",	--1603
		x"02",	--1604
		x"0e",	--1605
		x"3e",	--1606
		x"18",	--1607
		x"0f",	--1608
		x"2f",	--1609
		x"b0",	--1610
		x"98",	--1611
		x"0e",	--1612
		x"3e",	--1613
		x"10",	--1614
		x"0f",	--1615
		x"b0",	--1616
		x"98",	--1617
		x"0d",	--1618
		x"3d",	--1619
		x"0e",	--1620
		x"3e",	--1621
		x"10",	--1622
		x"0f",	--1623
		x"3f",	--1624
		x"18",	--1625
		x"b0",	--1626
		x"e4",	--1627
		x"b0",	--1628
		x"ba",	--1629
		x"31",	--1630
		x"20",	--1631
		x"30",	--1632
		x"31",	--1633
		x"e0",	--1634
		x"81",	--1635
		x"04",	--1636
		x"81",	--1637
		x"06",	--1638
		x"81",	--1639
		x"00",	--1640
		x"81",	--1641
		x"02",	--1642
		x"0e",	--1643
		x"3e",	--1644
		x"18",	--1645
		x"0f",	--1646
		x"2f",	--1647
		x"b0",	--1648
		x"98",	--1649
		x"0e",	--1650
		x"3e",	--1651
		x"10",	--1652
		x"0f",	--1653
		x"b0",	--1654
		x"98",	--1655
		x"d1",	--1656
		x"11",	--1657
		x"0d",	--1658
		x"3d",	--1659
		x"0e",	--1660
		x"3e",	--1661
		x"10",	--1662
		x"0f",	--1663
		x"3f",	--1664
		x"18",	--1665
		x"b0",	--1666
		x"e4",	--1667
		x"b0",	--1668
		x"ba",	--1669
		x"31",	--1670
		x"20",	--1671
		x"30",	--1672
		x"0b",	--1673
		x"0a",	--1674
		x"09",	--1675
		x"08",	--1676
		x"07",	--1677
		x"06",	--1678
		x"05",	--1679
		x"04",	--1680
		x"31",	--1681
		x"dc",	--1682
		x"81",	--1683
		x"04",	--1684
		x"81",	--1685
		x"06",	--1686
		x"81",	--1687
		x"00",	--1688
		x"81",	--1689
		x"02",	--1690
		x"0e",	--1691
		x"3e",	--1692
		x"18",	--1693
		x"0f",	--1694
		x"2f",	--1695
		x"b0",	--1696
		x"98",	--1697
		x"0e",	--1698
		x"3e",	--1699
		x"10",	--1700
		x"0f",	--1701
		x"b0",	--1702
		x"98",	--1703
		x"5f",	--1704
		x"18",	--1705
		x"6f",	--1706
		x"b6",	--1707
		x"5e",	--1708
		x"10",	--1709
		x"6e",	--1710
		x"d9",	--1711
		x"6f",	--1712
		x"ae",	--1713
		x"6e",	--1714
		x"e2",	--1715
		x"6f",	--1716
		x"ac",	--1717
		x"6e",	--1718
		x"d1",	--1719
		x"14",	--1720
		x"1c",	--1721
		x"15",	--1722
		x"1e",	--1723
		x"18",	--1724
		x"14",	--1725
		x"19",	--1726
		x"16",	--1727
		x"3c",	--1728
		x"20",	--1729
		x"0e",	--1730
		x"0f",	--1731
		x"06",	--1732
		x"07",	--1733
		x"81",	--1734
		x"20",	--1735
		x"81",	--1736
		x"22",	--1737
		x"0a",	--1738
		x"0b",	--1739
		x"81",	--1740
		x"20",	--1741
		x"08",	--1742
		x"08",	--1743
		x"09",	--1744
		x"12",	--1745
		x"05",	--1746
		x"04",	--1747
		x"b1",	--1748
		x"20",	--1749
		x"19",	--1750
		x"14",	--1751
		x"0d",	--1752
		x"0a",	--1753
		x"0b",	--1754
		x"0e",	--1755
		x"0f",	--1756
		x"1c",	--1757
		x"0d",	--1758
		x"0b",	--1759
		x"03",	--1760
		x"0b",	--1761
		x"0c",	--1762
		x"0d",	--1763
		x"0e",	--1764
		x"0f",	--1765
		x"06",	--1766
		x"07",	--1767
		x"09",	--1768
		x"e5",	--1769
		x"16",	--1770
		x"07",	--1771
		x"e2",	--1772
		x"0a",	--1773
		x"f5",	--1774
		x"f2",	--1775
		x"81",	--1776
		x"20",	--1777
		x"81",	--1778
		x"22",	--1779
		x"0c",	--1780
		x"1a",	--1781
		x"1a",	--1782
		x"1a",	--1783
		x"12",	--1784
		x"06",	--1785
		x"26",	--1786
		x"81",	--1787
		x"0a",	--1788
		x"5d",	--1789
		x"d1",	--1790
		x"11",	--1791
		x"19",	--1792
		x"83",	--1793
		x"c1",	--1794
		x"09",	--1795
		x"0c",	--1796
		x"3c",	--1797
		x"3f",	--1798
		x"00",	--1799
		x"18",	--1800
		x"1d",	--1801
		x"0a",	--1802
		x"3d",	--1803
		x"1a",	--1804
		x"20",	--1805
		x"1b",	--1806
		x"22",	--1807
		x"0c",	--1808
		x"0e",	--1809
		x"0f",	--1810
		x"0b",	--1811
		x"2a",	--1812
		x"0a",	--1813
		x"0b",	--1814
		x"3d",	--1815
		x"3f",	--1816
		x"00",	--1817
		x"f5",	--1818
		x"81",	--1819
		x"20",	--1820
		x"81",	--1821
		x"22",	--1822
		x"81",	--1823
		x"0a",	--1824
		x"0c",	--1825
		x"0d",	--1826
		x"3c",	--1827
		x"7f",	--1828
		x"0d",	--1829
		x"3c",	--1830
		x"40",	--1831
		x"44",	--1832
		x"81",	--1833
		x"0c",	--1834
		x"81",	--1835
		x"0e",	--1836
		x"f1",	--1837
		x"03",	--1838
		x"08",	--1839
		x"0f",	--1840
		x"3f",	--1841
		x"b0",	--1842
		x"ba",	--1843
		x"31",	--1844
		x"24",	--1845
		x"34",	--1846
		x"35",	--1847
		x"36",	--1848
		x"37",	--1849
		x"38",	--1850
		x"39",	--1851
		x"3a",	--1852
		x"3b",	--1853
		x"30",	--1854
		x"1e",	--1855
		x"0f",	--1856
		x"d3",	--1857
		x"3a",	--1858
		x"03",	--1859
		x"08",	--1860
		x"1e",	--1861
		x"10",	--1862
		x"1c",	--1863
		x"20",	--1864
		x"1d",	--1865
		x"22",	--1866
		x"12",	--1867
		x"0d",	--1868
		x"0c",	--1869
		x"06",	--1870
		x"07",	--1871
		x"06",	--1872
		x"37",	--1873
		x"00",	--1874
		x"81",	--1875
		x"20",	--1876
		x"81",	--1877
		x"22",	--1878
		x"12",	--1879
		x"0f",	--1880
		x"0e",	--1881
		x"1a",	--1882
		x"0f",	--1883
		x"e7",	--1884
		x"81",	--1885
		x"0a",	--1886
		x"a6",	--1887
		x"6e",	--1888
		x"36",	--1889
		x"5f",	--1890
		x"d1",	--1891
		x"11",	--1892
		x"19",	--1893
		x"20",	--1894
		x"c1",	--1895
		x"19",	--1896
		x"0f",	--1897
		x"3f",	--1898
		x"18",	--1899
		x"c5",	--1900
		x"0d",	--1901
		x"ba",	--1902
		x"0c",	--1903
		x"0d",	--1904
		x"3c",	--1905
		x"80",	--1906
		x"0d",	--1907
		x"0c",	--1908
		x"b3",	--1909
		x"0d",	--1910
		x"b1",	--1911
		x"81",	--1912
		x"20",	--1913
		x"03",	--1914
		x"81",	--1915
		x"22",	--1916
		x"ab",	--1917
		x"3e",	--1918
		x"40",	--1919
		x"0f",	--1920
		x"3e",	--1921
		x"80",	--1922
		x"3f",	--1923
		x"a4",	--1924
		x"4d",	--1925
		x"7b",	--1926
		x"4f",	--1927
		x"de",	--1928
		x"5f",	--1929
		x"d1",	--1930
		x"11",	--1931
		x"19",	--1932
		x"06",	--1933
		x"c1",	--1934
		x"11",	--1935
		x"0f",	--1936
		x"3f",	--1937
		x"10",	--1938
		x"9e",	--1939
		x"4f",	--1940
		x"f8",	--1941
		x"6f",	--1942
		x"f1",	--1943
		x"3f",	--1944
		x"56",	--1945
		x"97",	--1946
		x"0b",	--1947
		x"0a",	--1948
		x"09",	--1949
		x"08",	--1950
		x"07",	--1951
		x"31",	--1952
		x"e8",	--1953
		x"81",	--1954
		x"04",	--1955
		x"81",	--1956
		x"06",	--1957
		x"81",	--1958
		x"00",	--1959
		x"81",	--1960
		x"02",	--1961
		x"0e",	--1962
		x"3e",	--1963
		x"10",	--1964
		x"0f",	--1965
		x"2f",	--1966
		x"b0",	--1967
		x"98",	--1968
		x"0e",	--1969
		x"3e",	--1970
		x"0f",	--1971
		x"b0",	--1972
		x"98",	--1973
		x"5f",	--1974
		x"10",	--1975
		x"6f",	--1976
		x"5d",	--1977
		x"5e",	--1978
		x"08",	--1979
		x"6e",	--1980
		x"82",	--1981
		x"d1",	--1982
		x"09",	--1983
		x"11",	--1984
		x"6f",	--1985
		x"58",	--1986
		x"6f",	--1987
		x"56",	--1988
		x"6e",	--1989
		x"6f",	--1990
		x"6e",	--1991
		x"4c",	--1992
		x"1d",	--1993
		x"12",	--1994
		x"1d",	--1995
		x"0a",	--1996
		x"81",	--1997
		x"12",	--1998
		x"1e",	--1999
		x"14",	--2000
		x"1f",	--2001
		x"16",	--2002
		x"18",	--2003
		x"0c",	--2004
		x"19",	--2005
		x"0e",	--2006
		x"0f",	--2007
		x"1e",	--2008
		x"0e",	--2009
		x"0f",	--2010
		x"3d",	--2011
		x"81",	--2012
		x"12",	--2013
		x"37",	--2014
		x"1f",	--2015
		x"0c",	--2016
		x"3d",	--2017
		x"00",	--2018
		x"0a",	--2019
		x"0b",	--2020
		x"0b",	--2021
		x"0a",	--2022
		x"0b",	--2023
		x"0e",	--2024
		x"0f",	--2025
		x"12",	--2026
		x"0d",	--2027
		x"0c",	--2028
		x"0e",	--2029
		x"0f",	--2030
		x"37",	--2031
		x"0b",	--2032
		x"0f",	--2033
		x"f7",	--2034
		x"f2",	--2035
		x"0e",	--2036
		x"f4",	--2037
		x"ef",	--2038
		x"09",	--2039
		x"e5",	--2040
		x"0e",	--2041
		x"e3",	--2042
		x"dd",	--2043
		x"0c",	--2044
		x"0d",	--2045
		x"3c",	--2046
		x"7f",	--2047
		x"0d",	--2048
		x"3c",	--2049
		x"40",	--2050
		x"1c",	--2051
		x"81",	--2052
		x"14",	--2053
		x"81",	--2054
		x"16",	--2055
		x"0f",	--2056
		x"3f",	--2057
		x"10",	--2058
		x"b0",	--2059
		x"ba",	--2060
		x"31",	--2061
		x"18",	--2062
		x"37",	--2063
		x"38",	--2064
		x"39",	--2065
		x"3a",	--2066
		x"3b",	--2067
		x"30",	--2068
		x"e1",	--2069
		x"10",	--2070
		x"0f",	--2071
		x"3f",	--2072
		x"10",	--2073
		x"f0",	--2074
		x"4f",	--2075
		x"fa",	--2076
		x"3f",	--2077
		x"56",	--2078
		x"eb",	--2079
		x"0d",	--2080
		x"e2",	--2081
		x"0c",	--2082
		x"0d",	--2083
		x"3c",	--2084
		x"80",	--2085
		x"0d",	--2086
		x"0c",	--2087
		x"db",	--2088
		x"0d",	--2089
		x"d9",	--2090
		x"0e",	--2091
		x"02",	--2092
		x"0f",	--2093
		x"d5",	--2094
		x"3a",	--2095
		x"40",	--2096
		x"0b",	--2097
		x"3a",	--2098
		x"80",	--2099
		x"3b",	--2100
		x"ce",	--2101
		x"81",	--2102
		x"14",	--2103
		x"81",	--2104
		x"16",	--2105
		x"81",	--2106
		x"12",	--2107
		x"0f",	--2108
		x"3f",	--2109
		x"10",	--2110
		x"cb",	--2111
		x"0f",	--2112
		x"3f",	--2113
		x"c8",	--2114
		x"31",	--2115
		x"e8",	--2116
		x"81",	--2117
		x"04",	--2118
		x"81",	--2119
		x"06",	--2120
		x"81",	--2121
		x"00",	--2122
		x"81",	--2123
		x"02",	--2124
		x"0e",	--2125
		x"3e",	--2126
		x"10",	--2127
		x"0f",	--2128
		x"2f",	--2129
		x"b0",	--2130
		x"98",	--2131
		x"0e",	--2132
		x"3e",	--2133
		x"0f",	--2134
		x"b0",	--2135
		x"98",	--2136
		x"e1",	--2137
		x"10",	--2138
		x"0d",	--2139
		x"e1",	--2140
		x"08",	--2141
		x"0a",	--2142
		x"0e",	--2143
		x"3e",	--2144
		x"0f",	--2145
		x"3f",	--2146
		x"10",	--2147
		x"b0",	--2148
		x"bc",	--2149
		x"31",	--2150
		x"18",	--2151
		x"30",	--2152
		x"3f",	--2153
		x"fb",	--2154
		x"31",	--2155
		x"f4",	--2156
		x"81",	--2157
		x"00",	--2158
		x"81",	--2159
		x"02",	--2160
		x"0e",	--2161
		x"2e",	--2162
		x"0f",	--2163
		x"b0",	--2164
		x"98",	--2165
		x"5f",	--2166
		x"04",	--2167
		x"6f",	--2168
		x"28",	--2169
		x"27",	--2170
		x"6f",	--2171
		x"07",	--2172
		x"1d",	--2173
		x"06",	--2174
		x"0d",	--2175
		x"21",	--2176
		x"3d",	--2177
		x"1f",	--2178
		x"09",	--2179
		x"c1",	--2180
		x"05",	--2181
		x"26",	--2182
		x"3e",	--2183
		x"3f",	--2184
		x"ff",	--2185
		x"31",	--2186
		x"0c",	--2187
		x"30",	--2188
		x"1e",	--2189
		x"08",	--2190
		x"1f",	--2191
		x"0a",	--2192
		x"3c",	--2193
		x"1e",	--2194
		x"4c",	--2195
		x"4d",	--2196
		x"7d",	--2197
		x"1f",	--2198
		x"0f",	--2199
		x"c1",	--2200
		x"05",	--2201
		x"ef",	--2202
		x"3e",	--2203
		x"3f",	--2204
		x"1e",	--2205
		x"0f",	--2206
		x"31",	--2207
		x"0c",	--2208
		x"30",	--2209
		x"0e",	--2210
		x"0f",	--2211
		x"31",	--2212
		x"0c",	--2213
		x"30",	--2214
		x"12",	--2215
		x"0f",	--2216
		x"0e",	--2217
		x"7d",	--2218
		x"fb",	--2219
		x"eb",	--2220
		x"0e",	--2221
		x"3f",	--2222
		x"00",	--2223
		x"31",	--2224
		x"0c",	--2225
		x"30",	--2226
		x"0b",	--2227
		x"0a",	--2228
		x"09",	--2229
		x"08",	--2230
		x"31",	--2231
		x"0a",	--2232
		x"0b",	--2233
		x"c1",	--2234
		x"01",	--2235
		x"0e",	--2236
		x"0d",	--2237
		x"0b",	--2238
		x"0b",	--2239
		x"e1",	--2240
		x"00",	--2241
		x"0f",	--2242
		x"b0",	--2243
		x"ba",	--2244
		x"31",	--2245
		x"38",	--2246
		x"39",	--2247
		x"3a",	--2248
		x"3b",	--2249
		x"30",	--2250
		x"f1",	--2251
		x"03",	--2252
		x"00",	--2253
		x"b1",	--2254
		x"1e",	--2255
		x"02",	--2256
		x"81",	--2257
		x"04",	--2258
		x"81",	--2259
		x"06",	--2260
		x"0e",	--2261
		x"0f",	--2262
		x"b0",	--2263
		x"48",	--2264
		x"3f",	--2265
		x"0f",	--2266
		x"18",	--2267
		x"e5",	--2268
		x"81",	--2269
		x"04",	--2270
		x"81",	--2271
		x"06",	--2272
		x"4e",	--2273
		x"7e",	--2274
		x"1f",	--2275
		x"06",	--2276
		x"3e",	--2277
		x"1e",	--2278
		x"0e",	--2279
		x"81",	--2280
		x"02",	--2281
		x"d7",	--2282
		x"91",	--2283
		x"04",	--2284
		x"04",	--2285
		x"91",	--2286
		x"06",	--2287
		x"06",	--2288
		x"7e",	--2289
		x"f8",	--2290
		x"f1",	--2291
		x"0e",	--2292
		x"3e",	--2293
		x"1e",	--2294
		x"1c",	--2295
		x"0d",	--2296
		x"48",	--2297
		x"78",	--2298
		x"1f",	--2299
		x"04",	--2300
		x"0c",	--2301
		x"0d",	--2302
		x"78",	--2303
		x"fc",	--2304
		x"3c",	--2305
		x"3d",	--2306
		x"0c",	--2307
		x"0d",	--2308
		x"18",	--2309
		x"09",	--2310
		x"0c",	--2311
		x"04",	--2312
		x"0d",	--2313
		x"02",	--2314
		x"08",	--2315
		x"09",	--2316
		x"7e",	--2317
		x"1f",	--2318
		x"0e",	--2319
		x"0d",	--2320
		x"0e",	--2321
		x"0d",	--2322
		x"0e",	--2323
		x"81",	--2324
		x"04",	--2325
		x"81",	--2326
		x"06",	--2327
		x"3e",	--2328
		x"1e",	--2329
		x"0e",	--2330
		x"81",	--2331
		x"02",	--2332
		x"a4",	--2333
		x"12",	--2334
		x"0b",	--2335
		x"0a",	--2336
		x"7e",	--2337
		x"fb",	--2338
		x"ec",	--2339
		x"0b",	--2340
		x"0a",	--2341
		x"09",	--2342
		x"1f",	--2343
		x"17",	--2344
		x"3e",	--2345
		x"00",	--2346
		x"2c",	--2347
		x"3a",	--2348
		x"18",	--2349
		x"0b",	--2350
		x"39",	--2351
		x"0c",	--2352
		x"0d",	--2353
		x"4f",	--2354
		x"4f",	--2355
		x"17",	--2356
		x"3c",	--2357
		x"5e",	--2358
		x"6e",	--2359
		x"0f",	--2360
		x"0a",	--2361
		x"0b",	--2362
		x"0f",	--2363
		x"39",	--2364
		x"3a",	--2365
		x"3b",	--2366
		x"30",	--2367
		x"3f",	--2368
		x"00",	--2369
		x"0f",	--2370
		x"3a",	--2371
		x"0b",	--2372
		x"39",	--2373
		x"18",	--2374
		x"0c",	--2375
		x"0d",	--2376
		x"4f",	--2377
		x"4f",	--2378
		x"e9",	--2379
		x"12",	--2380
		x"0d",	--2381
		x"0c",	--2382
		x"7f",	--2383
		x"fb",	--2384
		x"e3",	--2385
		x"3a",	--2386
		x"10",	--2387
		x"0b",	--2388
		x"39",	--2389
		x"10",	--2390
		x"ef",	--2391
		x"3a",	--2392
		x"20",	--2393
		x"0b",	--2394
		x"09",	--2395
		x"ea",	--2396
		x"0b",	--2397
		x"0a",	--2398
		x"09",	--2399
		x"08",	--2400
		x"07",	--2401
		x"0d",	--2402
		x"1e",	--2403
		x"04",	--2404
		x"1f",	--2405
		x"06",	--2406
		x"5a",	--2407
		x"01",	--2408
		x"6c",	--2409
		x"6c",	--2410
		x"70",	--2411
		x"6c",	--2412
		x"6a",	--2413
		x"6c",	--2414
		x"36",	--2415
		x"0e",	--2416
		x"32",	--2417
		x"1b",	--2418
		x"02",	--2419
		x"3b",	--2420
		x"82",	--2421
		x"6d",	--2422
		x"3b",	--2423
		x"80",	--2424
		x"5e",	--2425
		x"0c",	--2426
		x"0d",	--2427
		x"3c",	--2428
		x"7f",	--2429
		x"0d",	--2430
		x"3c",	--2431
		x"40",	--2432
		x"40",	--2433
		x"3e",	--2434
		x"3f",	--2435
		x"0f",	--2436
		x"0f",	--2437
		x"4a",	--2438
		x"0d",	--2439
		x"3d",	--2440
		x"7f",	--2441
		x"12",	--2442
		x"0f",	--2443
		x"0e",	--2444
		x"12",	--2445
		x"0f",	--2446
		x"0e",	--2447
		x"12",	--2448
		x"0f",	--2449
		x"0e",	--2450
		x"12",	--2451
		x"0f",	--2452
		x"0e",	--2453
		x"12",	--2454
		x"0f",	--2455
		x"0e",	--2456
		x"12",	--2457
		x"0f",	--2458
		x"0e",	--2459
		x"12",	--2460
		x"0f",	--2461
		x"0e",	--2462
		x"3e",	--2463
		x"3f",	--2464
		x"7f",	--2465
		x"4d",	--2466
		x"05",	--2467
		x"0f",	--2468
		x"cc",	--2469
		x"4d",	--2470
		x"0e",	--2471
		x"0f",	--2472
		x"4d",	--2473
		x"0d",	--2474
		x"0d",	--2475
		x"0d",	--2476
		x"0d",	--2477
		x"0d",	--2478
		x"0d",	--2479
		x"0d",	--2480
		x"0c",	--2481
		x"3c",	--2482
		x"7f",	--2483
		x"0c",	--2484
		x"4f",	--2485
		x"0f",	--2486
		x"0f",	--2487
		x"0f",	--2488
		x"0d",	--2489
		x"0d",	--2490
		x"0f",	--2491
		x"37",	--2492
		x"38",	--2493
		x"39",	--2494
		x"3a",	--2495
		x"3b",	--2496
		x"30",	--2497
		x"0d",	--2498
		x"be",	--2499
		x"0c",	--2500
		x"0d",	--2501
		x"3c",	--2502
		x"80",	--2503
		x"0d",	--2504
		x"0c",	--2505
		x"02",	--2506
		x"0d",	--2507
		x"b8",	--2508
		x"3e",	--2509
		x"40",	--2510
		x"0f",	--2511
		x"b4",	--2512
		x"12",	--2513
		x"0f",	--2514
		x"0e",	--2515
		x"0d",	--2516
		x"3d",	--2517
		x"80",	--2518
		x"b2",	--2519
		x"7d",	--2520
		x"0e",	--2521
		x"0f",	--2522
		x"cd",	--2523
		x"0e",	--2524
		x"3f",	--2525
		x"10",	--2526
		x"3e",	--2527
		x"3f",	--2528
		x"7f",	--2529
		x"7d",	--2530
		x"c5",	--2531
		x"37",	--2532
		x"82",	--2533
		x"07",	--2534
		x"37",	--2535
		x"1a",	--2536
		x"4f",	--2537
		x"0c",	--2538
		x"0d",	--2539
		x"4b",	--2540
		x"7b",	--2541
		x"1f",	--2542
		x"05",	--2543
		x"12",	--2544
		x"0d",	--2545
		x"0c",	--2546
		x"7b",	--2547
		x"fb",	--2548
		x"18",	--2549
		x"09",	--2550
		x"77",	--2551
		x"1f",	--2552
		x"04",	--2553
		x"08",	--2554
		x"09",	--2555
		x"77",	--2556
		x"fc",	--2557
		x"38",	--2558
		x"39",	--2559
		x"08",	--2560
		x"09",	--2561
		x"1e",	--2562
		x"0f",	--2563
		x"08",	--2564
		x"04",	--2565
		x"09",	--2566
		x"02",	--2567
		x"0e",	--2568
		x"0f",	--2569
		x"08",	--2570
		x"09",	--2571
		x"08",	--2572
		x"09",	--2573
		x"0e",	--2574
		x"0f",	--2575
		x"3e",	--2576
		x"7f",	--2577
		x"0f",	--2578
		x"3e",	--2579
		x"40",	--2580
		x"26",	--2581
		x"38",	--2582
		x"3f",	--2583
		x"09",	--2584
		x"0e",	--2585
		x"0f",	--2586
		x"12",	--2587
		x"0f",	--2588
		x"0e",	--2589
		x"12",	--2590
		x"0f",	--2591
		x"0e",	--2592
		x"12",	--2593
		x"0f",	--2594
		x"0e",	--2595
		x"12",	--2596
		x"0f",	--2597
		x"0e",	--2598
		x"12",	--2599
		x"0f",	--2600
		x"0e",	--2601
		x"12",	--2602
		x"0f",	--2603
		x"0e",	--2604
		x"12",	--2605
		x"0f",	--2606
		x"0e",	--2607
		x"3e",	--2608
		x"3f",	--2609
		x"7f",	--2610
		x"5d",	--2611
		x"39",	--2612
		x"00",	--2613
		x"72",	--2614
		x"4d",	--2615
		x"70",	--2616
		x"08",	--2617
		x"09",	--2618
		x"da",	--2619
		x"0f",	--2620
		x"d8",	--2621
		x"0e",	--2622
		x"0f",	--2623
		x"3e",	--2624
		x"80",	--2625
		x"0f",	--2626
		x"0e",	--2627
		x"04",	--2628
		x"38",	--2629
		x"40",	--2630
		x"09",	--2631
		x"d0",	--2632
		x"0f",	--2633
		x"ce",	--2634
		x"f9",	--2635
		x"0b",	--2636
		x"0a",	--2637
		x"2a",	--2638
		x"5b",	--2639
		x"02",	--2640
		x"3b",	--2641
		x"7f",	--2642
		x"1d",	--2643
		x"02",	--2644
		x"12",	--2645
		x"0d",	--2646
		x"12",	--2647
		x"0d",	--2648
		x"12",	--2649
		x"0d",	--2650
		x"12",	--2651
		x"0d",	--2652
		x"12",	--2653
		x"0d",	--2654
		x"12",	--2655
		x"0d",	--2656
		x"12",	--2657
		x"0d",	--2658
		x"4d",	--2659
		x"5f",	--2660
		x"03",	--2661
		x"3f",	--2662
		x"80",	--2663
		x"0f",	--2664
		x"0f",	--2665
		x"ce",	--2666
		x"01",	--2667
		x"0d",	--2668
		x"2d",	--2669
		x"0a",	--2670
		x"51",	--2671
		x"be",	--2672
		x"82",	--2673
		x"02",	--2674
		x"0c",	--2675
		x"0d",	--2676
		x"0c",	--2677
		x"0d",	--2678
		x"0c",	--2679
		x"0d",	--2680
		x"0c",	--2681
		x"0d",	--2682
		x"0c",	--2683
		x"0d",	--2684
		x"0c",	--2685
		x"0d",	--2686
		x"0c",	--2687
		x"0d",	--2688
		x"0c",	--2689
		x"0d",	--2690
		x"fe",	--2691
		x"03",	--2692
		x"00",	--2693
		x"3d",	--2694
		x"00",	--2695
		x"0b",	--2696
		x"3f",	--2697
		x"81",	--2698
		x"0c",	--2699
		x"0d",	--2700
		x"0a",	--2701
		x"3f",	--2702
		x"3d",	--2703
		x"00",	--2704
		x"f9",	--2705
		x"8e",	--2706
		x"02",	--2707
		x"8e",	--2708
		x"04",	--2709
		x"8e",	--2710
		x"06",	--2711
		x"3a",	--2712
		x"3b",	--2713
		x"30",	--2714
		x"3d",	--2715
		x"ff",	--2716
		x"2a",	--2717
		x"3d",	--2718
		x"81",	--2719
		x"8e",	--2720
		x"02",	--2721
		x"fe",	--2722
		x"03",	--2723
		x"00",	--2724
		x"0c",	--2725
		x"0d",	--2726
		x"0c",	--2727
		x"0d",	--2728
		x"0c",	--2729
		x"0d",	--2730
		x"0c",	--2731
		x"0d",	--2732
		x"0c",	--2733
		x"0d",	--2734
		x"0c",	--2735
		x"0d",	--2736
		x"0c",	--2737
		x"0d",	--2738
		x"0c",	--2739
		x"0d",	--2740
		x"0a",	--2741
		x"0b",	--2742
		x"0a",	--2743
		x"3b",	--2744
		x"00",	--2745
		x"8e",	--2746
		x"04",	--2747
		x"8e",	--2748
		x"06",	--2749
		x"3a",	--2750
		x"3b",	--2751
		x"30",	--2752
		x"0b",	--2753
		x"ad",	--2754
		x"ee",	--2755
		x"00",	--2756
		x"3a",	--2757
		x"3b",	--2758
		x"30",	--2759
		x"0a",	--2760
		x"0c",	--2761
		x"0c",	--2762
		x"0d",	--2763
		x"0c",	--2764
		x"3d",	--2765
		x"10",	--2766
		x"0c",	--2767
		x"02",	--2768
		x"0d",	--2769
		x"08",	--2770
		x"de",	--2771
		x"00",	--2772
		x"e4",	--2773
		x"0b",	--2774
		x"f2",	--2775
		x"ee",	--2776
		x"00",	--2777
		x"e3",	--2778
		x"ce",	--2779
		x"00",	--2780
		x"dc",	--2781
		x"0b",	--2782
		x"6d",	--2783
		x"6d",	--2784
		x"12",	--2785
		x"6c",	--2786
		x"6c",	--2787
		x"0f",	--2788
		x"6d",	--2789
		x"41",	--2790
		x"6c",	--2791
		x"11",	--2792
		x"6d",	--2793
		x"0d",	--2794
		x"6c",	--2795
		x"14",	--2796
		x"5d",	--2797
		x"01",	--2798
		x"5d",	--2799
		x"01",	--2800
		x"14",	--2801
		x"4d",	--2802
		x"09",	--2803
		x"1e",	--2804
		x"0f",	--2805
		x"3b",	--2806
		x"30",	--2807
		x"6c",	--2808
		x"28",	--2809
		x"ce",	--2810
		x"01",	--2811
		x"f7",	--2812
		x"3e",	--2813
		x"0f",	--2814
		x"3b",	--2815
		x"30",	--2816
		x"cf",	--2817
		x"01",	--2818
		x"f0",	--2819
		x"3e",	--2820
		x"f8",	--2821
		x"1b",	--2822
		x"02",	--2823
		x"1c",	--2824
		x"02",	--2825
		x"0c",	--2826
		x"e6",	--2827
		x"0b",	--2828
		x"16",	--2829
		x"1b",	--2830
		x"04",	--2831
		x"1f",	--2832
		x"06",	--2833
		x"1c",	--2834
		x"04",	--2835
		x"1e",	--2836
		x"06",	--2837
		x"0e",	--2838
		x"da",	--2839
		x"0f",	--2840
		x"02",	--2841
		x"0c",	--2842
		x"d6",	--2843
		x"0f",	--2844
		x"06",	--2845
		x"0e",	--2846
		x"02",	--2847
		x"0b",	--2848
		x"02",	--2849
		x"0e",	--2850
		x"d1",	--2851
		x"4d",	--2852
		x"ce",	--2853
		x"3e",	--2854
		x"d6",	--2855
		x"6c",	--2856
		x"d7",	--2857
		x"5e",	--2858
		x"01",	--2859
		x"5f",	--2860
		x"01",	--2861
		x"0e",	--2862
		x"c5",	--2863
		x"0d",	--2864
		x"0f",	--2865
		x"04",	--2866
		x"3d",	--2867
		x"03",	--2868
		x"3f",	--2869
		x"1f",	--2870
		x"0e",	--2871
		x"03",	--2872
		x"5d",	--2873
		x"3e",	--2874
		x"1e",	--2875
		x"0d",	--2876
		x"b0",	--2877
		x"e6",	--2878
		x"3d",	--2879
		x"6d",	--2880
		x"02",	--2881
		x"3e",	--2882
		x"1e",	--2883
		x"5d",	--2884
		x"02",	--2885
		x"3f",	--2886
		x"1f",	--2887
		x"30",	--2888
		x"b0",	--2889
		x"60",	--2890
		x"0f",	--2891
		x"30",	--2892
		x"0b",	--2893
		x"0b",	--2894
		x"0f",	--2895
		x"06",	--2896
		x"3b",	--2897
		x"03",	--2898
		x"3e",	--2899
		x"3f",	--2900
		x"1e",	--2901
		x"0f",	--2902
		x"0d",	--2903
		x"05",	--2904
		x"5b",	--2905
		x"3c",	--2906
		x"3d",	--2907
		x"1c",	--2908
		x"0d",	--2909
		x"b0",	--2910
		x"08",	--2911
		x"6b",	--2912
		x"04",	--2913
		x"3c",	--2914
		x"3d",	--2915
		x"1c",	--2916
		x"0d",	--2917
		x"5b",	--2918
		x"04",	--2919
		x"3e",	--2920
		x"3f",	--2921
		x"1e",	--2922
		x"0f",	--2923
		x"3b",	--2924
		x"30",	--2925
		x"b0",	--2926
		x"9a",	--2927
		x"0e",	--2928
		x"0f",	--2929
		x"30",	--2930
		x"7c",	--2931
		x"10",	--2932
		x"0d",	--2933
		x"0e",	--2934
		x"0f",	--2935
		x"0e",	--2936
		x"0e",	--2937
		x"02",	--2938
		x"0e",	--2939
		x"1f",	--2940
		x"1c",	--2941
		x"f8",	--2942
		x"30",	--2943
		x"b0",	--2944
		x"e6",	--2945
		x"0f",	--2946
		x"30",	--2947
		x"0b",	--2948
		x"0a",	--2949
		x"09",	--2950
		x"79",	--2951
		x"20",	--2952
		x"0a",	--2953
		x"0b",	--2954
		x"0c",	--2955
		x"0d",	--2956
		x"0e",	--2957
		x"0f",	--2958
		x"0c",	--2959
		x"0d",	--2960
		x"0d",	--2961
		x"06",	--2962
		x"02",	--2963
		x"0c",	--2964
		x"03",	--2965
		x"0c",	--2966
		x"0d",	--2967
		x"1e",	--2968
		x"19",	--2969
		x"f2",	--2970
		x"39",	--2971
		x"3a",	--2972
		x"3b",	--2973
		x"30",	--2974
		x"b0",	--2975
		x"08",	--2976
		x"0e",	--2977
		x"0f",	--2978
		x"30",	--2979
		x"00",	--2980
		x"32",	--2981
		x"f0",	--2982
		x"fd",	--2983
		x"63",	--2984
		x"72",	--2985
		x"65",	--2986
		x"74",	--2987
		x"75",	--2988
		x"61",	--2989
		x"65",	--2990
		x"0d",	--2991
		x"00",	--2992
		x"25",	--2993
		x"20",	--2994
		x"45",	--2995
		x"54",	--2996
		x"52",	--2997
		x"47",	--2998
		x"54",	--2999
		x"0a",	--3000
		x"53",	--3001
		x"6d",	--3002
		x"74",	--3003
		x"69",	--3004
		x"67",	--3005
		x"77",	--3006
		x"6e",	--3007
		x"20",	--3008
		x"65",	--3009
		x"72",	--3010
		x"62",	--3011
		x"79",	--3012
		x"77",	--3013
		x"6f",	--3014
		x"67",	--3015
		x"0a",	--3016
		x"0d",	--3017
		x"3d",	--3018
		x"3d",	--3019
		x"3d",	--3020
		x"20",	--3021
		x"70",	--3022
		x"6e",	--3023
		x"53",	--3024
		x"34",	--3025
		x"30",	--3026
		x"69",	--3027
		x"20",	--3028
		x"63",	--3029
		x"69",	--3030
		x"6e",	--3031
		x"3d",	--3032
		x"3d",	--3033
		x"3d",	--3034
		x"0d",	--3035
		x"00",	--3036
		x"0a",	--3037
		x"69",	--3038
		x"70",	--3039
		x"65",	--3040
		x"4c",	--3041
		x"6e",	--3042
		x"20",	--3043
		x"64",	--3044
		x"74",	--3045
		x"72",	--3046
		x"52",	--3047
		x"61",	--3048
		x"79",	--3049
		x"0a",	--3050
		x"0d",	--3051
		x"42",	--3052
		x"55",	--3053
		x"3d",	--3054
		x"64",	--3055
		x"0a",	--3056
		x"0d",	--3057
		x"74",	--3058
		x"73",	--3059
		x"3d",	--3060
		x"63",	--3061
		x"0a",	--3062
		x"3e",	--3063
		x"00",	--3064
		x"0a",	--3065
		x"3a",	--3066
		x"73",	--3067
		x"0a",	--3068
		x"08",	--3069
		x"08",	--3070
		x"25",	--3071
		x"00",	--3072
		x"72",	--3073
		x"74",	--3074
		x"0a",	--3075
		x"00",	--3076
		x"6f",	--3077
		x"72",	--3078
		x"63",	--3079
		x"20",	--3080
		x"73",	--3081
		x"67",	--3082
		x"3a",	--3083
		x"0a",	--3084
		x"09",	--3085
		x"63",	--3086
		x"52",	--3087
		x"47",	--3088
		x"53",	--3089
		x"45",	--3090
		x"20",	--3091
		x"41",	--3092
		x"55",	--3093
		x"0d",	--3094
		x"00",	--3095
		x"6f",	--3096
		x"65",	--3097
		x"68",	--3098
		x"6e",	--3099
		x"20",	--3100
		x"65",	--3101
		x"74",	--3102
		x"74",	--3103
		x"72",	--3104
		x"69",	--3105
		x"6c",	--3106
		x"20",	--3107
		x"72",	--3108
		x"6e",	--3109
		x"0d",	--3110
		x"00",	--3111
		x"3d",	--3112
		x"64",	--3113
		x"76",	--3114
		x"25",	--3115
		x"0d",	--3116
		x"00",	--3117
		x"65",	--3118
		x"64",	--3119
		x"0d",	--3120
		x"09",	--3121
		x"63",	--3122
		x"52",	--3123
		x"47",	--3124
		x"53",	--3125
		x"45",	--3126
		x"0d",	--3127
		x"00",	--3128
		x"63",	--3129
		x"69",	--3130
		x"20",	--3131
		x"6f",	--3132
		x"20",	--3133
		x"20",	--3134
		x"75",	--3135
		x"62",	--3136
		x"72",	--3137
		x"0a",	--3138
		x"25",	--3139
		x"3a",	--3140
		x"6e",	--3141
		x"20",	--3142
		x"75",	--3143
		x"68",	--3144
		x"63",	--3145
		x"6d",	--3146
		x"61",	--3147
		x"64",	--3148
		x"0a",	--3149
		x"ea",	--3150
		x"18",	--3151
		x"18",	--3152
		x"18",	--3153
		x"18",	--3154
		x"18",	--3155
		x"18",	--3156
		x"18",	--3157
		x"18",	--3158
		x"18",	--3159
		x"18",	--3160
		x"18",	--3161
		x"18",	--3162
		x"18",	--3163
		x"18",	--3164
		x"18",	--3165
		x"18",	--3166
		x"18",	--3167
		x"18",	--3168
		x"18",	--3169
		x"18",	--3170
		x"18",	--3171
		x"18",	--3172
		x"18",	--3173
		x"18",	--3174
		x"18",	--3175
		x"18",	--3176
		x"18",	--3177
		x"18",	--3178
		x"dc",	--3179
		x"18",	--3180
		x"18",	--3181
		x"18",	--3182
		x"18",	--3183
		x"18",	--3184
		x"18",	--3185
		x"18",	--3186
		x"18",	--3187
		x"18",	--3188
		x"18",	--3189
		x"18",	--3190
		x"18",	--3191
		x"18",	--3192
		x"18",	--3193
		x"18",	--3194
		x"18",	--3195
		x"18",	--3196
		x"18",	--3197
		x"18",	--3198
		x"18",	--3199
		x"18",	--3200
		x"18",	--3201
		x"18",	--3202
		x"18",	--3203
		x"18",	--3204
		x"18",	--3205
		x"18",	--3206
		x"18",	--3207
		x"18",	--3208
		x"18",	--3209
		x"18",	--3210
		x"ce",	--3211
		x"c0",	--3212
		x"b2",	--3213
		x"18",	--3214
		x"18",	--3215
		x"18",	--3216
		x"18",	--3217
		x"18",	--3218
		x"18",	--3219
		x"18",	--3220
		x"9a",	--3221
		x"18",	--3222
		x"88",	--3223
		x"18",	--3224
		x"18",	--3225
		x"18",	--3226
		x"18",	--3227
		x"6c",	--3228
		x"18",	--3229
		x"18",	--3230
		x"18",	--3231
		x"5e",	--3232
		x"4c",	--3233
		x"30",	--3234
		x"32",	--3235
		x"34",	--3236
		x"36",	--3237
		x"38",	--3238
		x"61",	--3239
		x"63",	--3240
		x"65",	--3241
		x"00",	--3242
		x"00",	--3243
		x"00",	--3244
		x"00",	--3245
		x"00",	--3246
		x"00",	--3247
		x"02",	--3248
		x"03",	--3249
		x"03",	--3250
		x"04",	--3251
		x"04",	--3252
		x"04",	--3253
		x"04",	--3254
		x"05",	--3255
		x"05",	--3256
		x"05",	--3257
		x"05",	--3258
		x"05",	--3259
		x"05",	--3260
		x"05",	--3261
		x"05",	--3262
		x"06",	--3263
		x"06",	--3264
		x"06",	--3265
		x"06",	--3266
		x"06",	--3267
		x"06",	--3268
		x"06",	--3269
		x"06",	--3270
		x"06",	--3271
		x"06",	--3272
		x"06",	--3273
		x"06",	--3274
		x"06",	--3275
		x"06",	--3276
		x"06",	--3277
		x"06",	--3278
		x"07",	--3279
		x"07",	--3280
		x"07",	--3281
		x"07",	--3282
		x"07",	--3283
		x"07",	--3284
		x"07",	--3285
		x"07",	--3286
		x"07",	--3287
		x"07",	--3288
		x"07",	--3289
		x"07",	--3290
		x"07",	--3291
		x"07",	--3292
		x"07",	--3293
		x"07",	--3294
		x"07",	--3295
		x"07",	--3296
		x"07",	--3297
		x"07",	--3298
		x"07",	--3299
		x"07",	--3300
		x"07",	--3301
		x"07",	--3302
		x"07",	--3303
		x"07",	--3304
		x"07",	--3305
		x"07",	--3306
		x"07",	--3307
		x"07",	--3308
		x"07",	--3309
		x"07",	--3310
		x"08",	--3311
		x"08",	--3312
		x"08",	--3313
		x"08",	--3314
		x"08",	--3315
		x"08",	--3316
		x"08",	--3317
		x"08",	--3318
		x"08",	--3319
		x"08",	--3320
		x"08",	--3321
		x"08",	--3322
		x"08",	--3323
		x"08",	--3324
		x"08",	--3325
		x"08",	--3326
		x"08",	--3327
		x"08",	--3328
		x"08",	--3329
		x"08",	--3330
		x"08",	--3331
		x"08",	--3332
		x"08",	--3333
		x"08",	--3334
		x"08",	--3335
		x"08",	--3336
		x"08",	--3337
		x"08",	--3338
		x"08",	--3339
		x"08",	--3340
		x"08",	--3341
		x"08",	--3342
		x"08",	--3343
		x"08",	--3344
		x"08",	--3345
		x"08",	--3346
		x"08",	--3347
		x"08",	--3348
		x"08",	--3349
		x"08",	--3350
		x"08",	--3351
		x"08",	--3352
		x"08",	--3353
		x"08",	--3354
		x"08",	--3355
		x"08",	--3356
		x"08",	--3357
		x"08",	--3358
		x"08",	--3359
		x"08",	--3360
		x"08",	--3361
		x"08",	--3362
		x"08",	--3363
		x"08",	--3364
		x"08",	--3365
		x"08",	--3366
		x"08",	--3367
		x"08",	--3368
		x"08",	--3369
		x"08",	--3370
		x"08",	--3371
		x"08",	--3372
		x"08",	--3373
		x"08",	--3374
		x"ff",	--3375
		x"ff",	--3376
		x"ff",	--3377
		x"ff",	--3378
		x"ff",	--3379
		x"ff",	--3380
		x"ff",	--3381
		x"ff",	--3382
		x"ff",	--3383
		x"ff",	--3384
		x"ff",	--3385
		x"ff",	--3386
		x"ff",	--3387
		x"ff",	--3388
		x"ff",	--3389
		x"ff",	--3390
		x"ff",	--3391
		x"ff",	--3392
		x"ff",	--3393
		x"ff",	--3394
		x"ff",	--3395
		x"ff",	--3396
		x"ff",	--3397
		x"ff",	--3398
		x"ff",	--3399
		x"ff",	--3400
		x"ff",	--3401
		x"ff",	--3402
		x"ff",	--3403
		x"ff",	--3404
		x"ff",	--3405
		x"ff",	--3406
		x"ff",	--3407
		x"ff",	--3408
		x"ff",	--3409
		x"ff",	--3410
		x"ff",	--3411
		x"ff",	--3412
		x"ff",	--3413
		x"ff",	--3414
		x"ff",	--3415
		x"ff",	--3416
		x"ff",	--3417
		x"ff",	--3418
		x"ff",	--3419
		x"ff",	--3420
		x"ff",	--3421
		x"ff",	--3422
		x"ff",	--3423
		x"ff",	--3424
		x"ff",	--3425
		x"ff",	--3426
		x"ff",	--3427
		x"ff",	--3428
		x"ff",	--3429
		x"ff",	--3430
		x"ff",	--3431
		x"ff",	--3432
		x"ff",	--3433
		x"ff",	--3434
		x"ff",	--3435
		x"ff",	--3436
		x"ff",	--3437
		x"ff",	--3438
		x"ff",	--3439
		x"ff",	--3440
		x"ff",	--3441
		x"ff",	--3442
		x"ff",	--3443
		x"ff",	--3444
		x"ff",	--3445
		x"ff",	--3446
		x"ff",	--3447
		x"ff",	--3448
		x"ff",	--3449
		x"ff",	--3450
		x"ff",	--3451
		x"ff",	--3452
		x"ff",	--3453
		x"ff",	--3454
		x"ff",	--3455
		x"ff",	--3456
		x"ff",	--3457
		x"ff",	--3458
		x"ff",	--3459
		x"ff",	--3460
		x"ff",	--3461
		x"ff",	--3462
		x"ff",	--3463
		x"ff",	--3464
		x"ff",	--3465
		x"ff",	--3466
		x"ff",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"be",	--4080
		x"be",	--4081
		x"be",	--4082
		x"be",	--4083
		x"be",	--4084
		x"be",	--4085
		x"be",	--4086
		x"f4",	--4087
		x"be",	--4088
		x"be",	--4089
		x"be",	--4090
		x"be",	--4091
		x"be",	--4092
		x"be",	--4093
		x"be",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"03",	--5
		x"40",	--6
		x"06",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"03",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fa",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"01",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"03",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"43",	--40
		x"00",	--41
		x"40",	--42
		x"c2",	--43
		x"43",	--44
		x"12",	--45
		x"e9",	--46
		x"12",	--47
		x"e5",	--48
		x"43",	--49
		x"00",	--50
		x"12",	--51
		x"f7",	--52
		x"12",	--53
		x"e7",	--54
		x"40",	--55
		x"f7",	--56
		x"00",	--57
		x"12",	--58
		x"e7",	--59
		x"53",	--60
		x"12",	--61
		x"12",	--62
		x"00",	--63
		x"12",	--64
		x"f7",	--65
		x"12",	--66
		x"e7",	--67
		x"50",	--68
		x"00",	--69
		x"12",	--70
		x"00",	--71
		x"12",	--72
		x"f7",	--73
		x"12",	--74
		x"e7",	--75
		x"52",	--76
		x"40",	--77
		x"e2",	--78
		x"40",	--79
		x"00",	--80
		x"12",	--81
		x"e5",	--82
		x"40",	--83
		x"e3",	--84
		x"40",	--85
		x"00",	--86
		x"12",	--87
		x"e5",	--88
		x"40",	--89
		x"e1",	--90
		x"40",	--91
		x"00",	--92
		x"12",	--93
		x"e5",	--94
		x"43",	--95
		x"40",	--96
		x"4e",	--97
		x"40",	--98
		x"01",	--99
		x"41",	--100
		x"50",	--101
		x"00",	--102
		x"12",	--103
		x"e4",	--104
		x"41",	--105
		x"50",	--106
		x"00",	--107
		x"12",	--108
		x"e4",	--109
		x"43",	--110
		x"40",	--111
		x"4e",	--112
		x"40",	--113
		x"01",	--114
		x"41",	--115
		x"12",	--116
		x"e4",	--117
		x"41",	--118
		x"12",	--119
		x"e4",	--120
		x"41",	--121
		x"41",	--122
		x"50",	--123
		x"00",	--124
		x"12",	--125
		x"e1",	--126
		x"d2",	--127
		x"43",	--128
		x"12",	--129
		x"f7",	--130
		x"12",	--131
		x"e7",	--132
		x"53",	--133
		x"43",	--134
		x"d0",	--135
		x"00",	--136
		x"53",	--137
		x"90",	--138
		x"00",	--139
		x"24",	--140
		x"43",	--141
		x"4b",	--142
		x"f0",	--143
		x"00",	--144
		x"24",	--145
		x"5f",	--146
		x"53",	--147
		x"23",	--148
		x"4f",	--149
		x"3c",	--150
		x"43",	--151
		x"43",	--152
		x"4f",	--153
		x"00",	--154
		x"12",	--155
		x"e9",	--156
		x"93",	--157
		x"27",	--158
		x"12",	--159
		x"e9",	--160
		x"92",	--161
		x"24",	--162
		x"90",	--163
		x"00",	--164
		x"20",	--165
		x"12",	--166
		x"f7",	--167
		x"12",	--168
		x"e7",	--169
		x"53",	--170
		x"40",	--171
		x"00",	--172
		x"51",	--173
		x"5f",	--174
		x"43",	--175
		x"00",	--176
		x"12",	--177
		x"12",	--178
		x"f7",	--179
		x"12",	--180
		x"e7",	--181
		x"52",	--182
		x"41",	--183
		x"50",	--184
		x"00",	--185
		x"41",	--186
		x"00",	--187
		x"12",	--188
		x"e5",	--189
		x"3f",	--190
		x"93",	--191
		x"27",	--192
		x"53",	--193
		x"12",	--194
		x"f7",	--195
		x"12",	--196
		x"e7",	--197
		x"53",	--198
		x"3f",	--199
		x"90",	--200
		x"00",	--201
		x"2f",	--202
		x"4f",	--203
		x"11",	--204
		x"12",	--205
		x"12",	--206
		x"f7",	--207
		x"4f",	--208
		x"00",	--209
		x"12",	--210
		x"e7",	--211
		x"52",	--212
		x"40",	--213
		x"00",	--214
		x"51",	--215
		x"5a",	--216
		x"41",	--217
		x"00",	--218
		x"4f",	--219
		x"00",	--220
		x"53",	--221
		x"3f",	--222
		x"40",	--223
		x"f7",	--224
		x"4f",	--225
		x"02",	--226
		x"4e",	--227
		x"02",	--228
		x"41",	--229
		x"82",	--230
		x"90",	--231
		x"00",	--232
		x"00",	--233
		x"20",	--234
		x"93",	--235
		x"00",	--236
		x"24",	--237
		x"41",	--238
		x"4f",	--239
		x"53",	--240
		x"41",	--241
		x"52",	--242
		x"12",	--243
		x"e3",	--244
		x"93",	--245
		x"00",	--246
		x"24",	--247
		x"41",	--248
		x"4f",	--249
		x"41",	--250
		x"53",	--251
		x"12",	--252
		x"e3",	--253
		x"93",	--254
		x"00",	--255
		x"24",	--256
		x"41",	--257
		x"00",	--258
		x"43",	--259
		x"12",	--260
		x"f1",	--261
		x"43",	--262
		x"40",	--263
		x"42",	--264
		x"12",	--265
		x"ef",	--266
		x"4e",	--267
		x"4f",	--268
		x"42",	--269
		x"02",	--270
		x"12",	--271
		x"e5",	--272
		x"41",	--273
		x"00",	--274
		x"43",	--275
		x"12",	--276
		x"f1",	--277
		x"43",	--278
		x"40",	--279
		x"42",	--280
		x"12",	--281
		x"ef",	--282
		x"4e",	--283
		x"4f",	--284
		x"42",	--285
		x"02",	--286
		x"12",	--287
		x"e5",	--288
		x"43",	--289
		x"52",	--290
		x"41",	--291
		x"12",	--292
		x"f7",	--293
		x"4f",	--294
		x"00",	--295
		x"12",	--296
		x"e7",	--297
		x"41",	--298
		x"00",	--299
		x"4f",	--300
		x"11",	--301
		x"4f",	--302
		x"00",	--303
		x"12",	--304
		x"f7",	--305
		x"12",	--306
		x"e7",	--307
		x"52",	--308
		x"43",	--309
		x"52",	--310
		x"41",	--311
		x"12",	--312
		x"f7",	--313
		x"12",	--314
		x"e7",	--315
		x"53",	--316
		x"43",	--317
		x"3f",	--318
		x"12",	--319
		x"50",	--320
		x"ff",	--321
		x"4f",	--322
		x"12",	--323
		x"f8",	--324
		x"12",	--325
		x"e7",	--326
		x"53",	--327
		x"90",	--328
		x"00",	--329
		x"00",	--330
		x"20",	--331
		x"93",	--332
		x"00",	--333
		x"24",	--334
		x"41",	--335
		x"4b",	--336
		x"53",	--337
		x"41",	--338
		x"52",	--339
		x"12",	--340
		x"e3",	--341
		x"93",	--342
		x"00",	--343
		x"24",	--344
		x"41",	--345
		x"4f",	--346
		x"41",	--347
		x"53",	--348
		x"12",	--349
		x"e3",	--350
		x"93",	--351
		x"00",	--352
		x"24",	--353
		x"12",	--354
		x"00",	--355
		x"12",	--356
		x"00",	--357
		x"12",	--358
		x"f8",	--359
		x"12",	--360
		x"e7",	--361
		x"50",	--362
		x"00",	--363
		x"41",	--364
		x"00",	--365
		x"41",	--366
		x"00",	--367
		x"00",	--368
		x"43",	--369
		x"50",	--370
		x"00",	--371
		x"41",	--372
		x"41",	--373
		x"12",	--374
		x"f8",	--375
		x"12",	--376
		x"e7",	--377
		x"4b",	--378
		x"11",	--379
		x"4f",	--380
		x"00",	--381
		x"12",	--382
		x"f8",	--383
		x"12",	--384
		x"e7",	--385
		x"52",	--386
		x"43",	--387
		x"50",	--388
		x"00",	--389
		x"41",	--390
		x"41",	--391
		x"12",	--392
		x"f8",	--393
		x"12",	--394
		x"e7",	--395
		x"53",	--396
		x"43",	--397
		x"3f",	--398
		x"12",	--399
		x"82",	--400
		x"4f",	--401
		x"12",	--402
		x"f8",	--403
		x"12",	--404
		x"e7",	--405
		x"53",	--406
		x"90",	--407
		x"00",	--408
		x"00",	--409
		x"20",	--410
		x"93",	--411
		x"00",	--412
		x"24",	--413
		x"41",	--414
		x"4b",	--415
		x"53",	--416
		x"41",	--417
		x"53",	--418
		x"12",	--419
		x"e3",	--420
		x"93",	--421
		x"00",	--422
		x"24",	--423
		x"41",	--424
		x"00",	--425
		x"12",	--426
		x"12",	--427
		x"12",	--428
		x"f8",	--429
		x"12",	--430
		x"e7",	--431
		x"50",	--432
		x"00",	--433
		x"43",	--434
		x"52",	--435
		x"41",	--436
		x"41",	--437
		x"12",	--438
		x"f8",	--439
		x"12",	--440
		x"e7",	--441
		x"4b",	--442
		x"11",	--443
		x"4f",	--444
		x"00",	--445
		x"12",	--446
		x"f8",	--447
		x"12",	--448
		x"e7",	--449
		x"52",	--450
		x"43",	--451
		x"52",	--452
		x"41",	--453
		x"41",	--454
		x"12",	--455
		x"f8",	--456
		x"12",	--457
		x"e7",	--458
		x"53",	--459
		x"43",	--460
		x"3f",	--461
		x"12",	--462
		x"12",	--463
		x"12",	--464
		x"12",	--465
		x"12",	--466
		x"43",	--467
		x"00",	--468
		x"43",	--469
		x"00",	--470
		x"4e",	--471
		x"93",	--472
		x"24",	--473
		x"4e",	--474
		x"53",	--475
		x"4e",	--476
		x"43",	--477
		x"43",	--478
		x"43",	--479
		x"3c",	--480
		x"90",	--481
		x"00",	--482
		x"2c",	--483
		x"4f",	--484
		x"5c",	--485
		x"5c",	--486
		x"5c",	--487
		x"5c",	--488
		x"4c",	--489
		x"00",	--490
		x"50",	--491
		x"ff",	--492
		x"48",	--493
		x"11",	--494
		x"5a",	--495
		x"4c",	--496
		x"00",	--497
		x"43",	--498
		x"53",	--499
		x"49",	--500
		x"4b",	--501
		x"4b",	--502
		x"93",	--503
		x"24",	--504
		x"90",	--505
		x"00",	--506
		x"24",	--507
		x"90",	--508
		x"00",	--509
		x"24",	--510
		x"4c",	--511
		x"50",	--512
		x"ff",	--513
		x"93",	--514
		x"23",	--515
		x"90",	--516
		x"00",	--517
		x"2c",	--518
		x"4f",	--519
		x"5a",	--520
		x"4a",	--521
		x"5c",	--522
		x"5c",	--523
		x"5a",	--524
		x"4c",	--525
		x"00",	--526
		x"50",	--527
		x"ff",	--528
		x"48",	--529
		x"11",	--530
		x"58",	--531
		x"4c",	--532
		x"00",	--533
		x"3f",	--534
		x"43",	--535
		x"3f",	--536
		x"4c",	--537
		x"50",	--538
		x"ff",	--539
		x"90",	--540
		x"00",	--541
		x"2c",	--542
		x"4f",	--543
		x"5c",	--544
		x"5c",	--545
		x"5c",	--546
		x"5c",	--547
		x"4c",	--548
		x"00",	--549
		x"50",	--550
		x"ff",	--551
		x"3f",	--552
		x"4c",	--553
		x"50",	--554
		x"ff",	--555
		x"90",	--556
		x"00",	--557
		x"2c",	--558
		x"4f",	--559
		x"5c",	--560
		x"5c",	--561
		x"5c",	--562
		x"5c",	--563
		x"4c",	--564
		x"00",	--565
		x"50",	--566
		x"ff",	--567
		x"3f",	--568
		x"43",	--569
		x"00",	--570
		x"43",	--571
		x"41",	--572
		x"41",	--573
		x"41",	--574
		x"41",	--575
		x"41",	--576
		x"41",	--577
		x"43",	--578
		x"00",	--579
		x"4a",	--580
		x"53",	--581
		x"5e",	--582
		x"41",	--583
		x"41",	--584
		x"41",	--585
		x"41",	--586
		x"41",	--587
		x"41",	--588
		x"11",	--589
		x"12",	--590
		x"12",	--591
		x"f8",	--592
		x"12",	--593
		x"e7",	--594
		x"52",	--595
		x"43",	--596
		x"41",	--597
		x"41",	--598
		x"41",	--599
		x"41",	--600
		x"41",	--601
		x"41",	--602
		x"12",	--603
		x"12",	--604
		x"4e",	--605
		x"4c",	--606
		x"4e",	--607
		x"00",	--608
		x"4d",	--609
		x"00",	--610
		x"4c",	--611
		x"00",	--612
		x"4d",	--613
		x"43",	--614
		x"40",	--615
		x"36",	--616
		x"40",	--617
		x"01",	--618
		x"12",	--619
		x"f6",	--620
		x"4e",	--621
		x"00",	--622
		x"12",	--623
		x"c2",	--624
		x"43",	--625
		x"4a",	--626
		x"01",	--627
		x"40",	--628
		x"00",	--629
		x"01",	--630
		x"42",	--631
		x"01",	--632
		x"00",	--633
		x"41",	--634
		x"43",	--635
		x"41",	--636
		x"41",	--637
		x"41",	--638
		x"12",	--639
		x"12",	--640
		x"12",	--641
		x"43",	--642
		x"00",	--643
		x"40",	--644
		x"3f",	--645
		x"00",	--646
		x"4f",	--647
		x"4b",	--648
		x"00",	--649
		x"43",	--650
		x"12",	--651
		x"f1",	--652
		x"43",	--653
		x"40",	--654
		x"3f",	--655
		x"12",	--656
		x"ed",	--657
		x"4e",	--658
		x"4f",	--659
		x"4b",	--660
		x"00",	--661
		x"43",	--662
		x"12",	--663
		x"f1",	--664
		x"4e",	--665
		x"4f",	--666
		x"48",	--667
		x"49",	--668
		x"12",	--669
		x"ec",	--670
		x"12",	--671
		x"e9",	--672
		x"4e",	--673
		x"00",	--674
		x"43",	--675
		x"00",	--676
		x"41",	--677
		x"41",	--678
		x"41",	--679
		x"41",	--680
		x"12",	--681
		x"12",	--682
		x"12",	--683
		x"4d",	--684
		x"4e",	--685
		x"4d",	--686
		x"00",	--687
		x"4e",	--688
		x"00",	--689
		x"4f",	--690
		x"49",	--691
		x"00",	--692
		x"43",	--693
		x"12",	--694
		x"f1",	--695
		x"4e",	--696
		x"4f",	--697
		x"4a",	--698
		x"4b",	--699
		x"12",	--700
		x"ed",	--701
		x"4e",	--702
		x"4f",	--703
		x"49",	--704
		x"00",	--705
		x"43",	--706
		x"12",	--707
		x"f1",	--708
		x"4e",	--709
		x"4f",	--710
		x"4a",	--711
		x"4b",	--712
		x"12",	--713
		x"ec",	--714
		x"12",	--715
		x"e9",	--716
		x"4e",	--717
		x"00",	--718
		x"41",	--719
		x"41",	--720
		x"41",	--721
		x"41",	--722
		x"41",	--723
		x"42",	--724
		x"02",	--725
		x"90",	--726
		x"00",	--727
		x"34",	--728
		x"4c",	--729
		x"5d",	--730
		x"5d",	--731
		x"50",	--732
		x"02",	--733
		x"4f",	--734
		x"00",	--735
		x"4e",	--736
		x"00",	--737
		x"53",	--738
		x"4c",	--739
		x"02",	--740
		x"43",	--741
		x"41",	--742
		x"43",	--743
		x"41",	--744
		x"12",	--745
		x"42",	--746
		x"02",	--747
		x"93",	--748
		x"38",	--749
		x"92",	--750
		x"02",	--751
		x"24",	--752
		x"40",	--753
		x"02",	--754
		x"43",	--755
		x"3c",	--756
		x"52",	--757
		x"9f",	--758
		x"ff",	--759
		x"24",	--760
		x"53",	--761
		x"9b",	--762
		x"23",	--763
		x"12",	--764
		x"f8",	--765
		x"12",	--766
		x"e7",	--767
		x"53",	--768
		x"43",	--769
		x"41",	--770
		x"41",	--771
		x"43",	--772
		x"5c",	--773
		x"5c",	--774
		x"50",	--775
		x"02",	--776
		x"4e",	--777
		x"12",	--778
		x"00",	--779
		x"41",	--780
		x"41",	--781
		x"42",	--782
		x"00",	--783
		x"f2",	--784
		x"23",	--785
		x"4f",	--786
		x"00",	--787
		x"4f",	--788
		x"00",	--789
		x"43",	--790
		x"41",	--791
		x"f0",	--792
		x"00",	--793
		x"4f",	--794
		x"f9",	--795
		x"11",	--796
		x"12",	--797
		x"e6",	--798
		x"41",	--799
		x"12",	--800
		x"4f",	--801
		x"4f",	--802
		x"11",	--803
		x"11",	--804
		x"11",	--805
		x"11",	--806
		x"4e",	--807
		x"12",	--808
		x"e6",	--809
		x"4b",	--810
		x"12",	--811
		x"e6",	--812
		x"41",	--813
		x"41",	--814
		x"12",	--815
		x"12",	--816
		x"4f",	--817
		x"40",	--818
		x"00",	--819
		x"4a",	--820
		x"4b",	--821
		x"f0",	--822
		x"00",	--823
		x"24",	--824
		x"11",	--825
		x"53",	--826
		x"23",	--827
		x"f3",	--828
		x"24",	--829
		x"40",	--830
		x"00",	--831
		x"12",	--832
		x"e6",	--833
		x"53",	--834
		x"93",	--835
		x"23",	--836
		x"41",	--837
		x"41",	--838
		x"41",	--839
		x"40",	--840
		x"00",	--841
		x"3f",	--842
		x"12",	--843
		x"4f",	--844
		x"4f",	--845
		x"10",	--846
		x"11",	--847
		x"4e",	--848
		x"12",	--849
		x"e6",	--850
		x"4b",	--851
		x"12",	--852
		x"e6",	--853
		x"41",	--854
		x"41",	--855
		x"12",	--856
		x"12",	--857
		x"4e",	--858
		x"4f",	--859
		x"4f",	--860
		x"10",	--861
		x"11",	--862
		x"4d",	--863
		x"12",	--864
		x"e6",	--865
		x"4b",	--866
		x"12",	--867
		x"e6",	--868
		x"4b",	--869
		x"4a",	--870
		x"10",	--871
		x"10",	--872
		x"ec",	--873
		x"ec",	--874
		x"4d",	--875
		x"12",	--876
		x"e6",	--877
		x"4a",	--878
		x"12",	--879
		x"e6",	--880
		x"41",	--881
		x"41",	--882
		x"41",	--883
		x"12",	--884
		x"12",	--885
		x"12",	--886
		x"4f",	--887
		x"93",	--888
		x"24",	--889
		x"4e",	--890
		x"53",	--891
		x"43",	--892
		x"4a",	--893
		x"5b",	--894
		x"4d",	--895
		x"11",	--896
		x"12",	--897
		x"e6",	--898
		x"99",	--899
		x"24",	--900
		x"53",	--901
		x"b0",	--902
		x"00",	--903
		x"20",	--904
		x"40",	--905
		x"00",	--906
		x"12",	--907
		x"e6",	--908
		x"3f",	--909
		x"40",	--910
		x"00",	--911
		x"12",	--912
		x"e6",	--913
		x"3f",	--914
		x"41",	--915
		x"41",	--916
		x"41",	--917
		x"41",	--918
		x"12",	--919
		x"12",	--920
		x"12",	--921
		x"4f",	--922
		x"93",	--923
		x"24",	--924
		x"4e",	--925
		x"53",	--926
		x"43",	--927
		x"4a",	--928
		x"11",	--929
		x"12",	--930
		x"e6",	--931
		x"99",	--932
		x"24",	--933
		x"53",	--934
		x"b0",	--935
		x"00",	--936
		x"23",	--937
		x"40",	--938
		x"00",	--939
		x"12",	--940
		x"e6",	--941
		x"4a",	--942
		x"11",	--943
		x"12",	--944
		x"e6",	--945
		x"99",	--946
		x"23",	--947
		x"41",	--948
		x"41",	--949
		x"41",	--950
		x"41",	--951
		x"12",	--952
		x"12",	--953
		x"12",	--954
		x"50",	--955
		x"ff",	--956
		x"4f",	--957
		x"93",	--958
		x"38",	--959
		x"90",	--960
		x"00",	--961
		x"38",	--962
		x"43",	--963
		x"41",	--964
		x"59",	--965
		x"40",	--966
		x"00",	--967
		x"4b",	--968
		x"12",	--969
		x"f6",	--970
		x"50",	--971
		x"00",	--972
		x"4f",	--973
		x"00",	--974
		x"53",	--975
		x"40",	--976
		x"00",	--977
		x"4b",	--978
		x"12",	--979
		x"f6",	--980
		x"4f",	--981
		x"90",	--982
		x"00",	--983
		x"37",	--984
		x"49",	--985
		x"53",	--986
		x"51",	--987
		x"40",	--988
		x"00",	--989
		x"4b",	--990
		x"12",	--991
		x"f6",	--992
		x"50",	--993
		x"00",	--994
		x"4f",	--995
		x"00",	--996
		x"53",	--997
		x"41",	--998
		x"5a",	--999
		x"4f",	--1000
		x"11",	--1001
		x"12",	--1002
		x"e6",	--1003
		x"93",	--1004
		x"23",	--1005
		x"50",	--1006
		x"00",	--1007
		x"41",	--1008
		x"41",	--1009
		x"41",	--1010
		x"41",	--1011
		x"40",	--1012
		x"00",	--1013
		x"12",	--1014
		x"e6",	--1015
		x"e3",	--1016
		x"53",	--1017
		x"3f",	--1018
		x"43",	--1019
		x"43",	--1020
		x"3f",	--1021
		x"12",	--1022
		x"12",	--1023
		x"12",	--1024
		x"41",	--1025
		x"52",	--1026
		x"4b",	--1027
		x"49",	--1028
		x"93",	--1029
		x"20",	--1030
		x"3c",	--1031
		x"11",	--1032
		x"12",	--1033
		x"e6",	--1034
		x"49",	--1035
		x"4a",	--1036
		x"53",	--1037
		x"4a",	--1038
		x"00",	--1039
		x"93",	--1040
		x"24",	--1041
		x"90",	--1042
		x"00",	--1043
		x"23",	--1044
		x"49",	--1045
		x"53",	--1046
		x"49",	--1047
		x"00",	--1048
		x"50",	--1049
		x"ff",	--1050
		x"90",	--1051
		x"00",	--1052
		x"2f",	--1053
		x"4f",	--1054
		x"5f",	--1055
		x"4f",	--1056
		x"f8",	--1057
		x"41",	--1058
		x"41",	--1059
		x"41",	--1060
		x"41",	--1061
		x"4b",	--1062
		x"52",	--1063
		x"4b",	--1064
		x"00",	--1065
		x"4b",	--1066
		x"12",	--1067
		x"e6",	--1068
		x"49",	--1069
		x"3f",	--1070
		x"4b",	--1071
		x"53",	--1072
		x"4b",	--1073
		x"12",	--1074
		x"e6",	--1075
		x"49",	--1076
		x"3f",	--1077
		x"4b",	--1078
		x"53",	--1079
		x"4f",	--1080
		x"49",	--1081
		x"93",	--1082
		x"27",	--1083
		x"53",	--1084
		x"11",	--1085
		x"12",	--1086
		x"e6",	--1087
		x"49",	--1088
		x"93",	--1089
		x"23",	--1090
		x"3f",	--1091
		x"4b",	--1092
		x"52",	--1093
		x"4b",	--1094
		x"00",	--1095
		x"4b",	--1096
		x"12",	--1097
		x"e7",	--1098
		x"49",	--1099
		x"3f",	--1100
		x"4b",	--1101
		x"53",	--1102
		x"4b",	--1103
		x"4e",	--1104
		x"10",	--1105
		x"11",	--1106
		x"10",	--1107
		x"11",	--1108
		x"12",	--1109
		x"e6",	--1110
		x"49",	--1111
		x"3f",	--1112
		x"4b",	--1113
		x"53",	--1114
		x"4b",	--1115
		x"12",	--1116
		x"e7",	--1117
		x"49",	--1118
		x"3f",	--1119
		x"4b",	--1120
		x"53",	--1121
		x"4b",	--1122
		x"12",	--1123
		x"e6",	--1124
		x"49",	--1125
		x"3f",	--1126
		x"4b",	--1127
		x"53",	--1128
		x"4b",	--1129
		x"12",	--1130
		x"e6",	--1131
		x"49",	--1132
		x"3f",	--1133
		x"4b",	--1134
		x"53",	--1135
		x"4b",	--1136
		x"12",	--1137
		x"e6",	--1138
		x"49",	--1139
		x"3f",	--1140
		x"40",	--1141
		x"00",	--1142
		x"12",	--1143
		x"e6",	--1144
		x"3f",	--1145
		x"12",	--1146
		x"12",	--1147
		x"42",	--1148
		x"02",	--1149
		x"42",	--1150
		x"00",	--1151
		x"03",	--1152
		x"42",	--1153
		x"02",	--1154
		x"90",	--1155
		x"00",	--1156
		x"34",	--1157
		x"53",	--1158
		x"02",	--1159
		x"42",	--1160
		x"02",	--1161
		x"42",	--1162
		x"02",	--1163
		x"9f",	--1164
		x"20",	--1165
		x"53",	--1166
		x"02",	--1167
		x"40",	--1168
		x"00",	--1169
		x"00",	--1170
		x"c0",	--1171
		x"00",	--1172
		x"00",	--1173
		x"41",	--1174
		x"41",	--1175
		x"c0",	--1176
		x"00",	--1177
		x"00",	--1178
		x"13",	--1179
		x"43",	--1180
		x"02",	--1181
		x"3f",	--1182
		x"40",	--1183
		x"09",	--1184
		x"00",	--1185
		x"40",	--1186
		x"00",	--1187
		x"00",	--1188
		x"41",	--1189
		x"42",	--1190
		x"02",	--1191
		x"42",	--1192
		x"02",	--1193
		x"9f",	--1194
		x"38",	--1195
		x"42",	--1196
		x"02",	--1197
		x"82",	--1198
		x"02",	--1199
		x"41",	--1200
		x"42",	--1201
		x"02",	--1202
		x"42",	--1203
		x"02",	--1204
		x"40",	--1205
		x"00",	--1206
		x"8d",	--1207
		x"8e",	--1208
		x"41",	--1209
		x"42",	--1210
		x"02",	--1211
		x"4f",	--1212
		x"03",	--1213
		x"42",	--1214
		x"02",	--1215
		x"42",	--1216
		x"02",	--1217
		x"9e",	--1218
		x"24",	--1219
		x"42",	--1220
		x"02",	--1221
		x"90",	--1222
		x"00",	--1223
		x"38",	--1224
		x"43",	--1225
		x"02",	--1226
		x"41",	--1227
		x"53",	--1228
		x"02",	--1229
		x"41",	--1230
		x"43",	--1231
		x"41",	--1232
		x"12",	--1233
		x"12",	--1234
		x"4e",	--1235
		x"4f",	--1236
		x"43",	--1237
		x"40",	--1238
		x"4f",	--1239
		x"12",	--1240
		x"f0",	--1241
		x"93",	--1242
		x"34",	--1243
		x"4a",	--1244
		x"4b",	--1245
		x"12",	--1246
		x"f0",	--1247
		x"41",	--1248
		x"41",	--1249
		x"41",	--1250
		x"43",	--1251
		x"40",	--1252
		x"4f",	--1253
		x"4a",	--1254
		x"4b",	--1255
		x"12",	--1256
		x"ec",	--1257
		x"12",	--1258
		x"f0",	--1259
		x"53",	--1260
		x"60",	--1261
		x"80",	--1262
		x"41",	--1263
		x"41",	--1264
		x"41",	--1265
		x"12",	--1266
		x"12",	--1267
		x"12",	--1268
		x"12",	--1269
		x"12",	--1270
		x"12",	--1271
		x"12",	--1272
		x"12",	--1273
		x"50",	--1274
		x"ff",	--1275
		x"4d",	--1276
		x"4f",	--1277
		x"93",	--1278
		x"28",	--1279
		x"4e",	--1280
		x"93",	--1281
		x"28",	--1282
		x"92",	--1283
		x"20",	--1284
		x"40",	--1285
		x"ec",	--1286
		x"92",	--1287
		x"24",	--1288
		x"93",	--1289
		x"24",	--1290
		x"93",	--1291
		x"24",	--1292
		x"4f",	--1293
		x"00",	--1294
		x"00",	--1295
		x"4e",	--1296
		x"00",	--1297
		x"4f",	--1298
		x"00",	--1299
		x"4f",	--1300
		x"00",	--1301
		x"4e",	--1302
		x"00",	--1303
		x"4e",	--1304
		x"00",	--1305
		x"41",	--1306
		x"8b",	--1307
		x"4c",	--1308
		x"93",	--1309
		x"38",	--1310
		x"90",	--1311
		x"00",	--1312
		x"34",	--1313
		x"93",	--1314
		x"38",	--1315
		x"46",	--1316
		x"00",	--1317
		x"47",	--1318
		x"00",	--1319
		x"49",	--1320
		x"f0",	--1321
		x"00",	--1322
		x"24",	--1323
		x"46",	--1324
		x"47",	--1325
		x"c3",	--1326
		x"10",	--1327
		x"10",	--1328
		x"53",	--1329
		x"23",	--1330
		x"4a",	--1331
		x"00",	--1332
		x"4b",	--1333
		x"00",	--1334
		x"43",	--1335
		x"43",	--1336
		x"f0",	--1337
		x"00",	--1338
		x"24",	--1339
		x"5c",	--1340
		x"6d",	--1341
		x"53",	--1342
		x"23",	--1343
		x"53",	--1344
		x"63",	--1345
		x"f6",	--1346
		x"f7",	--1347
		x"43",	--1348
		x"43",	--1349
		x"93",	--1350
		x"20",	--1351
		x"93",	--1352
		x"24",	--1353
		x"41",	--1354
		x"00",	--1355
		x"41",	--1356
		x"00",	--1357
		x"da",	--1358
		x"db",	--1359
		x"4f",	--1360
		x"00",	--1361
		x"9e",	--1362
		x"00",	--1363
		x"20",	--1364
		x"4f",	--1365
		x"00",	--1366
		x"41",	--1367
		x"00",	--1368
		x"46",	--1369
		x"47",	--1370
		x"54",	--1371
		x"65",	--1372
		x"4e",	--1373
		x"00",	--1374
		x"4f",	--1375
		x"00",	--1376
		x"40",	--1377
		x"00",	--1378
		x"00",	--1379
		x"93",	--1380
		x"38",	--1381
		x"48",	--1382
		x"50",	--1383
		x"00",	--1384
		x"41",	--1385
		x"41",	--1386
		x"41",	--1387
		x"41",	--1388
		x"41",	--1389
		x"41",	--1390
		x"41",	--1391
		x"41",	--1392
		x"41",	--1393
		x"91",	--1394
		x"38",	--1395
		x"4b",	--1396
		x"00",	--1397
		x"43",	--1398
		x"43",	--1399
		x"4f",	--1400
		x"00",	--1401
		x"9e",	--1402
		x"00",	--1403
		x"27",	--1404
		x"93",	--1405
		x"24",	--1406
		x"46",	--1407
		x"47",	--1408
		x"84",	--1409
		x"75",	--1410
		x"93",	--1411
		x"38",	--1412
		x"43",	--1413
		x"00",	--1414
		x"41",	--1415
		x"00",	--1416
		x"4e",	--1417
		x"00",	--1418
		x"4f",	--1419
		x"00",	--1420
		x"4e",	--1421
		x"4f",	--1422
		x"53",	--1423
		x"63",	--1424
		x"90",	--1425
		x"3f",	--1426
		x"28",	--1427
		x"90",	--1428
		x"40",	--1429
		x"2c",	--1430
		x"93",	--1431
		x"2c",	--1432
		x"48",	--1433
		x"00",	--1434
		x"53",	--1435
		x"5e",	--1436
		x"6f",	--1437
		x"4b",	--1438
		x"53",	--1439
		x"4e",	--1440
		x"4f",	--1441
		x"53",	--1442
		x"63",	--1443
		x"90",	--1444
		x"3f",	--1445
		x"2b",	--1446
		x"24",	--1447
		x"4e",	--1448
		x"00",	--1449
		x"4f",	--1450
		x"00",	--1451
		x"4a",	--1452
		x"00",	--1453
		x"40",	--1454
		x"00",	--1455
		x"00",	--1456
		x"93",	--1457
		x"37",	--1458
		x"4e",	--1459
		x"4f",	--1460
		x"f3",	--1461
		x"f3",	--1462
		x"c3",	--1463
		x"10",	--1464
		x"10",	--1465
		x"4c",	--1466
		x"4d",	--1467
		x"de",	--1468
		x"df",	--1469
		x"4a",	--1470
		x"00",	--1471
		x"4b",	--1472
		x"00",	--1473
		x"53",	--1474
		x"00",	--1475
		x"48",	--1476
		x"3f",	--1477
		x"93",	--1478
		x"23",	--1479
		x"4f",	--1480
		x"00",	--1481
		x"4f",	--1482
		x"00",	--1483
		x"00",	--1484
		x"4f",	--1485
		x"00",	--1486
		x"00",	--1487
		x"4f",	--1488
		x"00",	--1489
		x"00",	--1490
		x"4e",	--1491
		x"00",	--1492
		x"ff",	--1493
		x"00",	--1494
		x"4e",	--1495
		x"00",	--1496
		x"4d",	--1497
		x"3f",	--1498
		x"43",	--1499
		x"43",	--1500
		x"3f",	--1501
		x"e3",	--1502
		x"53",	--1503
		x"90",	--1504
		x"00",	--1505
		x"37",	--1506
		x"3f",	--1507
		x"93",	--1508
		x"2b",	--1509
		x"3f",	--1510
		x"44",	--1511
		x"45",	--1512
		x"86",	--1513
		x"77",	--1514
		x"3f",	--1515
		x"4e",	--1516
		x"3f",	--1517
		x"43",	--1518
		x"00",	--1519
		x"41",	--1520
		x"00",	--1521
		x"e3",	--1522
		x"e3",	--1523
		x"53",	--1524
		x"63",	--1525
		x"4e",	--1526
		x"00",	--1527
		x"4f",	--1528
		x"00",	--1529
		x"3f",	--1530
		x"93",	--1531
		x"27",	--1532
		x"59",	--1533
		x"00",	--1534
		x"44",	--1535
		x"00",	--1536
		x"45",	--1537
		x"00",	--1538
		x"49",	--1539
		x"f0",	--1540
		x"00",	--1541
		x"24",	--1542
		x"4d",	--1543
		x"44",	--1544
		x"45",	--1545
		x"c3",	--1546
		x"10",	--1547
		x"10",	--1548
		x"53",	--1549
		x"23",	--1550
		x"4c",	--1551
		x"00",	--1552
		x"4d",	--1553
		x"00",	--1554
		x"43",	--1555
		x"43",	--1556
		x"f0",	--1557
		x"00",	--1558
		x"24",	--1559
		x"5c",	--1560
		x"6d",	--1561
		x"53",	--1562
		x"23",	--1563
		x"53",	--1564
		x"63",	--1565
		x"f4",	--1566
		x"f5",	--1567
		x"43",	--1568
		x"43",	--1569
		x"93",	--1570
		x"20",	--1571
		x"93",	--1572
		x"20",	--1573
		x"43",	--1574
		x"43",	--1575
		x"41",	--1576
		x"00",	--1577
		x"41",	--1578
		x"00",	--1579
		x"da",	--1580
		x"db",	--1581
		x"3f",	--1582
		x"43",	--1583
		x"43",	--1584
		x"3f",	--1585
		x"92",	--1586
		x"23",	--1587
		x"9e",	--1588
		x"00",	--1589
		x"00",	--1590
		x"27",	--1591
		x"40",	--1592
		x"f9",	--1593
		x"3f",	--1594
		x"50",	--1595
		x"ff",	--1596
		x"4e",	--1597
		x"00",	--1598
		x"4f",	--1599
		x"00",	--1600
		x"4c",	--1601
		x"00",	--1602
		x"4d",	--1603
		x"00",	--1604
		x"41",	--1605
		x"50",	--1606
		x"00",	--1607
		x"41",	--1608
		x"52",	--1609
		x"12",	--1610
		x"f4",	--1611
		x"41",	--1612
		x"50",	--1613
		x"00",	--1614
		x"41",	--1615
		x"12",	--1616
		x"f4",	--1617
		x"41",	--1618
		x"52",	--1619
		x"41",	--1620
		x"50",	--1621
		x"00",	--1622
		x"41",	--1623
		x"50",	--1624
		x"00",	--1625
		x"12",	--1626
		x"e9",	--1627
		x"12",	--1628
		x"f2",	--1629
		x"50",	--1630
		x"00",	--1631
		x"41",	--1632
		x"50",	--1633
		x"ff",	--1634
		x"4e",	--1635
		x"00",	--1636
		x"4f",	--1637
		x"00",	--1638
		x"4c",	--1639
		x"00",	--1640
		x"4d",	--1641
		x"00",	--1642
		x"41",	--1643
		x"50",	--1644
		x"00",	--1645
		x"41",	--1646
		x"52",	--1647
		x"12",	--1648
		x"f4",	--1649
		x"41",	--1650
		x"50",	--1651
		x"00",	--1652
		x"41",	--1653
		x"12",	--1654
		x"f4",	--1655
		x"e3",	--1656
		x"00",	--1657
		x"41",	--1658
		x"52",	--1659
		x"41",	--1660
		x"50",	--1661
		x"00",	--1662
		x"41",	--1663
		x"50",	--1664
		x"00",	--1665
		x"12",	--1666
		x"e9",	--1667
		x"12",	--1668
		x"f2",	--1669
		x"50",	--1670
		x"00",	--1671
		x"41",	--1672
		x"12",	--1673
		x"12",	--1674
		x"12",	--1675
		x"12",	--1676
		x"12",	--1677
		x"12",	--1678
		x"12",	--1679
		x"12",	--1680
		x"50",	--1681
		x"ff",	--1682
		x"4e",	--1683
		x"00",	--1684
		x"4f",	--1685
		x"00",	--1686
		x"4c",	--1687
		x"00",	--1688
		x"4d",	--1689
		x"00",	--1690
		x"41",	--1691
		x"50",	--1692
		x"00",	--1693
		x"41",	--1694
		x"52",	--1695
		x"12",	--1696
		x"f4",	--1697
		x"41",	--1698
		x"50",	--1699
		x"00",	--1700
		x"41",	--1701
		x"12",	--1702
		x"f4",	--1703
		x"41",	--1704
		x"00",	--1705
		x"93",	--1706
		x"28",	--1707
		x"41",	--1708
		x"00",	--1709
		x"93",	--1710
		x"28",	--1711
		x"92",	--1712
		x"24",	--1713
		x"92",	--1714
		x"24",	--1715
		x"93",	--1716
		x"24",	--1717
		x"93",	--1718
		x"24",	--1719
		x"41",	--1720
		x"00",	--1721
		x"41",	--1722
		x"00",	--1723
		x"41",	--1724
		x"00",	--1725
		x"41",	--1726
		x"00",	--1727
		x"40",	--1728
		x"00",	--1729
		x"43",	--1730
		x"43",	--1731
		x"43",	--1732
		x"43",	--1733
		x"43",	--1734
		x"00",	--1735
		x"43",	--1736
		x"00",	--1737
		x"43",	--1738
		x"43",	--1739
		x"4c",	--1740
		x"00",	--1741
		x"3c",	--1742
		x"58",	--1743
		x"69",	--1744
		x"c3",	--1745
		x"10",	--1746
		x"10",	--1747
		x"53",	--1748
		x"00",	--1749
		x"24",	--1750
		x"b3",	--1751
		x"24",	--1752
		x"58",	--1753
		x"69",	--1754
		x"56",	--1755
		x"67",	--1756
		x"43",	--1757
		x"43",	--1758
		x"99",	--1759
		x"28",	--1760
		x"24",	--1761
		x"43",	--1762
		x"43",	--1763
		x"5c",	--1764
		x"6d",	--1765
		x"56",	--1766
		x"67",	--1767
		x"93",	--1768
		x"37",	--1769
		x"d3",	--1770
		x"d3",	--1771
		x"3f",	--1772
		x"98",	--1773
		x"2b",	--1774
		x"3f",	--1775
		x"4a",	--1776
		x"00",	--1777
		x"4b",	--1778
		x"00",	--1779
		x"4f",	--1780
		x"41",	--1781
		x"00",	--1782
		x"51",	--1783
		x"00",	--1784
		x"4a",	--1785
		x"53",	--1786
		x"46",	--1787
		x"00",	--1788
		x"43",	--1789
		x"91",	--1790
		x"00",	--1791
		x"00",	--1792
		x"24",	--1793
		x"4d",	--1794
		x"00",	--1795
		x"93",	--1796
		x"38",	--1797
		x"90",	--1798
		x"40",	--1799
		x"2c",	--1800
		x"41",	--1801
		x"00",	--1802
		x"53",	--1803
		x"41",	--1804
		x"00",	--1805
		x"41",	--1806
		x"00",	--1807
		x"4d",	--1808
		x"5e",	--1809
		x"6f",	--1810
		x"93",	--1811
		x"38",	--1812
		x"5a",	--1813
		x"6b",	--1814
		x"53",	--1815
		x"90",	--1816
		x"40",	--1817
		x"2b",	--1818
		x"4a",	--1819
		x"00",	--1820
		x"4b",	--1821
		x"00",	--1822
		x"4c",	--1823
		x"00",	--1824
		x"4e",	--1825
		x"4f",	--1826
		x"f0",	--1827
		x"00",	--1828
		x"f3",	--1829
		x"90",	--1830
		x"00",	--1831
		x"24",	--1832
		x"4e",	--1833
		x"00",	--1834
		x"4f",	--1835
		x"00",	--1836
		x"40",	--1837
		x"00",	--1838
		x"00",	--1839
		x"41",	--1840
		x"52",	--1841
		x"12",	--1842
		x"f2",	--1843
		x"50",	--1844
		x"00",	--1845
		x"41",	--1846
		x"41",	--1847
		x"41",	--1848
		x"41",	--1849
		x"41",	--1850
		x"41",	--1851
		x"41",	--1852
		x"41",	--1853
		x"41",	--1854
		x"d3",	--1855
		x"d3",	--1856
		x"3f",	--1857
		x"50",	--1858
		x"00",	--1859
		x"4a",	--1860
		x"b3",	--1861
		x"24",	--1862
		x"41",	--1863
		x"00",	--1864
		x"41",	--1865
		x"00",	--1866
		x"c3",	--1867
		x"10",	--1868
		x"10",	--1869
		x"4c",	--1870
		x"4d",	--1871
		x"d3",	--1872
		x"d0",	--1873
		x"80",	--1874
		x"46",	--1875
		x"00",	--1876
		x"47",	--1877
		x"00",	--1878
		x"c3",	--1879
		x"10",	--1880
		x"10",	--1881
		x"53",	--1882
		x"93",	--1883
		x"3b",	--1884
		x"48",	--1885
		x"00",	--1886
		x"3f",	--1887
		x"93",	--1888
		x"24",	--1889
		x"43",	--1890
		x"91",	--1891
		x"00",	--1892
		x"00",	--1893
		x"24",	--1894
		x"4f",	--1895
		x"00",	--1896
		x"41",	--1897
		x"50",	--1898
		x"00",	--1899
		x"3f",	--1900
		x"93",	--1901
		x"23",	--1902
		x"4e",	--1903
		x"4f",	--1904
		x"f0",	--1905
		x"00",	--1906
		x"f3",	--1907
		x"93",	--1908
		x"23",	--1909
		x"93",	--1910
		x"23",	--1911
		x"93",	--1912
		x"00",	--1913
		x"20",	--1914
		x"93",	--1915
		x"00",	--1916
		x"27",	--1917
		x"50",	--1918
		x"00",	--1919
		x"63",	--1920
		x"f0",	--1921
		x"ff",	--1922
		x"f3",	--1923
		x"3f",	--1924
		x"43",	--1925
		x"3f",	--1926
		x"43",	--1927
		x"3f",	--1928
		x"43",	--1929
		x"91",	--1930
		x"00",	--1931
		x"00",	--1932
		x"24",	--1933
		x"4f",	--1934
		x"00",	--1935
		x"41",	--1936
		x"50",	--1937
		x"00",	--1938
		x"3f",	--1939
		x"43",	--1940
		x"3f",	--1941
		x"93",	--1942
		x"23",	--1943
		x"40",	--1944
		x"f9",	--1945
		x"3f",	--1946
		x"12",	--1947
		x"12",	--1948
		x"12",	--1949
		x"12",	--1950
		x"12",	--1951
		x"50",	--1952
		x"ff",	--1953
		x"4e",	--1954
		x"00",	--1955
		x"4f",	--1956
		x"00",	--1957
		x"4c",	--1958
		x"00",	--1959
		x"4d",	--1960
		x"00",	--1961
		x"41",	--1962
		x"50",	--1963
		x"00",	--1964
		x"41",	--1965
		x"52",	--1966
		x"12",	--1967
		x"f4",	--1968
		x"41",	--1969
		x"52",	--1970
		x"41",	--1971
		x"12",	--1972
		x"f4",	--1973
		x"41",	--1974
		x"00",	--1975
		x"93",	--1976
		x"28",	--1977
		x"41",	--1978
		x"00",	--1979
		x"93",	--1980
		x"28",	--1981
		x"e1",	--1982
		x"00",	--1983
		x"00",	--1984
		x"92",	--1985
		x"24",	--1986
		x"93",	--1987
		x"24",	--1988
		x"92",	--1989
		x"24",	--1990
		x"93",	--1991
		x"24",	--1992
		x"41",	--1993
		x"00",	--1994
		x"81",	--1995
		x"00",	--1996
		x"4d",	--1997
		x"00",	--1998
		x"41",	--1999
		x"00",	--2000
		x"41",	--2001
		x"00",	--2002
		x"41",	--2003
		x"00",	--2004
		x"41",	--2005
		x"00",	--2006
		x"99",	--2007
		x"2c",	--2008
		x"5e",	--2009
		x"6f",	--2010
		x"53",	--2011
		x"4d",	--2012
		x"00",	--2013
		x"40",	--2014
		x"00",	--2015
		x"43",	--2016
		x"40",	--2017
		x"40",	--2018
		x"43",	--2019
		x"43",	--2020
		x"3c",	--2021
		x"dc",	--2022
		x"dd",	--2023
		x"88",	--2024
		x"79",	--2025
		x"c3",	--2026
		x"10",	--2027
		x"10",	--2028
		x"5e",	--2029
		x"6f",	--2030
		x"53",	--2031
		x"24",	--2032
		x"99",	--2033
		x"2b",	--2034
		x"23",	--2035
		x"98",	--2036
		x"2b",	--2037
		x"3f",	--2038
		x"9f",	--2039
		x"2b",	--2040
		x"98",	--2041
		x"2f",	--2042
		x"3f",	--2043
		x"4a",	--2044
		x"4b",	--2045
		x"f0",	--2046
		x"00",	--2047
		x"f3",	--2048
		x"90",	--2049
		x"00",	--2050
		x"24",	--2051
		x"4a",	--2052
		x"00",	--2053
		x"4b",	--2054
		x"00",	--2055
		x"41",	--2056
		x"50",	--2057
		x"00",	--2058
		x"12",	--2059
		x"f2",	--2060
		x"50",	--2061
		x"00",	--2062
		x"41",	--2063
		x"41",	--2064
		x"41",	--2065
		x"41",	--2066
		x"41",	--2067
		x"41",	--2068
		x"42",	--2069
		x"00",	--2070
		x"41",	--2071
		x"50",	--2072
		x"00",	--2073
		x"3f",	--2074
		x"9e",	--2075
		x"23",	--2076
		x"40",	--2077
		x"f9",	--2078
		x"3f",	--2079
		x"93",	--2080
		x"23",	--2081
		x"4a",	--2082
		x"4b",	--2083
		x"f0",	--2084
		x"00",	--2085
		x"f3",	--2086
		x"93",	--2087
		x"23",	--2088
		x"93",	--2089
		x"23",	--2090
		x"93",	--2091
		x"20",	--2092
		x"93",	--2093
		x"27",	--2094
		x"50",	--2095
		x"00",	--2096
		x"63",	--2097
		x"f0",	--2098
		x"ff",	--2099
		x"f3",	--2100
		x"3f",	--2101
		x"43",	--2102
		x"00",	--2103
		x"43",	--2104
		x"00",	--2105
		x"43",	--2106
		x"00",	--2107
		x"41",	--2108
		x"50",	--2109
		x"00",	--2110
		x"3f",	--2111
		x"41",	--2112
		x"52",	--2113
		x"3f",	--2114
		x"50",	--2115
		x"ff",	--2116
		x"4e",	--2117
		x"00",	--2118
		x"4f",	--2119
		x"00",	--2120
		x"4c",	--2121
		x"00",	--2122
		x"4d",	--2123
		x"00",	--2124
		x"41",	--2125
		x"50",	--2126
		x"00",	--2127
		x"41",	--2128
		x"52",	--2129
		x"12",	--2130
		x"f4",	--2131
		x"41",	--2132
		x"52",	--2133
		x"41",	--2134
		x"12",	--2135
		x"f4",	--2136
		x"93",	--2137
		x"00",	--2138
		x"28",	--2139
		x"93",	--2140
		x"00",	--2141
		x"28",	--2142
		x"41",	--2143
		x"52",	--2144
		x"41",	--2145
		x"50",	--2146
		x"00",	--2147
		x"12",	--2148
		x"f5",	--2149
		x"50",	--2150
		x"00",	--2151
		x"41",	--2152
		x"43",	--2153
		x"3f",	--2154
		x"50",	--2155
		x"ff",	--2156
		x"4e",	--2157
		x"00",	--2158
		x"4f",	--2159
		x"00",	--2160
		x"41",	--2161
		x"52",	--2162
		x"41",	--2163
		x"12",	--2164
		x"f4",	--2165
		x"41",	--2166
		x"00",	--2167
		x"93",	--2168
		x"24",	--2169
		x"28",	--2170
		x"92",	--2171
		x"24",	--2172
		x"41",	--2173
		x"00",	--2174
		x"93",	--2175
		x"38",	--2176
		x"90",	--2177
		x"00",	--2178
		x"38",	--2179
		x"93",	--2180
		x"00",	--2181
		x"20",	--2182
		x"43",	--2183
		x"40",	--2184
		x"7f",	--2185
		x"50",	--2186
		x"00",	--2187
		x"41",	--2188
		x"41",	--2189
		x"00",	--2190
		x"41",	--2191
		x"00",	--2192
		x"40",	--2193
		x"00",	--2194
		x"8d",	--2195
		x"4c",	--2196
		x"f0",	--2197
		x"00",	--2198
		x"20",	--2199
		x"93",	--2200
		x"00",	--2201
		x"27",	--2202
		x"e3",	--2203
		x"e3",	--2204
		x"53",	--2205
		x"63",	--2206
		x"50",	--2207
		x"00",	--2208
		x"41",	--2209
		x"43",	--2210
		x"43",	--2211
		x"50",	--2212
		x"00",	--2213
		x"41",	--2214
		x"c3",	--2215
		x"10",	--2216
		x"10",	--2217
		x"53",	--2218
		x"23",	--2219
		x"3f",	--2220
		x"43",	--2221
		x"40",	--2222
		x"80",	--2223
		x"50",	--2224
		x"00",	--2225
		x"41",	--2226
		x"12",	--2227
		x"12",	--2228
		x"12",	--2229
		x"12",	--2230
		x"82",	--2231
		x"4e",	--2232
		x"4f",	--2233
		x"43",	--2234
		x"00",	--2235
		x"93",	--2236
		x"20",	--2237
		x"93",	--2238
		x"20",	--2239
		x"43",	--2240
		x"00",	--2241
		x"41",	--2242
		x"12",	--2243
		x"f2",	--2244
		x"52",	--2245
		x"41",	--2246
		x"41",	--2247
		x"41",	--2248
		x"41",	--2249
		x"41",	--2250
		x"40",	--2251
		x"00",	--2252
		x"00",	--2253
		x"40",	--2254
		x"00",	--2255
		x"00",	--2256
		x"4a",	--2257
		x"00",	--2258
		x"4b",	--2259
		x"00",	--2260
		x"4a",	--2261
		x"4b",	--2262
		x"12",	--2263
		x"f2",	--2264
		x"53",	--2265
		x"93",	--2266
		x"38",	--2267
		x"27",	--2268
		x"4a",	--2269
		x"00",	--2270
		x"4b",	--2271
		x"00",	--2272
		x"4f",	--2273
		x"f0",	--2274
		x"00",	--2275
		x"20",	--2276
		x"40",	--2277
		x"00",	--2278
		x"8f",	--2279
		x"4e",	--2280
		x"00",	--2281
		x"3f",	--2282
		x"51",	--2283
		x"00",	--2284
		x"00",	--2285
		x"61",	--2286
		x"00",	--2287
		x"00",	--2288
		x"53",	--2289
		x"23",	--2290
		x"3f",	--2291
		x"4f",	--2292
		x"e3",	--2293
		x"53",	--2294
		x"43",	--2295
		x"43",	--2296
		x"4e",	--2297
		x"f0",	--2298
		x"00",	--2299
		x"24",	--2300
		x"5c",	--2301
		x"6d",	--2302
		x"53",	--2303
		x"23",	--2304
		x"53",	--2305
		x"63",	--2306
		x"fa",	--2307
		x"fb",	--2308
		x"43",	--2309
		x"43",	--2310
		x"93",	--2311
		x"20",	--2312
		x"93",	--2313
		x"20",	--2314
		x"43",	--2315
		x"43",	--2316
		x"f0",	--2317
		x"00",	--2318
		x"20",	--2319
		x"48",	--2320
		x"49",	--2321
		x"da",	--2322
		x"db",	--2323
		x"4d",	--2324
		x"00",	--2325
		x"4e",	--2326
		x"00",	--2327
		x"40",	--2328
		x"00",	--2329
		x"8f",	--2330
		x"4e",	--2331
		x"00",	--2332
		x"3f",	--2333
		x"c3",	--2334
		x"10",	--2335
		x"10",	--2336
		x"53",	--2337
		x"23",	--2338
		x"3f",	--2339
		x"12",	--2340
		x"12",	--2341
		x"12",	--2342
		x"93",	--2343
		x"2c",	--2344
		x"90",	--2345
		x"01",	--2346
		x"28",	--2347
		x"40",	--2348
		x"00",	--2349
		x"43",	--2350
		x"42",	--2351
		x"4e",	--2352
		x"4f",	--2353
		x"49",	--2354
		x"93",	--2355
		x"20",	--2356
		x"50",	--2357
		x"f9",	--2358
		x"4c",	--2359
		x"43",	--2360
		x"8e",	--2361
		x"7f",	--2362
		x"4a",	--2363
		x"41",	--2364
		x"41",	--2365
		x"41",	--2366
		x"41",	--2367
		x"90",	--2368
		x"01",	--2369
		x"28",	--2370
		x"42",	--2371
		x"43",	--2372
		x"40",	--2373
		x"00",	--2374
		x"4e",	--2375
		x"4f",	--2376
		x"49",	--2377
		x"93",	--2378
		x"27",	--2379
		x"c3",	--2380
		x"10",	--2381
		x"10",	--2382
		x"53",	--2383
		x"23",	--2384
		x"3f",	--2385
		x"40",	--2386
		x"00",	--2387
		x"43",	--2388
		x"40",	--2389
		x"00",	--2390
		x"3f",	--2391
		x"40",	--2392
		x"00",	--2393
		x"43",	--2394
		x"43",	--2395
		x"3f",	--2396
		x"12",	--2397
		x"12",	--2398
		x"12",	--2399
		x"12",	--2400
		x"12",	--2401
		x"4f",	--2402
		x"4f",	--2403
		x"00",	--2404
		x"4f",	--2405
		x"00",	--2406
		x"4d",	--2407
		x"00",	--2408
		x"4d",	--2409
		x"93",	--2410
		x"28",	--2411
		x"92",	--2412
		x"24",	--2413
		x"93",	--2414
		x"24",	--2415
		x"93",	--2416
		x"24",	--2417
		x"4d",	--2418
		x"00",	--2419
		x"90",	--2420
		x"ff",	--2421
		x"38",	--2422
		x"90",	--2423
		x"00",	--2424
		x"34",	--2425
		x"4e",	--2426
		x"4f",	--2427
		x"f0",	--2428
		x"00",	--2429
		x"f3",	--2430
		x"90",	--2431
		x"00",	--2432
		x"24",	--2433
		x"50",	--2434
		x"00",	--2435
		x"63",	--2436
		x"93",	--2437
		x"38",	--2438
		x"4b",	--2439
		x"50",	--2440
		x"00",	--2441
		x"c3",	--2442
		x"10",	--2443
		x"10",	--2444
		x"c3",	--2445
		x"10",	--2446
		x"10",	--2447
		x"c3",	--2448
		x"10",	--2449
		x"10",	--2450
		x"c3",	--2451
		x"10",	--2452
		x"10",	--2453
		x"c3",	--2454
		x"10",	--2455
		x"10",	--2456
		x"c3",	--2457
		x"10",	--2458
		x"10",	--2459
		x"c3",	--2460
		x"10",	--2461
		x"10",	--2462
		x"f3",	--2463
		x"f0",	--2464
		x"00",	--2465
		x"4d",	--2466
		x"3c",	--2467
		x"93",	--2468
		x"23",	--2469
		x"43",	--2470
		x"43",	--2471
		x"43",	--2472
		x"4d",	--2473
		x"5d",	--2474
		x"5d",	--2475
		x"5d",	--2476
		x"5d",	--2477
		x"5d",	--2478
		x"5d",	--2479
		x"5d",	--2480
		x"4f",	--2481
		x"f0",	--2482
		x"00",	--2483
		x"dd",	--2484
		x"4a",	--2485
		x"11",	--2486
		x"43",	--2487
		x"10",	--2488
		x"4c",	--2489
		x"df",	--2490
		x"4d",	--2491
		x"41",	--2492
		x"41",	--2493
		x"41",	--2494
		x"41",	--2495
		x"41",	--2496
		x"41",	--2497
		x"93",	--2498
		x"23",	--2499
		x"4e",	--2500
		x"4f",	--2501
		x"f0",	--2502
		x"00",	--2503
		x"f3",	--2504
		x"93",	--2505
		x"20",	--2506
		x"93",	--2507
		x"27",	--2508
		x"50",	--2509
		x"00",	--2510
		x"63",	--2511
		x"3f",	--2512
		x"c3",	--2513
		x"10",	--2514
		x"10",	--2515
		x"4b",	--2516
		x"50",	--2517
		x"00",	--2518
		x"3f",	--2519
		x"43",	--2520
		x"43",	--2521
		x"43",	--2522
		x"3f",	--2523
		x"d3",	--2524
		x"d0",	--2525
		x"00",	--2526
		x"f3",	--2527
		x"f0",	--2528
		x"00",	--2529
		x"43",	--2530
		x"3f",	--2531
		x"40",	--2532
		x"ff",	--2533
		x"8b",	--2534
		x"90",	--2535
		x"00",	--2536
		x"34",	--2537
		x"4e",	--2538
		x"4f",	--2539
		x"47",	--2540
		x"f0",	--2541
		x"00",	--2542
		x"24",	--2543
		x"c3",	--2544
		x"10",	--2545
		x"10",	--2546
		x"53",	--2547
		x"23",	--2548
		x"43",	--2549
		x"43",	--2550
		x"f0",	--2551
		x"00",	--2552
		x"24",	--2553
		x"58",	--2554
		x"69",	--2555
		x"53",	--2556
		x"23",	--2557
		x"53",	--2558
		x"63",	--2559
		x"fe",	--2560
		x"ff",	--2561
		x"43",	--2562
		x"43",	--2563
		x"93",	--2564
		x"20",	--2565
		x"93",	--2566
		x"20",	--2567
		x"43",	--2568
		x"43",	--2569
		x"4e",	--2570
		x"4f",	--2571
		x"dc",	--2572
		x"dd",	--2573
		x"48",	--2574
		x"49",	--2575
		x"f0",	--2576
		x"00",	--2577
		x"f3",	--2578
		x"90",	--2579
		x"00",	--2580
		x"24",	--2581
		x"50",	--2582
		x"00",	--2583
		x"63",	--2584
		x"48",	--2585
		x"49",	--2586
		x"c3",	--2587
		x"10",	--2588
		x"10",	--2589
		x"c3",	--2590
		x"10",	--2591
		x"10",	--2592
		x"c3",	--2593
		x"10",	--2594
		x"10",	--2595
		x"c3",	--2596
		x"10",	--2597
		x"10",	--2598
		x"c3",	--2599
		x"10",	--2600
		x"10",	--2601
		x"c3",	--2602
		x"10",	--2603
		x"10",	--2604
		x"c3",	--2605
		x"10",	--2606
		x"10",	--2607
		x"f3",	--2608
		x"f0",	--2609
		x"00",	--2610
		x"43",	--2611
		x"90",	--2612
		x"40",	--2613
		x"2f",	--2614
		x"43",	--2615
		x"3f",	--2616
		x"43",	--2617
		x"43",	--2618
		x"3f",	--2619
		x"93",	--2620
		x"23",	--2621
		x"48",	--2622
		x"49",	--2623
		x"f0",	--2624
		x"00",	--2625
		x"f3",	--2626
		x"93",	--2627
		x"24",	--2628
		x"50",	--2629
		x"00",	--2630
		x"63",	--2631
		x"3f",	--2632
		x"93",	--2633
		x"27",	--2634
		x"3f",	--2635
		x"12",	--2636
		x"12",	--2637
		x"4f",	--2638
		x"4f",	--2639
		x"00",	--2640
		x"f0",	--2641
		x"00",	--2642
		x"4f",	--2643
		x"00",	--2644
		x"c3",	--2645
		x"10",	--2646
		x"c3",	--2647
		x"10",	--2648
		x"c3",	--2649
		x"10",	--2650
		x"c3",	--2651
		x"10",	--2652
		x"c3",	--2653
		x"10",	--2654
		x"c3",	--2655
		x"10",	--2656
		x"c3",	--2657
		x"10",	--2658
		x"4d",	--2659
		x"4f",	--2660
		x"00",	--2661
		x"b0",	--2662
		x"00",	--2663
		x"43",	--2664
		x"6f",	--2665
		x"4f",	--2666
		x"00",	--2667
		x"93",	--2668
		x"20",	--2669
		x"93",	--2670
		x"24",	--2671
		x"40",	--2672
		x"ff",	--2673
		x"00",	--2674
		x"4a",	--2675
		x"4b",	--2676
		x"5c",	--2677
		x"6d",	--2678
		x"5c",	--2679
		x"6d",	--2680
		x"5c",	--2681
		x"6d",	--2682
		x"5c",	--2683
		x"6d",	--2684
		x"5c",	--2685
		x"6d",	--2686
		x"5c",	--2687
		x"6d",	--2688
		x"5c",	--2689
		x"6d",	--2690
		x"40",	--2691
		x"00",	--2692
		x"00",	--2693
		x"90",	--2694
		x"40",	--2695
		x"2c",	--2696
		x"40",	--2697
		x"ff",	--2698
		x"5c",	--2699
		x"6d",	--2700
		x"4f",	--2701
		x"53",	--2702
		x"90",	--2703
		x"40",	--2704
		x"2b",	--2705
		x"4a",	--2706
		x"00",	--2707
		x"4c",	--2708
		x"00",	--2709
		x"4d",	--2710
		x"00",	--2711
		x"41",	--2712
		x"41",	--2713
		x"41",	--2714
		x"90",	--2715
		x"00",	--2716
		x"24",	--2717
		x"50",	--2718
		x"ff",	--2719
		x"4d",	--2720
		x"00",	--2721
		x"40",	--2722
		x"00",	--2723
		x"00",	--2724
		x"4a",	--2725
		x"4b",	--2726
		x"5c",	--2727
		x"6d",	--2728
		x"5c",	--2729
		x"6d",	--2730
		x"5c",	--2731
		x"6d",	--2732
		x"5c",	--2733
		x"6d",	--2734
		x"5c",	--2735
		x"6d",	--2736
		x"5c",	--2737
		x"6d",	--2738
		x"5c",	--2739
		x"6d",	--2740
		x"4c",	--2741
		x"4d",	--2742
		x"d3",	--2743
		x"d0",	--2744
		x"40",	--2745
		x"4a",	--2746
		x"00",	--2747
		x"4b",	--2748
		x"00",	--2749
		x"41",	--2750
		x"41",	--2751
		x"41",	--2752
		x"93",	--2753
		x"23",	--2754
		x"43",	--2755
		x"00",	--2756
		x"41",	--2757
		x"41",	--2758
		x"41",	--2759
		x"93",	--2760
		x"24",	--2761
		x"4a",	--2762
		x"4b",	--2763
		x"f3",	--2764
		x"f0",	--2765
		x"00",	--2766
		x"93",	--2767
		x"20",	--2768
		x"93",	--2769
		x"24",	--2770
		x"43",	--2771
		x"00",	--2772
		x"3f",	--2773
		x"93",	--2774
		x"23",	--2775
		x"42",	--2776
		x"00",	--2777
		x"3f",	--2778
		x"43",	--2779
		x"00",	--2780
		x"3f",	--2781
		x"12",	--2782
		x"4f",	--2783
		x"93",	--2784
		x"28",	--2785
		x"4e",	--2786
		x"93",	--2787
		x"28",	--2788
		x"92",	--2789
		x"24",	--2790
		x"92",	--2791
		x"24",	--2792
		x"93",	--2793
		x"24",	--2794
		x"93",	--2795
		x"24",	--2796
		x"4f",	--2797
		x"00",	--2798
		x"9e",	--2799
		x"00",	--2800
		x"24",	--2801
		x"93",	--2802
		x"20",	--2803
		x"43",	--2804
		x"4e",	--2805
		x"41",	--2806
		x"41",	--2807
		x"93",	--2808
		x"24",	--2809
		x"93",	--2810
		x"00",	--2811
		x"23",	--2812
		x"43",	--2813
		x"4e",	--2814
		x"41",	--2815
		x"41",	--2816
		x"93",	--2817
		x"00",	--2818
		x"27",	--2819
		x"43",	--2820
		x"3f",	--2821
		x"4f",	--2822
		x"00",	--2823
		x"4e",	--2824
		x"00",	--2825
		x"9b",	--2826
		x"3b",	--2827
		x"9c",	--2828
		x"38",	--2829
		x"4f",	--2830
		x"00",	--2831
		x"4f",	--2832
		x"00",	--2833
		x"4e",	--2834
		x"00",	--2835
		x"4e",	--2836
		x"00",	--2837
		x"9f",	--2838
		x"2b",	--2839
		x"9e",	--2840
		x"28",	--2841
		x"9b",	--2842
		x"2b",	--2843
		x"9e",	--2844
		x"28",	--2845
		x"9f",	--2846
		x"28",	--2847
		x"9c",	--2848
		x"28",	--2849
		x"43",	--2850
		x"3f",	--2851
		x"93",	--2852
		x"23",	--2853
		x"43",	--2854
		x"3f",	--2855
		x"92",	--2856
		x"23",	--2857
		x"4e",	--2858
		x"00",	--2859
		x"4f",	--2860
		x"00",	--2861
		x"8f",	--2862
		x"3f",	--2863
		x"43",	--2864
		x"93",	--2865
		x"34",	--2866
		x"40",	--2867
		x"00",	--2868
		x"e3",	--2869
		x"53",	--2870
		x"93",	--2871
		x"34",	--2872
		x"e3",	--2873
		x"e3",	--2874
		x"53",	--2875
		x"12",	--2876
		x"12",	--2877
		x"f6",	--2878
		x"41",	--2879
		x"b3",	--2880
		x"24",	--2881
		x"e3",	--2882
		x"53",	--2883
		x"b3",	--2884
		x"24",	--2885
		x"e3",	--2886
		x"53",	--2887
		x"41",	--2888
		x"12",	--2889
		x"f6",	--2890
		x"4e",	--2891
		x"41",	--2892
		x"12",	--2893
		x"43",	--2894
		x"93",	--2895
		x"34",	--2896
		x"40",	--2897
		x"00",	--2898
		x"e3",	--2899
		x"e3",	--2900
		x"53",	--2901
		x"63",	--2902
		x"93",	--2903
		x"34",	--2904
		x"e3",	--2905
		x"e3",	--2906
		x"e3",	--2907
		x"53",	--2908
		x"63",	--2909
		x"12",	--2910
		x"f7",	--2911
		x"b3",	--2912
		x"24",	--2913
		x"e3",	--2914
		x"e3",	--2915
		x"53",	--2916
		x"63",	--2917
		x"b3",	--2918
		x"24",	--2919
		x"e3",	--2920
		x"e3",	--2921
		x"53",	--2922
		x"63",	--2923
		x"41",	--2924
		x"41",	--2925
		x"12",	--2926
		x"f6",	--2927
		x"4c",	--2928
		x"4d",	--2929
		x"41",	--2930
		x"40",	--2931
		x"00",	--2932
		x"4e",	--2933
		x"43",	--2934
		x"5f",	--2935
		x"6e",	--2936
		x"9d",	--2937
		x"28",	--2938
		x"8d",	--2939
		x"d3",	--2940
		x"83",	--2941
		x"23",	--2942
		x"41",	--2943
		x"12",	--2944
		x"f6",	--2945
		x"4e",	--2946
		x"41",	--2947
		x"12",	--2948
		x"12",	--2949
		x"12",	--2950
		x"40",	--2951
		x"00",	--2952
		x"4c",	--2953
		x"4d",	--2954
		x"43",	--2955
		x"43",	--2956
		x"5e",	--2957
		x"6f",	--2958
		x"6c",	--2959
		x"6d",	--2960
		x"9b",	--2961
		x"28",	--2962
		x"20",	--2963
		x"9a",	--2964
		x"28",	--2965
		x"8a",	--2966
		x"7b",	--2967
		x"d3",	--2968
		x"83",	--2969
		x"23",	--2970
		x"41",	--2971
		x"41",	--2972
		x"41",	--2973
		x"41",	--2974
		x"12",	--2975
		x"f7",	--2976
		x"4c",	--2977
		x"4d",	--2978
		x"41",	--2979
		x"13",	--2980
		x"d0",	--2981
		x"00",	--2982
		x"3f",	--2983
		x"6f",	--2984
		x"72",	--2985
		x"63",	--2986
		x"20",	--2987
		x"73",	--2988
		x"67",	--2989
		x"3a",	--2990
		x"0a",	--2991
		x"09",	--2992
		x"63",	--2993
		x"4c",	--2994
		x"46",	--2995
		x"20",	--2996
		x"49",	--2997
		x"48",	--2998
		x"0d",	--2999
		x"00",	--3000
		x"6f",	--3001
		x"65",	--3002
		x"68",	--3003
		x"6e",	--3004
		x"20",	--3005
		x"65",	--3006
		x"74",	--3007
		x"74",	--3008
		x"72",	--3009
		x"69",	--3010
		x"6c",	--3011
		x"20",	--3012
		x"72",	--3013
		x"6e",	--3014
		x"0d",	--3015
		x"00",	--3016
		x"0a",	--3017
		x"3d",	--3018
		x"3d",	--3019
		x"3d",	--3020
		x"6f",	--3021
		x"65",	--3022
		x"4d",	--3023
		x"50",	--3024
		x"33",	--3025
		x"20",	--3026
		x"6e",	--3027
		x"61",	--3028
		x"74",	--3029
		x"6f",	--3030
		x"20",	--3031
		x"3d",	--3032
		x"3d",	--3033
		x"3d",	--3034
		x"0a",	--3035
		x"0d",	--3036
		x"53",	--3037
		x"6d",	--3038
		x"6c",	--3039
		x"20",	--3040
		x"69",	--3041
		x"65",	--3042
		x"45",	--3043
		x"69",	--3044
		x"6f",	--3045
		x"20",	--3046
		x"65",	--3047
		x"64",	--3048
		x"0d",	--3049
		x"00",	--3050
		x"0a",	--3051
		x"41",	--3052
		x"44",	--3053
		x"25",	--3054
		x"0d",	--3055
		x"00",	--3056
		x"0a",	--3057
		x"65",	--3058
		x"74",	--3059
		x"25",	--3060
		x"0d",	--3061
		x"00",	--3062
		x"20",	--3063
		x"0d",	--3064
		x"00",	--3065
		x"25",	--3066
		x"0d",	--3067
		x"00",	--3068
		x"20",	--3069
		x"00",	--3070
		x"63",	--3071
		x"77",	--3072
		x"69",	--3073
		x"65",	--3074
		x"0d",	--3075
		x"63",	--3076
		x"72",	--3077
		x"65",	--3078
		x"74",	--3079
		x"75",	--3080
		x"61",	--3081
		x"65",	--3082
		x"0d",	--3083
		x"00",	--3084
		x"25",	--3085
		x"20",	--3086
		x"45",	--3087
		x"49",	--3088
		x"54",	--3089
		x"52",	--3090
		x"56",	--3091
		x"4c",	--3092
		x"45",	--3093
		x"0a",	--3094
		x"53",	--3095
		x"6d",	--3096
		x"74",	--3097
		x"69",	--3098
		x"67",	--3099
		x"77",	--3100
		x"6e",	--3101
		x"20",	--3102
		x"65",	--3103
		x"72",	--3104
		x"62",	--3105
		x"79",	--3106
		x"77",	--3107
		x"6f",	--3108
		x"67",	--3109
		x"0a",	--3110
		x"72",	--3111
		x"25",	--3112
		x"20",	--3113
		x"3d",	--3114
		x"64",	--3115
		x"0a",	--3116
		x"72",	--3117
		x"61",	--3118
		x"0a",	--3119
		x"00",	--3120
		x"25",	--3121
		x"20",	--3122
		x"45",	--3123
		x"49",	--3124
		x"54",	--3125
		x"52",	--3126
		x"0a",	--3127
		x"25",	--3128
		x"20",	--3129
		x"73",	--3130
		x"6e",	--3131
		x"74",	--3132
		x"61",	--3133
		x"6e",	--3134
		x"6d",	--3135
		x"65",	--3136
		x"0d",	--3137
		x"00",	--3138
		x"63",	--3139
		x"20",	--3140
		x"6f",	--3141
		x"73",	--3142
		x"63",	--3143
		x"20",	--3144
		x"6f",	--3145
		x"6d",	--3146
		x"6e",	--3147
		x"0d",	--3148
		x"00",	--3149
		x"e8",	--3150
		x"e8",	--3151
		x"e8",	--3152
		x"e8",	--3153
		x"e8",	--3154
		x"e8",	--3155
		x"e8",	--3156
		x"e8",	--3157
		x"e8",	--3158
		x"e8",	--3159
		x"e8",	--3160
		x"e8",	--3161
		x"e8",	--3162
		x"e8",	--3163
		x"e8",	--3164
		x"e8",	--3165
		x"e8",	--3166
		x"e8",	--3167
		x"e8",	--3168
		x"e8",	--3169
		x"e8",	--3170
		x"e8",	--3171
		x"e8",	--3172
		x"e8",	--3173
		x"e8",	--3174
		x"e8",	--3175
		x"e8",	--3176
		x"e8",	--3177
		x"e8",	--3178
		x"e8",	--3179
		x"e8",	--3180
		x"e8",	--3181
		x"e8",	--3182
		x"e8",	--3183
		x"e8",	--3184
		x"e8",	--3185
		x"e8",	--3186
		x"e8",	--3187
		x"e8",	--3188
		x"e8",	--3189
		x"e8",	--3190
		x"e8",	--3191
		x"e8",	--3192
		x"e8",	--3193
		x"e8",	--3194
		x"e8",	--3195
		x"e8",	--3196
		x"e8",	--3197
		x"e8",	--3198
		x"e8",	--3199
		x"e8",	--3200
		x"e8",	--3201
		x"e8",	--3202
		x"e8",	--3203
		x"e8",	--3204
		x"e8",	--3205
		x"e8",	--3206
		x"e8",	--3207
		x"e8",	--3208
		x"e8",	--3209
		x"e8",	--3210
		x"e8",	--3211
		x"e8",	--3212
		x"e8",	--3213
		x"e8",	--3214
		x"e8",	--3215
		x"e8",	--3216
		x"e8",	--3217
		x"e8",	--3218
		x"e8",	--3219
		x"e8",	--3220
		x"e8",	--3221
		x"e8",	--3222
		x"e8",	--3223
		x"e8",	--3224
		x"e8",	--3225
		x"e8",	--3226
		x"e8",	--3227
		x"e8",	--3228
		x"e8",	--3229
		x"e8",	--3230
		x"e8",	--3231
		x"e8",	--3232
		x"e8",	--3233
		x"31",	--3234
		x"33",	--3235
		x"35",	--3236
		x"37",	--3237
		x"39",	--3238
		x"62",	--3239
		x"64",	--3240
		x"66",	--3241
		x"00",	--3242
		x"00",	--3243
		x"00",	--3244
		x"00",	--3245
		x"00",	--3246
		x"01",	--3247
		x"02",	--3248
		x"03",	--3249
		x"03",	--3250
		x"04",	--3251
		x"04",	--3252
		x"04",	--3253
		x"04",	--3254
		x"05",	--3255
		x"05",	--3256
		x"05",	--3257
		x"05",	--3258
		x"05",	--3259
		x"05",	--3260
		x"05",	--3261
		x"05",	--3262
		x"06",	--3263
		x"06",	--3264
		x"06",	--3265
		x"06",	--3266
		x"06",	--3267
		x"06",	--3268
		x"06",	--3269
		x"06",	--3270
		x"06",	--3271
		x"06",	--3272
		x"06",	--3273
		x"06",	--3274
		x"06",	--3275
		x"06",	--3276
		x"06",	--3277
		x"06",	--3278
		x"07",	--3279
		x"07",	--3280
		x"07",	--3281
		x"07",	--3282
		x"07",	--3283
		x"07",	--3284
		x"07",	--3285
		x"07",	--3286
		x"07",	--3287
		x"07",	--3288
		x"07",	--3289
		x"07",	--3290
		x"07",	--3291
		x"07",	--3292
		x"07",	--3293
		x"07",	--3294
		x"07",	--3295
		x"07",	--3296
		x"07",	--3297
		x"07",	--3298
		x"07",	--3299
		x"07",	--3300
		x"07",	--3301
		x"07",	--3302
		x"07",	--3303
		x"07",	--3304
		x"07",	--3305
		x"07",	--3306
		x"07",	--3307
		x"07",	--3308
		x"07",	--3309
		x"07",	--3310
		x"08",	--3311
		x"08",	--3312
		x"08",	--3313
		x"08",	--3314
		x"08",	--3315
		x"08",	--3316
		x"08",	--3317
		x"08",	--3318
		x"08",	--3319
		x"08",	--3320
		x"08",	--3321
		x"08",	--3322
		x"08",	--3323
		x"08",	--3324
		x"08",	--3325
		x"08",	--3326
		x"08",	--3327
		x"08",	--3328
		x"08",	--3329
		x"08",	--3330
		x"08",	--3331
		x"08",	--3332
		x"08",	--3333
		x"08",	--3334
		x"08",	--3335
		x"08",	--3336
		x"08",	--3337
		x"08",	--3338
		x"08",	--3339
		x"08",	--3340
		x"08",	--3341
		x"08",	--3342
		x"08",	--3343
		x"08",	--3344
		x"08",	--3345
		x"08",	--3346
		x"08",	--3347
		x"08",	--3348
		x"08",	--3349
		x"08",	--3350
		x"08",	--3351
		x"08",	--3352
		x"08",	--3353
		x"08",	--3354
		x"08",	--3355
		x"08",	--3356
		x"08",	--3357
		x"08",	--3358
		x"08",	--3359
		x"08",	--3360
		x"08",	--3361
		x"08",	--3362
		x"08",	--3363
		x"08",	--3364
		x"08",	--3365
		x"08",	--3366
		x"08",	--3367
		x"08",	--3368
		x"08",	--3369
		x"08",	--3370
		x"08",	--3371
		x"08",	--3372
		x"08",	--3373
		x"08",	--3374
		x"ff",	--3375
		x"ff",	--3376
		x"ff",	--3377
		x"ff",	--3378
		x"ff",	--3379
		x"ff",	--3380
		x"ff",	--3381
		x"ff",	--3382
		x"ff",	--3383
		x"ff",	--3384
		x"ff",	--3385
		x"ff",	--3386
		x"ff",	--3387
		x"ff",	--3388
		x"ff",	--3389
		x"ff",	--3390
		x"ff",	--3391
		x"ff",	--3392
		x"ff",	--3393
		x"ff",	--3394
		x"ff",	--3395
		x"ff",	--3396
		x"ff",	--3397
		x"ff",	--3398
		x"ff",	--3399
		x"ff",	--3400
		x"ff",	--3401
		x"ff",	--3402
		x"ff",	--3403
		x"ff",	--3404
		x"ff",	--3405
		x"ff",	--3406
		x"ff",	--3407
		x"ff",	--3408
		x"ff",	--3409
		x"ff",	--3410
		x"ff",	--3411
		x"ff",	--3412
		x"ff",	--3413
		x"ff",	--3414
		x"ff",	--3415
		x"ff",	--3416
		x"ff",	--3417
		x"ff",	--3418
		x"ff",	--3419
		x"ff",	--3420
		x"ff",	--3421
		x"ff",	--3422
		x"ff",	--3423
		x"ff",	--3424
		x"ff",	--3425
		x"ff",	--3426
		x"ff",	--3427
		x"ff",	--3428
		x"ff",	--3429
		x"ff",	--3430
		x"ff",	--3431
		x"ff",	--3432
		x"ff",	--3433
		x"ff",	--3434
		x"ff",	--3435
		x"ff",	--3436
		x"ff",	--3437
		x"ff",	--3438
		x"ff",	--3439
		x"ff",	--3440
		x"ff",	--3441
		x"ff",	--3442
		x"ff",	--3443
		x"ff",	--3444
		x"ff",	--3445
		x"ff",	--3446
		x"ff",	--3447
		x"ff",	--3448
		x"ff",	--3449
		x"ff",	--3450
		x"ff",	--3451
		x"ff",	--3452
		x"ff",	--3453
		x"ff",	--3454
		x"ff",	--3455
		x"ff",	--3456
		x"ff",	--3457
		x"ff",	--3458
		x"ff",	--3459
		x"ff",	--3460
		x"ff",	--3461
		x"ff",	--3462
		x"ff",	--3463
		x"ff",	--3464
		x"ff",	--3465
		x"ff",	--3466
		x"ff",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"e8",	--4087
		x"e1",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
