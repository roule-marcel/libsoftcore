library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"34",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"10",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"34",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"a0",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"24",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"34",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"10",	--29
		x"f9",	--30
		x"31",	--31
		x"62",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"3c",	--44
		x"b0",	--45
		x"78",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"90",	--50
		x"b0",	--51
		x"00",	--52
		x"21",	--53
		x"3d",	--54
		x"ad",	--55
		x"3e",	--56
		x"ea",	--57
		x"7f",	--58
		x"69",	--59
		x"b0",	--60
		x"a8",	--61
		x"3d",	--62
		x"be",	--63
		x"3e",	--64
		x"28",	--65
		x"7f",	--66
		x"77",	--67
		x"b0",	--68
		x"a8",	--69
		x"3d",	--70
		x"c4",	--71
		x"3e",	--72
		x"9c",	--73
		x"7f",	--74
		x"72",	--75
		x"b0",	--76
		x"a8",	--77
		x"3d",	--78
		x"c9",	--79
		x"3e",	--80
		x"18",	--81
		x"7f",	--82
		x"61",	--83
		x"b0",	--84
		x"a8",	--85
		x"3d",	--86
		x"d0",	--87
		x"3e",	--88
		x"a0",	--89
		x"7f",	--90
		x"70",	--91
		x"b0",	--92
		x"a8",	--93
		x"3d",	--94
		x"d4",	--95
		x"3e",	--96
		x"e0",	--97
		x"7f",	--98
		x"65",	--99
		x"b0",	--100
		x"a8",	--101
		x"3d",	--102
		x"dc",	--103
		x"3e",	--104
		x"be",	--105
		x"7f",	--106
		x"73",	--107
		x"b0",	--108
		x"a8",	--109
		x"3d",	--110
		x"ed",	--111
		x"3e",	--112
		x"e6",	--113
		x"7f",	--114
		x"63",	--115
		x"b0",	--116
		x"a8",	--117
		x"3d",	--118
		x"01",	--119
		x"3e",	--120
		x"a4",	--121
		x"7f",	--122
		x"64",	--123
		x"b0",	--124
		x"a8",	--125
		x"3d",	--126
		x"07",	--127
		x"3e",	--128
		x"f4",	--129
		x"7f",	--130
		x"62",	--131
		x"b0",	--132
		x"a8",	--133
		x"0e",	--134
		x"0f",	--135
		x"b0",	--136
		x"3e",	--137
		x"2c",	--138
		x"3d",	--139
		x"20",	--140
		x"3e",	--141
		x"80",	--142
		x"0f",	--143
		x"3f",	--144
		x"12",	--145
		x"b0",	--146
		x"46",	--147
		x"0f",	--148
		x"3f",	--149
		x"12",	--150
		x"b0",	--151
		x"8e",	--152
		x"2c",	--153
		x"3d",	--154
		x"20",	--155
		x"3e",	--156
		x"88",	--157
		x"0f",	--158
		x"3f",	--159
		x"b0",	--160
		x"46",	--161
		x"0f",	--162
		x"3f",	--163
		x"b0",	--164
		x"8e",	--165
		x"0e",	--166
		x"3e",	--167
		x"0f",	--168
		x"3f",	--169
		x"12",	--170
		x"b0",	--171
		x"96",	--172
		x"3e",	--173
		x"98",	--174
		x"0f",	--175
		x"3f",	--176
		x"06",	--177
		x"b0",	--178
		x"e2",	--179
		x"3e",	--180
		x"9c",	--181
		x"0f",	--182
		x"2f",	--183
		x"b0",	--184
		x"e2",	--185
		x"0e",	--186
		x"2e",	--187
		x"0f",	--188
		x"3f",	--189
		x"06",	--190
		x"b0",	--191
		x"cc",	--192
		x"0e",	--193
		x"3e",	--194
		x"0f",	--195
		x"3f",	--196
		x"12",	--197
		x"b0",	--198
		x"d6",	--199
		x"b0",	--200
		x"ba",	--201
		x"3e",	--202
		x"a0",	--203
		x"0f",	--204
		x"2f",	--205
		x"b0",	--206
		x"fa",	--207
		x"0f",	--208
		x"2f",	--209
		x"b0",	--210
		x"12",	--211
		x"3d",	--212
		x"64",	--213
		x"3e",	--214
		x"2a",	--215
		x"0f",	--216
		x"2f",	--217
		x"b0",	--218
		x"0e",	--219
		x"3e",	--220
		x"b0",	--221
		x"0f",	--222
		x"b0",	--223
		x"74",	--224
		x"0f",	--225
		x"b0",	--226
		x"9e",	--227
		x"30",	--228
		x"a0",	--229
		x"03",	--230
		x"03",	--231
		x"03",	--232
		x"30",	--233
		x"d1",	--234
		x"30",	--235
		x"17",	--236
		x"30",	--237
		x"1d",	--238
		x"30",	--239
		x"52",	--240
		x"3c",	--241
		x"32",	--242
		x"0d",	--243
		x"3d",	--244
		x"16",	--245
		x"0e",	--246
		x"3e",	--247
		x"22",	--248
		x"0f",	--249
		x"3f",	--250
		x"80",	--251
		x"b0",	--252
		x"ae",	--253
		x"31",	--254
		x"10",	--255
		x"30",	--256
		x"a0",	--257
		x"03",	--258
		x"03",	--259
		x"03",	--260
		x"30",	--261
		x"d1",	--262
		x"30",	--263
		x"17",	--264
		x"30",	--265
		x"1d",	--266
		x"30",	--267
		x"52",	--268
		x"3c",	--269
		x"32",	--270
		x"0d",	--271
		x"3d",	--272
		x"14",	--273
		x"0e",	--274
		x"3e",	--275
		x"18",	--276
		x"0f",	--277
		x"3f",	--278
		x"54",	--279
		x"b0",	--280
		x"ae",	--281
		x"31",	--282
		x"10",	--283
		x"0e",	--284
		x"3e",	--285
		x"44",	--286
		x"0f",	--287
		x"3f",	--288
		x"70",	--289
		x"b0",	--290
		x"b4",	--291
		x"b0",	--292
		x"8c",	--293
		x"f2",	--294
		x"80",	--295
		x"19",	--296
		x"32",	--297
		x"0b",	--298
		x"0a",	--299
		x"05",	--300
		x"1b",	--301
		x"03",	--302
		x"2b",	--303
		x"01",	--304
		x"0b",	--305
		x"b0",	--306
		x"5a",	--307
		x"0f",	--308
		x"fc",	--309
		x"b0",	--310
		x"82",	--311
		x"0b",	--312
		x"3e",	--313
		x"7f",	--314
		x"0d",	--315
		x"06",	--316
		x"7f",	--317
		x"1b",	--318
		x"ed",	--319
		x"7f",	--320
		x"1c",	--321
		x"12",	--322
		x"30",	--323
		x"12",	--324
		x"b0",	--325
		x"00",	--326
		x"21",	--327
		x"3f",	--328
		x"1c",	--329
		x"0f",	--330
		x"0a",	--331
		x"ca",	--332
		x"00",	--333
		x"0e",	--334
		x"5f",	--335
		x"1c",	--336
		x"b0",	--337
		x"dc",	--338
		x"0a",	--339
		x"dd",	--340
		x"0a",	--341
		x"db",	--342
		x"3a",	--343
		x"30",	--344
		x"15",	--345
		x"b0",	--346
		x"00",	--347
		x"21",	--348
		x"d4",	--349
		x"3a",	--350
		x"28",	--351
		x"d1",	--352
		x"82",	--353
		x"14",	--354
		x"0c",	--355
		x"4e",	--356
		x"8e",	--357
		x"0e",	--358
		x"30",	--359
		x"19",	--360
		x"81",	--361
		x"a0",	--362
		x"b0",	--363
		x"00",	--364
		x"21",	--365
		x"1f",	--366
		x"9c",	--367
		x"3e",	--368
		x"1c",	--369
		x"0e",	--370
		x"0e",	--371
		x"ce",	--372
		x"00",	--373
		x"1a",	--374
		x"ba",	--375
		x"1b",	--376
		x"04",	--377
		x"7f",	--378
		x"5b",	--379
		x"b5",	--380
		x"b1",	--381
		x"2b",	--382
		x"b2",	--383
		x"7f",	--384
		x"42",	--385
		x"17",	--386
		x"7f",	--387
		x"43",	--388
		x"04",	--389
		x"7f",	--390
		x"41",	--391
		x"a8",	--392
		x"07",	--393
		x"7f",	--394
		x"43",	--395
		x"16",	--396
		x"7f",	--397
		x"44",	--398
		x"a1",	--399
		x"1b",	--400
		x"30",	--401
		x"1c",	--402
		x"b0",	--403
		x"00",	--404
		x"21",	--405
		x"b0",	--406
		x"46",	--407
		x"0b",	--408
		x"98",	--409
		x"30",	--410
		x"21",	--411
		x"b0",	--412
		x"00",	--413
		x"21",	--414
		x"b0",	--415
		x"6e",	--416
		x"0b",	--417
		x"8f",	--418
		x"30",	--419
		x"28",	--420
		x"b0",	--421
		x"00",	--422
		x"21",	--423
		x"b0",	--424
		x"96",	--425
		x"0b",	--426
		x"86",	--427
		x"30",	--428
		x"30",	--429
		x"b0",	--430
		x"00",	--431
		x"21",	--432
		x"b0",	--433
		x"be",	--434
		x"0b",	--435
		x"7d",	--436
		x"30",	--437
		x"7e",	--438
		x"0b",	--439
		x"0b",	--440
		x"0e",	--441
		x"1f",	--442
		x"24",	--443
		x"b0",	--444
		x"84",	--445
		x"0f",	--446
		x"30",	--447
		x"86",	--448
		x"b0",	--449
		x"00",	--450
		x"21",	--451
		x"1b",	--452
		x"3b",	--453
		x"05",	--454
		x"f1",	--455
		x"30",	--456
		x"8a",	--457
		x"b0",	--458
		x"00",	--459
		x"21",	--460
		x"3b",	--461
		x"30",	--462
		x"82",	--463
		x"24",	--464
		x"30",	--465
		x"0b",	--466
		x"21",	--467
		x"0b",	--468
		x"81",	--469
		x"00",	--470
		x"1f",	--471
		x"14",	--472
		x"b2",	--473
		x"00",	--474
		x"25",	--475
		x"92",	--476
		x"10",	--477
		x"0e",	--478
		x"1f",	--479
		x"02",	--480
		x"b0",	--481
		x"f8",	--482
		x"0d",	--483
		x"0e",	--484
		x"1f",	--485
		x"00",	--486
		x"b0",	--487
		x"0e",	--488
		x"0f",	--489
		x"21",	--490
		x"3b",	--491
		x"30",	--492
		x"82",	--493
		x"10",	--494
		x"0a",	--495
		x"82",	--496
		x"10",	--497
		x"1f",	--498
		x"00",	--499
		x"b0",	--500
		x"36",	--501
		x"0f",	--502
		x"21",	--503
		x"3b",	--504
		x"30",	--505
		x"0f",	--506
		x"b0",	--507
		x"6e",	--508
		x"0f",	--509
		x"21",	--510
		x"3b",	--511
		x"30",	--512
		x"0e",	--513
		x"3f",	--514
		x"6e",	--515
		x"b0",	--516
		x"ca",	--517
		x"82",	--518
		x"00",	--519
		x"d3",	--520
		x"82",	--521
		x"26",	--522
		x"30",	--523
		x"0b",	--524
		x"0a",	--525
		x"21",	--526
		x"0a",	--527
		x"0b",	--528
		x"2f",	--529
		x"1b",	--530
		x"0e",	--531
		x"1f",	--532
		x"02",	--533
		x"b0",	--534
		x"f8",	--535
		x"0d",	--536
		x"2a",	--537
		x"18",	--538
		x"0e",	--539
		x"1f",	--540
		x"04",	--541
		x"81",	--542
		x"02",	--543
		x"b0",	--544
		x"f8",	--545
		x"0e",	--546
		x"1d",	--547
		x"02",	--548
		x"1f",	--549
		x"26",	--550
		x"b0",	--551
		x"0e",	--552
		x"0f",	--553
		x"21",	--554
		x"3a",	--555
		x"3b",	--556
		x"30",	--557
		x"3d",	--558
		x"64",	--559
		x"3e",	--560
		x"2a",	--561
		x"f2",	--562
		x"3e",	--563
		x"2a",	--564
		x"ef",	--565
		x"0e",	--566
		x"1f",	--567
		x"2a",	--568
		x"b0",	--569
		x"42",	--570
		x"0e",	--571
		x"1f",	--572
		x"28",	--573
		x"b0",	--574
		x"42",	--575
		x"30",	--576
		x"8d",	--577
		x"b0",	--578
		x"00",	--579
		x"21",	--580
		x"30",	--581
		x"b2",	--582
		x"02",	--583
		x"09",	--584
		x"1f",	--585
		x"2a",	--586
		x"b0",	--587
		x"fe",	--588
		x"1f",	--589
		x"28",	--590
		x"b0",	--591
		x"fe",	--592
		x"30",	--593
		x"0e",	--594
		x"3f",	--595
		x"6c",	--596
		x"b0",	--597
		x"ca",	--598
		x"82",	--599
		x"02",	--600
		x"ef",	--601
		x"82",	--602
		x"2a",	--603
		x"82",	--604
		x"28",	--605
		x"30",	--606
		x"0b",	--607
		x"0a",	--608
		x"21",	--609
		x"0b",	--610
		x"3f",	--611
		x"03",	--612
		x"30",	--613
		x"23",	--614
		x"0e",	--615
		x"1f",	--616
		x"02",	--617
		x"b0",	--618
		x"c6",	--619
		x"0a",	--620
		x"0e",	--621
		x"1f",	--622
		x"04",	--623
		x"b0",	--624
		x"c6",	--625
		x"0b",	--626
		x"0f",	--627
		x"0a",	--628
		x"30",	--629
		x"c0",	--630
		x"b0",	--631
		x"00",	--632
		x"31",	--633
		x"06",	--634
		x"0e",	--635
		x"1f",	--636
		x"2a",	--637
		x"b0",	--638
		x"42",	--639
		x"0e",	--640
		x"1f",	--641
		x"28",	--642
		x"b0",	--643
		x"42",	--644
		x"0f",	--645
		x"21",	--646
		x"3a",	--647
		x"3b",	--648
		x"30",	--649
		x"0e",	--650
		x"1f",	--651
		x"06",	--652
		x"b0",	--653
		x"f8",	--654
		x"1d",	--655
		x"0e",	--656
		x"1f",	--657
		x"02",	--658
		x"b0",	--659
		x"0e",	--660
		x"d1",	--661
		x"30",	--662
		x"94",	--663
		x"b0",	--664
		x"00",	--665
		x"a1",	--666
		x"00",	--667
		x"30",	--668
		x"a5",	--669
		x"b0",	--670
		x"00",	--671
		x"21",	--672
		x"3f",	--673
		x"e3",	--674
		x"3e",	--675
		x"9c",	--676
		x"1f",	--677
		x"2a",	--678
		x"b0",	--679
		x"42",	--680
		x"3e",	--681
		x"64",	--682
		x"1f",	--683
		x"28",	--684
		x"b0",	--685
		x"42",	--686
		x"1d",	--687
		x"3e",	--688
		x"c8",	--689
		x"1f",	--690
		x"02",	--691
		x"b0",	--692
		x"0e",	--693
		x"30",	--694
		x"3e",	--695
		x"64",	--696
		x"1f",	--697
		x"2a",	--698
		x"b0",	--699
		x"42",	--700
		x"3e",	--701
		x"9c",	--702
		x"1f",	--703
		x"28",	--704
		x"b0",	--705
		x"42",	--706
		x"1d",	--707
		x"3e",	--708
		x"c8",	--709
		x"1f",	--710
		x"02",	--711
		x"b0",	--712
		x"0e",	--713
		x"30",	--714
		x"3e",	--715
		x"c4",	--716
		x"1f",	--717
		x"2a",	--718
		x"b0",	--719
		x"42",	--720
		x"3e",	--721
		x"c4",	--722
		x"1f",	--723
		x"28",	--724
		x"b0",	--725
		x"42",	--726
		x"1d",	--727
		x"3e",	--728
		x"c8",	--729
		x"1f",	--730
		x"02",	--731
		x"b0",	--732
		x"0e",	--733
		x"30",	--734
		x"3e",	--735
		x"3c",	--736
		x"1f",	--737
		x"2a",	--738
		x"b0",	--739
		x"42",	--740
		x"3e",	--741
		x"3c",	--742
		x"1f",	--743
		x"28",	--744
		x"b0",	--745
		x"42",	--746
		x"1d",	--747
		x"3e",	--748
		x"c8",	--749
		x"1f",	--750
		x"02",	--751
		x"b0",	--752
		x"0e",	--753
		x"30",	--754
		x"30",	--755
		x"c8",	--756
		x"b0",	--757
		x"00",	--758
		x"21",	--759
		x"0f",	--760
		x"30",	--761
		x"b2",	--762
		x"00",	--763
		x"92",	--764
		x"b2",	--765
		x"30",	--766
		x"94",	--767
		x"b2",	--768
		x"41",	--769
		x"96",	--770
		x"30",	--771
		x"de",	--772
		x"b0",	--773
		x"00",	--774
		x"92",	--775
		x"90",	--776
		x"b1",	--777
		x"fc",	--778
		x"00",	--779
		x"b0",	--780
		x"00",	--781
		x"21",	--782
		x"0f",	--783
		x"30",	--784
		x"0b",	--785
		x"0a",	--786
		x"09",	--787
		x"09",	--788
		x"1f",	--789
		x"22",	--790
		x"b0",	--791
		x"ea",	--792
		x"0a",	--793
		x"0b",	--794
		x"1e",	--795
		x"24",	--796
		x"1f",	--797
		x"26",	--798
		x"b0",	--799
		x"84",	--800
		x"89",	--801
		x"24",	--802
		x"89",	--803
		x"26",	--804
		x"0d",	--805
		x"0e",	--806
		x"0f",	--807
		x"b0",	--808
		x"0a",	--809
		x"0c",	--810
		x"3d",	--811
		x"00",	--812
		x"b0",	--813
		x"84",	--814
		x"0a",	--815
		x"0b",	--816
		x"3c",	--817
		x"66",	--818
		x"3d",	--819
		x"66",	--820
		x"b0",	--821
		x"94",	--822
		x"0f",	--823
		x"01",	--824
		x"18",	--825
		x"3c",	--826
		x"cd",	--827
		x"3d",	--828
		x"cc",	--829
		x"0e",	--830
		x"0f",	--831
		x"b0",	--832
		x"34",	--833
		x"0f",	--834
		x"04",	--835
		x"3a",	--836
		x"cd",	--837
		x"3b",	--838
		x"cc",	--839
		x"0d",	--840
		x"0e",	--841
		x"1f",	--842
		x"20",	--843
		x"b0",	--844
		x"e2",	--845
		x"39",	--846
		x"3a",	--847
		x"3b",	--848
		x"30",	--849
		x"3a",	--850
		x"66",	--851
		x"3b",	--852
		x"66",	--853
		x"f1",	--854
		x"0b",	--855
		x"0a",	--856
		x"0b",	--857
		x"0a",	--858
		x"8f",	--859
		x"20",	--860
		x"8f",	--861
		x"22",	--862
		x"11",	--863
		x"16",	--864
		x"11",	--865
		x"16",	--866
		x"11",	--867
		x"16",	--868
		x"11",	--869
		x"16",	--870
		x"11",	--871
		x"16",	--872
		x"11",	--873
		x"16",	--874
		x"1d",	--875
		x"12",	--876
		x"1e",	--877
		x"14",	--878
		x"b0",	--879
		x"70",	--880
		x"31",	--881
		x"0c",	--882
		x"8b",	--883
		x"28",	--884
		x"0e",	--885
		x"3f",	--886
		x"22",	--887
		x"b0",	--888
		x"ca",	--889
		x"8b",	--890
		x"2a",	--891
		x"3a",	--892
		x"3b",	--893
		x"30",	--894
		x"0b",	--895
		x"0b",	--896
		x"1f",	--897
		x"22",	--898
		x"b0",	--899
		x"ea",	--900
		x"8b",	--901
		x"24",	--902
		x"8b",	--903
		x"26",	--904
		x"0d",	--905
		x"1e",	--906
		x"28",	--907
		x"1f",	--908
		x"2a",	--909
		x"b0",	--910
		x"0e",	--911
		x"3b",	--912
		x"30",	--913
		x"0b",	--914
		x"0b",	--915
		x"0d",	--916
		x"3e",	--917
		x"00",	--918
		x"1f",	--919
		x"20",	--920
		x"b0",	--921
		x"e2",	--922
		x"1f",	--923
		x"2a",	--924
		x"b0",	--925
		x"36",	--926
		x"3b",	--927
		x"30",	--928
		x"0b",	--929
		x"0b",	--930
		x"0d",	--931
		x"8d",	--932
		x"8d",	--933
		x"8d",	--934
		x"8d",	--935
		x"0f",	--936
		x"b0",	--937
		x"84",	--938
		x"0d",	--939
		x"0e",	--940
		x"0f",	--941
		x"b0",	--942
		x"f6",	--943
		x"3b",	--944
		x"30",	--945
		x"0b",	--946
		x"0a",	--947
		x"0a",	--948
		x"3b",	--949
		x"00",	--950
		x"0d",	--951
		x"0e",	--952
		x"1f",	--953
		x"6e",	--954
		x"b0",	--955
		x"e2",	--956
		x"0d",	--957
		x"0e",	--958
		x"1f",	--959
		x"6c",	--960
		x"b0",	--961
		x"e2",	--962
		x"30",	--963
		x"15",	--964
		x"b0",	--965
		x"00",	--966
		x"21",	--967
		x"3a",	--968
		x"3b",	--969
		x"30",	--970
		x"82",	--971
		x"6e",	--972
		x"82",	--973
		x"6c",	--974
		x"30",	--975
		x"0b",	--976
		x"0a",	--977
		x"21",	--978
		x"0a",	--979
		x"0b",	--980
		x"b2",	--981
		x"04",	--982
		x"4e",	--983
		x"3a",	--984
		x"03",	--985
		x"53",	--986
		x"3e",	--987
		x"0e",	--988
		x"1f",	--989
		x"02",	--990
		x"b0",	--991
		x"f8",	--992
		x"0a",	--993
		x"0e",	--994
		x"1f",	--995
		x"04",	--996
		x"b0",	--997
		x"f8",	--998
		x"0b",	--999
		x"0f",	--1000
		x"0a",	--1001
		x"30",	--1002
		x"62",	--1003
		x"b0",	--1004
		x"00",	--1005
		x"31",	--1006
		x"06",	--1007
		x"0e",	--1008
		x"0f",	--1009
		x"b0",	--1010
		x"ba",	--1011
		x"0c",	--1012
		x"3d",	--1013
		x"c8",	--1014
		x"b0",	--1015
		x"44",	--1016
		x"0c",	--1017
		x"0d",	--1018
		x"0e",	--1019
		x"3f",	--1020
		x"80",	--1021
		x"b0",	--1022
		x"d0",	--1023
		x"0d",	--1024
		x"0e",	--1025
		x"1f",	--1026
		x"6e",	--1027
		x"b0",	--1028
		x"e2",	--1029
		x"0e",	--1030
		x"0f",	--1031
		x"b0",	--1032
		x"ba",	--1033
		x"0c",	--1034
		x"3d",	--1035
		x"c8",	--1036
		x"b0",	--1037
		x"44",	--1038
		x"0d",	--1039
		x"0e",	--1040
		x"1f",	--1041
		x"6c",	--1042
		x"b0",	--1043
		x"e2",	--1044
		x"0f",	--1045
		x"21",	--1046
		x"3a",	--1047
		x"3b",	--1048
		x"30",	--1049
		x"0e",	--1050
		x"1f",	--1051
		x"06",	--1052
		x"b0",	--1053
		x"f8",	--1054
		x"1d",	--1055
		x"0e",	--1056
		x"1f",	--1057
		x"04",	--1058
		x"b0",	--1059
		x"0e",	--1060
		x"b6",	--1061
		x"0e",	--1062
		x"3f",	--1063
		x"64",	--1064
		x"b0",	--1065
		x"ca",	--1066
		x"82",	--1067
		x"04",	--1068
		x"aa",	--1069
		x"30",	--1070
		x"1c",	--1071
		x"b0",	--1072
		x"00",	--1073
		x"b1",	--1074
		x"36",	--1075
		x"00",	--1076
		x"b0",	--1077
		x"00",	--1078
		x"a1",	--1079
		x"00",	--1080
		x"30",	--1081
		x"47",	--1082
		x"b0",	--1083
		x"00",	--1084
		x"21",	--1085
		x"3f",	--1086
		x"d6",	--1087
		x"0b",	--1088
		x"0a",	--1089
		x"1f",	--1090
		x"72",	--1091
		x"b0",	--1092
		x"ea",	--1093
		x"0a",	--1094
		x"0b",	--1095
		x"1f",	--1096
		x"70",	--1097
		x"b0",	--1098
		x"ea",	--1099
		x"0b",	--1100
		x"0a",	--1101
		x"3e",	--1102
		x"3f",	--1103
		x"1e",	--1104
		x"0f",	--1105
		x"0f",	--1106
		x"0e",	--1107
		x"30",	--1108
		x"6a",	--1109
		x"30",	--1110
		x"2c",	--1111
		x"b0",	--1112
		x"12",	--1113
		x"31",	--1114
		x"0c",	--1115
		x"30",	--1116
		x"2c",	--1117
		x"30",	--1118
		x"72",	--1119
		x"b0",	--1120
		x"00",	--1121
		x"21",	--1122
		x"3a",	--1123
		x"3b",	--1124
		x"30",	--1125
		x"82",	--1126
		x"70",	--1127
		x"82",	--1128
		x"72",	--1129
		x"30",	--1130
		x"82",	--1131
		x"6e",	--1132
		x"82",	--1133
		x"6c",	--1134
		x"30",	--1135
		x"0b",	--1136
		x"0a",	--1137
		x"09",	--1138
		x"08",	--1139
		x"21",	--1140
		x"0a",	--1141
		x"0b",	--1142
		x"81",	--1143
		x"00",	--1144
		x"1f",	--1145
		x"1c",	--1146
		x"b2",	--1147
		x"06",	--1148
		x"6f",	--1149
		x"92",	--1150
		x"12",	--1151
		x"0e",	--1152
		x"1f",	--1153
		x"02",	--1154
		x"b0",	--1155
		x"f8",	--1156
		x"08",	--1157
		x"3a",	--1158
		x"03",	--1159
		x"1e",	--1160
		x"09",	--1161
		x"0d",	--1162
		x"0e",	--1163
		x"1f",	--1164
		x"06",	--1165
		x"b0",	--1166
		x"0e",	--1167
		x"0f",	--1168
		x"21",	--1169
		x"38",	--1170
		x"39",	--1171
		x"3a",	--1172
		x"3b",	--1173
		x"30",	--1174
		x"82",	--1175
		x"12",	--1176
		x"49",	--1177
		x"82",	--1178
		x"12",	--1179
		x"1f",	--1180
		x"06",	--1181
		x"b0",	--1182
		x"36",	--1183
		x"0f",	--1184
		x"21",	--1185
		x"38",	--1186
		x"39",	--1187
		x"3a",	--1188
		x"3b",	--1189
		x"30",	--1190
		x"0e",	--1191
		x"1f",	--1192
		x"04",	--1193
		x"b0",	--1194
		x"f8",	--1195
		x"09",	--1196
		x"3a",	--1197
		x"05",	--1198
		x"da",	--1199
		x"0e",	--1200
		x"1f",	--1201
		x"06",	--1202
		x"b0",	--1203
		x"f8",	--1204
		x"0a",	--1205
		x"0e",	--1206
		x"1f",	--1207
		x"08",	--1208
		x"b0",	--1209
		x"f8",	--1210
		x"0b",	--1211
		x"0f",	--1212
		x"0a",	--1213
		x"30",	--1214
		x"77",	--1215
		x"b0",	--1216
		x"00",	--1217
		x"31",	--1218
		x"06",	--1219
		x"0e",	--1220
		x"0f",	--1221
		x"b0",	--1222
		x"ba",	--1223
		x"0c",	--1224
		x"3d",	--1225
		x"c8",	--1226
		x"b0",	--1227
		x"44",	--1228
		x"0d",	--1229
		x"0e",	--1230
		x"1f",	--1231
		x"6e",	--1232
		x"b0",	--1233
		x"e2",	--1234
		x"0e",	--1235
		x"0f",	--1236
		x"b0",	--1237
		x"ba",	--1238
		x"0c",	--1239
		x"3d",	--1240
		x"c8",	--1241
		x"b0",	--1242
		x"44",	--1243
		x"0d",	--1244
		x"0e",	--1245
		x"1f",	--1246
		x"6c",	--1247
		x"b0",	--1248
		x"e2",	--1249
		x"a7",	--1250
		x"0f",	--1251
		x"b0",	--1252
		x"80",	--1253
		x"0f",	--1254
		x"21",	--1255
		x"38",	--1256
		x"39",	--1257
		x"3a",	--1258
		x"3b",	--1259
		x"30",	--1260
		x"0e",	--1261
		x"3f",	--1262
		x"80",	--1263
		x"b0",	--1264
		x"ca",	--1265
		x"82",	--1266
		x"06",	--1267
		x"89",	--1268
		x"1f",	--1269
		x"82",	--1270
		x"14",	--1271
		x"01",	--1272
		x"0f",	--1273
		x"82",	--1274
		x"14",	--1275
		x"0f",	--1276
		x"30",	--1277
		x"5e",	--1278
		x"19",	--1279
		x"4e",	--1280
		x"0f",	--1281
		x"03",	--1282
		x"c2",	--1283
		x"19",	--1284
		x"30",	--1285
		x"c2",	--1286
		x"19",	--1287
		x"30",	--1288
		x"1e",	--1289
		x"16",	--1290
		x"3e",	--1291
		x"06",	--1292
		x"0f",	--1293
		x"0f",	--1294
		x"10",	--1295
		x"80",	--1296
		x"c2",	--1297
		x"19",	--1298
		x"3e",	--1299
		x"07",	--1300
		x"03",	--1301
		x"82",	--1302
		x"16",	--1303
		x"30",	--1304
		x"1e",	--1305
		x"82",	--1306
		x"16",	--1307
		x"30",	--1308
		x"f2",	--1309
		x"0e",	--1310
		x"19",	--1311
		x"f2",	--1312
		x"f2",	--1313
		x"0a",	--1314
		x"19",	--1315
		x"ee",	--1316
		x"e2",	--1317
		x"19",	--1318
		x"eb",	--1319
		x"f2",	--1320
		x"0d",	--1321
		x"19",	--1322
		x"e7",	--1323
		x"f2",	--1324
		x"09",	--1325
		x"19",	--1326
		x"e3",	--1327
		x"f2",	--1328
		x"03",	--1329
		x"19",	--1330
		x"df",	--1331
		x"f2",	--1332
		x"07",	--1333
		x"19",	--1334
		x"db",	--1335
		x"8f",	--1336
		x"00",	--1337
		x"8f",	--1338
		x"02",	--1339
		x"9f",	--1340
		x"02",	--1341
		x"04",	--1342
		x"9f",	--1343
		x"04",	--1344
		x"06",	--1345
		x"9f",	--1346
		x"06",	--1347
		x"08",	--1348
		x"9f",	--1349
		x"08",	--1350
		x"0a",	--1351
		x"9f",	--1352
		x"0a",	--1353
		x"10",	--1354
		x"9f",	--1355
		x"0c",	--1356
		x"12",	--1357
		x"8f",	--1358
		x"14",	--1359
		x"8f",	--1360
		x"16",	--1361
		x"8f",	--1362
		x"0c",	--1363
		x"8f",	--1364
		x"0e",	--1365
		x"8f",	--1366
		x"18",	--1367
		x"8f",	--1368
		x"1a",	--1369
		x"8f",	--1370
		x"1c",	--1371
		x"8f",	--1372
		x"1e",	--1373
		x"30",	--1374
		x"8f",	--1375
		x"0c",	--1376
		x"8f",	--1377
		x"0e",	--1378
		x"8f",	--1379
		x"18",	--1380
		x"8f",	--1381
		x"1a",	--1382
		x"8f",	--1383
		x"1c",	--1384
		x"8f",	--1385
		x"1e",	--1386
		x"30",	--1387
		x"8f",	--1388
		x"00",	--1389
		x"8f",	--1390
		x"02",	--1391
		x"30",	--1392
		x"8f",	--1393
		x"04",	--1394
		x"8f",	--1395
		x"06",	--1396
		x"30",	--1397
		x"8f",	--1398
		x"08",	--1399
		x"8f",	--1400
		x"0a",	--1401
		x"30",	--1402
		x"8f",	--1403
		x"0c",	--1404
		x"8f",	--1405
		x"0e",	--1406
		x"30",	--1407
		x"8f",	--1408
		x"10",	--1409
		x"8f",	--1410
		x"12",	--1411
		x"30",	--1412
		x"0b",	--1413
		x"0a",	--1414
		x"09",	--1415
		x"07",	--1416
		x"06",	--1417
		x"05",	--1418
		x"04",	--1419
		x"09",	--1420
		x"04",	--1421
		x"05",	--1422
		x"16",	--1423
		x"14",	--1424
		x"17",	--1425
		x"16",	--1426
		x"1a",	--1427
		x"0c",	--1428
		x"1b",	--1429
		x"0e",	--1430
		x"0c",	--1431
		x"0d",	--1432
		x"0e",	--1433
		x"0f",	--1434
		x"b0",	--1435
		x"34",	--1436
		x"1c",	--1437
		x"10",	--1438
		x"1d",	--1439
		x"12",	--1440
		x"0f",	--1441
		x"5b",	--1442
		x"0e",	--1443
		x"0f",	--1444
		x"b0",	--1445
		x"84",	--1446
		x"06",	--1447
		x"07",	--1448
		x"89",	--1449
		x"14",	--1450
		x"89",	--1451
		x"16",	--1452
		x"0c",	--1453
		x"0d",	--1454
		x"0e",	--1455
		x"0f",	--1456
		x"b0",	--1457
		x"34",	--1458
		x"0f",	--1459
		x"5c",	--1460
		x"89",	--1461
		x"14",	--1462
		x"89",	--1463
		x"16",	--1464
		x"0c",	--1465
		x"0d",	--1466
		x"0e",	--1467
		x"0f",	--1468
		x"b0",	--1469
		x"d0",	--1470
		x"0a",	--1471
		x"0b",	--1472
		x"1c",	--1473
		x"18",	--1474
		x"1d",	--1475
		x"1a",	--1476
		x"b0",	--1477
		x"84",	--1478
		x"06",	--1479
		x"07",	--1480
		x"89",	--1481
		x"18",	--1482
		x"89",	--1483
		x"1a",	--1484
		x"2c",	--1485
		x"1d",	--1486
		x"02",	--1487
		x"0e",	--1488
		x"0f",	--1489
		x"b0",	--1490
		x"20",	--1491
		x"04",	--1492
		x"05",	--1493
		x"1c",	--1494
		x"04",	--1495
		x"1d",	--1496
		x"06",	--1497
		x"0e",	--1498
		x"0f",	--1499
		x"b0",	--1500
		x"20",	--1501
		x"0c",	--1502
		x"0d",	--1503
		x"b0",	--1504
		x"84",	--1505
		x"06",	--1506
		x"07",	--1507
		x"1c",	--1508
		x"1c",	--1509
		x"1d",	--1510
		x"1e",	--1511
		x"0e",	--1512
		x"0f",	--1513
		x"b0",	--1514
		x"d0",	--1515
		x"1c",	--1516
		x"08",	--1517
		x"1d",	--1518
		x"0a",	--1519
		x"b0",	--1520
		x"20",	--1521
		x"0c",	--1522
		x"0d",	--1523
		x"b0",	--1524
		x"84",	--1525
		x"34",	--1526
		x"35",	--1527
		x"36",	--1528
		x"37",	--1529
		x"39",	--1530
		x"3a",	--1531
		x"3b",	--1532
		x"30",	--1533
		x"0e",	--1534
		x"0f",	--1535
		x"b0",	--1536
		x"d0",	--1537
		x"06",	--1538
		x"07",	--1539
		x"89",	--1540
		x"14",	--1541
		x"89",	--1542
		x"16",	--1543
		x"0c",	--1544
		x"0d",	--1545
		x"0e",	--1546
		x"0f",	--1547
		x"b0",	--1548
		x"94",	--1549
		x"0f",	--1550
		x"01",	--1551
		x"a4",	--1552
		x"0a",	--1553
		x"0b",	--1554
		x"a5",	--1555
		x"0b",	--1556
		x"0a",	--1557
		x"21",	--1558
		x"0a",	--1559
		x"0b",	--1560
		x"30",	--1561
		x"38",	--1562
		x"b0",	--1563
		x"00",	--1564
		x"21",	--1565
		x"3a",	--1566
		x"03",	--1567
		x"1b",	--1568
		x"0e",	--1569
		x"1f",	--1570
		x"02",	--1571
		x"b0",	--1572
		x"f8",	--1573
		x"0a",	--1574
		x"0e",	--1575
		x"1f",	--1576
		x"04",	--1577
		x"b0",	--1578
		x"f8",	--1579
		x"0b",	--1580
		x"0f",	--1581
		x"0a",	--1582
		x"30",	--1583
		x"80",	--1584
		x"b0",	--1585
		x"00",	--1586
		x"31",	--1587
		x"06",	--1588
		x"8a",	--1589
		x"00",	--1590
		x"0f",	--1591
		x"21",	--1592
		x"3a",	--1593
		x"3b",	--1594
		x"30",	--1595
		x"30",	--1596
		x"40",	--1597
		x"b0",	--1598
		x"00",	--1599
		x"b1",	--1600
		x"5a",	--1601
		x"00",	--1602
		x"b0",	--1603
		x"00",	--1604
		x"a1",	--1605
		x"00",	--1606
		x"30",	--1607
		x"6b",	--1608
		x"b0",	--1609
		x"00",	--1610
		x"21",	--1611
		x"3f",	--1612
		x"ea",	--1613
		x"0b",	--1614
		x"21",	--1615
		x"0b",	--1616
		x"1f",	--1617
		x"17",	--1618
		x"16",	--1619
		x"30",	--1620
		x"9b",	--1621
		x"b0",	--1622
		x"00",	--1623
		x"21",	--1624
		x"0e",	--1625
		x"1f",	--1626
		x"02",	--1627
		x"b0",	--1628
		x"f8",	--1629
		x"2f",	--1630
		x"0f",	--1631
		x"30",	--1632
		x"80",	--1633
		x"b0",	--1634
		x"00",	--1635
		x"31",	--1636
		x"06",	--1637
		x"0f",	--1638
		x"21",	--1639
		x"3b",	--1640
		x"30",	--1641
		x"30",	--1642
		x"40",	--1643
		x"b0",	--1644
		x"00",	--1645
		x"b1",	--1646
		x"5a",	--1647
		x"00",	--1648
		x"b0",	--1649
		x"00",	--1650
		x"a1",	--1651
		x"00",	--1652
		x"30",	--1653
		x"8c",	--1654
		x"b0",	--1655
		x"00",	--1656
		x"21",	--1657
		x"3f",	--1658
		x"eb",	--1659
		x"0b",	--1660
		x"0a",	--1661
		x"8e",	--1662
		x"00",	--1663
		x"6d",	--1664
		x"4d",	--1665
		x"5e",	--1666
		x"1f",	--1667
		x"0a",	--1668
		x"0c",	--1669
		x"0f",	--1670
		x"7b",	--1671
		x"0a",	--1672
		x"2b",	--1673
		x"0c",	--1674
		x"0c",	--1675
		x"0c",	--1676
		x"0c",	--1677
		x"8d",	--1678
		x"0c",	--1679
		x"3c",	--1680
		x"d0",	--1681
		x"1a",	--1682
		x"7d",	--1683
		x"4d",	--1684
		x"17",	--1685
		x"7d",	--1686
		x"78",	--1687
		x"1a",	--1688
		x"4b",	--1689
		x"7b",	--1690
		x"d0",	--1691
		x"0a",	--1692
		x"e9",	--1693
		x"7b",	--1694
		x"0a",	--1695
		x"34",	--1696
		x"0c",	--1697
		x"0b",	--1698
		x"0b",	--1699
		x"0b",	--1700
		x"0c",	--1701
		x"8d",	--1702
		x"0c",	--1703
		x"3c",	--1704
		x"d0",	--1705
		x"7d",	--1706
		x"4d",	--1707
		x"e9",	--1708
		x"9e",	--1709
		x"00",	--1710
		x"0f",	--1711
		x"3a",	--1712
		x"3b",	--1713
		x"30",	--1714
		x"1a",	--1715
		x"de",	--1716
		x"4b",	--1717
		x"7b",	--1718
		x"9f",	--1719
		x"7b",	--1720
		x"06",	--1721
		x"0a",	--1722
		x"0c",	--1723
		x"0c",	--1724
		x"0c",	--1725
		x"0c",	--1726
		x"8d",	--1727
		x"0c",	--1728
		x"3c",	--1729
		x"a9",	--1730
		x"1a",	--1731
		x"ce",	--1732
		x"4b",	--1733
		x"7b",	--1734
		x"bf",	--1735
		x"7b",	--1736
		x"06",	--1737
		x"0a",	--1738
		x"0c",	--1739
		x"0c",	--1740
		x"0c",	--1741
		x"0c",	--1742
		x"8d",	--1743
		x"0c",	--1744
		x"3c",	--1745
		x"c9",	--1746
		x"1a",	--1747
		x"be",	--1748
		x"8d",	--1749
		x"0d",	--1750
		x"30",	--1751
		x"a2",	--1752
		x"b0",	--1753
		x"00",	--1754
		x"21",	--1755
		x"0c",	--1756
		x"0f",	--1757
		x"3a",	--1758
		x"3b",	--1759
		x"30",	--1760
		x"0c",	--1761
		x"ca",	--1762
		x"0b",	--1763
		x"0a",	--1764
		x"8e",	--1765
		x"00",	--1766
		x"6b",	--1767
		x"4b",	--1768
		x"37",	--1769
		x"1f",	--1770
		x"1a",	--1771
		x"0c",	--1772
		x"12",	--1773
		x"4d",	--1774
		x"7d",	--1775
		x"d0",	--1776
		x"7d",	--1777
		x"0a",	--1778
		x"22",	--1779
		x"0c",	--1780
		x"0d",	--1781
		x"0d",	--1782
		x"0d",	--1783
		x"0c",	--1784
		x"8b",	--1785
		x"0c",	--1786
		x"3c",	--1787
		x"d0",	--1788
		x"7b",	--1789
		x"4b",	--1790
		x"07",	--1791
		x"7b",	--1792
		x"2d",	--1793
		x"eb",	--1794
		x"3a",	--1795
		x"7b",	--1796
		x"4b",	--1797
		x"f9",	--1798
		x"02",	--1799
		x"32",	--1800
		x"03",	--1801
		x"82",	--1802
		x"32",	--1803
		x"82",	--1804
		x"38",	--1805
		x"1f",	--1806
		x"3a",	--1807
		x"32",	--1808
		x"9e",	--1809
		x"00",	--1810
		x"3a",	--1811
		x"3b",	--1812
		x"30",	--1813
		x"8b",	--1814
		x"0b",	--1815
		x"30",	--1816
		x"a2",	--1817
		x"b0",	--1818
		x"00",	--1819
		x"21",	--1820
		x"0f",	--1821
		x"3a",	--1822
		x"3b",	--1823
		x"30",	--1824
		x"0f",	--1825
		x"ee",	--1826
		x"0b",	--1827
		x"0a",	--1828
		x"0b",	--1829
		x"0a",	--1830
		x"8f",	--1831
		x"00",	--1832
		x"8f",	--1833
		x"02",	--1834
		x"8f",	--1835
		x"04",	--1836
		x"0c",	--1837
		x"0d",	--1838
		x"3e",	--1839
		x"00",	--1840
		x"3f",	--1841
		x"6e",	--1842
		x"b0",	--1843
		x"20",	--1844
		x"8b",	--1845
		x"02",	--1846
		x"02",	--1847
		x"32",	--1848
		x"03",	--1849
		x"82",	--1850
		x"32",	--1851
		x"b2",	--1852
		x"18",	--1853
		x"38",	--1854
		x"9b",	--1855
		x"3a",	--1856
		x"06",	--1857
		x"32",	--1858
		x"0f",	--1859
		x"3a",	--1860
		x"3b",	--1861
		x"30",	--1862
		x"0b",	--1863
		x"09",	--1864
		x"08",	--1865
		x"8f",	--1866
		x"06",	--1867
		x"bf",	--1868
		x"00",	--1869
		x"08",	--1870
		x"2b",	--1871
		x"1e",	--1872
		x"02",	--1873
		x"0f",	--1874
		x"b0",	--1875
		x"ba",	--1876
		x"0c",	--1877
		x"3d",	--1878
		x"00",	--1879
		x"b0",	--1880
		x"20",	--1881
		x"08",	--1882
		x"09",	--1883
		x"1e",	--1884
		x"06",	--1885
		x"0f",	--1886
		x"b0",	--1887
		x"ba",	--1888
		x"0c",	--1889
		x"0d",	--1890
		x"0e",	--1891
		x"0f",	--1892
		x"b0",	--1893
		x"d0",	--1894
		x"b0",	--1895
		x"b0",	--1896
		x"8b",	--1897
		x"04",	--1898
		x"9b",	--1899
		x"00",	--1900
		x"38",	--1901
		x"39",	--1902
		x"3b",	--1903
		x"30",	--1904
		x"0b",	--1905
		x"0a",	--1906
		x"09",	--1907
		x"0a",	--1908
		x"0b",	--1909
		x"8f",	--1910
		x"06",	--1911
		x"8f",	--1912
		x"08",	--1913
		x"29",	--1914
		x"1e",	--1915
		x"02",	--1916
		x"0f",	--1917
		x"b0",	--1918
		x"ba",	--1919
		x"0c",	--1920
		x"0d",	--1921
		x"0e",	--1922
		x"0f",	--1923
		x"b0",	--1924
		x"20",	--1925
		x"0a",	--1926
		x"0b",	--1927
		x"1e",	--1928
		x"06",	--1929
		x"0f",	--1930
		x"b0",	--1931
		x"ba",	--1932
		x"0c",	--1933
		x"0d",	--1934
		x"0e",	--1935
		x"0f",	--1936
		x"b0",	--1937
		x"d0",	--1938
		x"b0",	--1939
		x"b0",	--1940
		x"89",	--1941
		x"04",	--1942
		x"39",	--1943
		x"3a",	--1944
		x"3b",	--1945
		x"30",	--1946
		x"2f",	--1947
		x"8f",	--1948
		x"04",	--1949
		x"30",	--1950
		x"0b",	--1951
		x"0a",	--1952
		x"92",	--1953
		x"18",	--1954
		x"14",	--1955
		x"3b",	--1956
		x"78",	--1957
		x"0a",	--1958
		x"2b",	--1959
		x"5f",	--1960
		x"fc",	--1961
		x"8f",	--1962
		x"0f",	--1963
		x"30",	--1964
		x"b7",	--1965
		x"b0",	--1966
		x"00",	--1967
		x"31",	--1968
		x"06",	--1969
		x"1a",	--1970
		x"3b",	--1971
		x"06",	--1972
		x"1a",	--1973
		x"18",	--1974
		x"ef",	--1975
		x"0f",	--1976
		x"3a",	--1977
		x"3b",	--1978
		x"30",	--1979
		x"1e",	--1980
		x"18",	--1981
		x"3e",	--1982
		x"20",	--1983
		x"12",	--1984
		x"0f",	--1985
		x"0f",	--1986
		x"0f",	--1987
		x"0f",	--1988
		x"3f",	--1989
		x"74",	--1990
		x"ff",	--1991
		x"68",	--1992
		x"00",	--1993
		x"bf",	--1994
		x"3e",	--1995
		x"02",	--1996
		x"bf",	--1997
		x"08",	--1998
		x"04",	--1999
		x"1e",	--2000
		x"82",	--2001
		x"18",	--2002
		x"30",	--2003
		x"0b",	--2004
		x"1b",	--2005
		x"18",	--2006
		x"3b",	--2007
		x"20",	--2008
		x"12",	--2009
		x"0c",	--2010
		x"0c",	--2011
		x"0c",	--2012
		x"0c",	--2013
		x"3c",	--2014
		x"74",	--2015
		x"cc",	--2016
		x"00",	--2017
		x"8c",	--2018
		x"02",	--2019
		x"8c",	--2020
		x"04",	--2021
		x"1b",	--2022
		x"82",	--2023
		x"18",	--2024
		x"0f",	--2025
		x"3b",	--2026
		x"30",	--2027
		x"3f",	--2028
		x"fc",	--2029
		x"0b",	--2030
		x"31",	--2031
		x"f0",	--2032
		x"1b",	--2033
		x"18",	--2034
		x"1b",	--2035
		x"0f",	--2036
		x"5f",	--2037
		x"74",	--2038
		x"16",	--2039
		x"3d",	--2040
		x"7a",	--2041
		x"0c",	--2042
		x"05",	--2043
		x"3d",	--2044
		x"06",	--2045
		x"cd",	--2046
		x"fa",	--2047
		x"0e",	--2048
		x"1c",	--2049
		x"0c",	--2050
		x"f8",	--2051
		x"30",	--2052
		x"bf",	--2053
		x"b0",	--2054
		x"00",	--2055
		x"21",	--2056
		x"3f",	--2057
		x"31",	--2058
		x"10",	--2059
		x"3b",	--2060
		x"30",	--2061
		x"0c",	--2062
		x"81",	--2063
		x"00",	--2064
		x"6d",	--2065
		x"4d",	--2066
		x"24",	--2067
		x"1e",	--2068
		x"1f",	--2069
		x"06",	--2070
		x"6d",	--2071
		x"4d",	--2072
		x"11",	--2073
		x"1e",	--2074
		x"3f",	--2075
		x"0e",	--2076
		x"7d",	--2077
		x"20",	--2078
		x"f7",	--2079
		x"ce",	--2080
		x"ff",	--2081
		x"0d",	--2082
		x"0d",	--2083
		x"0d",	--2084
		x"8d",	--2085
		x"00",	--2086
		x"1f",	--2087
		x"6d",	--2088
		x"4d",	--2089
		x"ef",	--2090
		x"0e",	--2091
		x"0e",	--2092
		x"0c",	--2093
		x"0c",	--2094
		x"3c",	--2095
		x"74",	--2096
		x"0e",	--2097
		x"9c",	--2098
		x"02",	--2099
		x"31",	--2100
		x"10",	--2101
		x"3b",	--2102
		x"30",	--2103
		x"1f",	--2104
		x"f1",	--2105
		x"8f",	--2106
		x"00",	--2107
		x"0f",	--2108
		x"30",	--2109
		x"0e",	--2110
		x"2e",	--2111
		x"2f",	--2112
		x"30",	--2113
		x"0b",	--2114
		x"0a",	--2115
		x"0e",	--2116
		x"2e",	--2117
		x"2c",	--2118
		x"0d",	--2119
		x"0e",	--2120
		x"0f",	--2121
		x"0e",	--2122
		x"0f",	--2123
		x"0a",	--2124
		x"0b",	--2125
		x"0a",	--2126
		x"0b",	--2127
		x"0a",	--2128
		x"0b",	--2129
		x"3c",	--2130
		x"3a",	--2131
		x"0d",	--2132
		x"0e",	--2133
		x"0f",	--2134
		x"b0",	--2135
		x"e0",	--2136
		x"0f",	--2137
		x"3a",	--2138
		x"3b",	--2139
		x"30",	--2140
		x"b2",	--2141
		x"d2",	--2142
		x"60",	--2143
		x"b2",	--2144
		x"b8",	--2145
		x"72",	--2146
		x"0f",	--2147
		x"30",	--2148
		x"0b",	--2149
		x"0b",	--2150
		x"1f",	--2151
		x"1a",	--2152
		x"3f",	--2153
		x"20",	--2154
		x"19",	--2155
		x"0c",	--2156
		x"0c",	--2157
		x"0d",	--2158
		x"0d",	--2159
		x"0d",	--2160
		x"0d",	--2161
		x"0d",	--2162
		x"3d",	--2163
		x"34",	--2164
		x"8d",	--2165
		x"00",	--2166
		x"8d",	--2167
		x"02",	--2168
		x"8d",	--2169
		x"08",	--2170
		x"8d",	--2171
		x"0a",	--2172
		x"8d",	--2173
		x"0c",	--2174
		x"0e",	--2175
		x"1e",	--2176
		x"82",	--2177
		x"1a",	--2178
		x"3b",	--2179
		x"30",	--2180
		x"3f",	--2181
		x"fc",	--2182
		x"0f",	--2183
		x"0c",	--2184
		x"0c",	--2185
		x"0c",	--2186
		x"0c",	--2187
		x"0c",	--2188
		x"3c",	--2189
		x"34",	--2190
		x"8c",	--2191
		x"02",	--2192
		x"8c",	--2193
		x"04",	--2194
		x"8c",	--2195
		x"06",	--2196
		x"8c",	--2197
		x"08",	--2198
		x"9c",	--2199
		x"00",	--2200
		x"0f",	--2201
		x"30",	--2202
		x"0f",	--2203
		x"0e",	--2204
		x"0e",	--2205
		x"0e",	--2206
		x"0e",	--2207
		x"0e",	--2208
		x"8e",	--2209
		x"34",	--2210
		x"0f",	--2211
		x"30",	--2212
		x"0f",	--2213
		x"0e",	--2214
		x"0d",	--2215
		x"0c",	--2216
		x"0b",	--2217
		x"0a",	--2218
		x"09",	--2219
		x"08",	--2220
		x"07",	--2221
		x"92",	--2222
		x"1a",	--2223
		x"33",	--2224
		x"3a",	--2225
		x"34",	--2226
		x"0b",	--2227
		x"2b",	--2228
		x"08",	--2229
		x"38",	--2230
		x"07",	--2231
		x"37",	--2232
		x"06",	--2233
		x"09",	--2234
		x"0f",	--2235
		x"1f",	--2236
		x"8b",	--2237
		x"00",	--2238
		x"19",	--2239
		x"3a",	--2240
		x"0e",	--2241
		x"3b",	--2242
		x"0e",	--2243
		x"38",	--2244
		x"0e",	--2245
		x"37",	--2246
		x"0e",	--2247
		x"19",	--2248
		x"1a",	--2249
		x"19",	--2250
		x"8a",	--2251
		x"00",	--2252
		x"f1",	--2253
		x"2f",	--2254
		x"1f",	--2255
		x"02",	--2256
		x"ea",	--2257
		x"8b",	--2258
		x"00",	--2259
		x"1f",	--2260
		x"0a",	--2261
		x"9b",	--2262
		x"08",	--2263
		x"88",	--2264
		x"00",	--2265
		x"e4",	--2266
		x"2f",	--2267
		x"1f",	--2268
		x"87",	--2269
		x"00",	--2270
		x"2f",	--2271
		x"de",	--2272
		x"8a",	--2273
		x"00",	--2274
		x"db",	--2275
		x"b2",	--2276
		x"fe",	--2277
		x"60",	--2278
		x"37",	--2279
		x"38",	--2280
		x"39",	--2281
		x"3a",	--2282
		x"3b",	--2283
		x"3c",	--2284
		x"3d",	--2285
		x"3e",	--2286
		x"3f",	--2287
		x"00",	--2288
		x"8f",	--2289
		x"00",	--2290
		x"0f",	--2291
		x"30",	--2292
		x"2f",	--2293
		x"2e",	--2294
		x"1f",	--2295
		x"02",	--2296
		x"30",	--2297
		x"8f",	--2298
		x"00",	--2299
		x"30",	--2300
		x"8f",	--2301
		x"00",	--2302
		x"3f",	--2303
		x"f4",	--2304
		x"b0",	--2305
		x"ca",	--2306
		x"82",	--2307
		x"0e",	--2308
		x"0f",	--2309
		x"30",	--2310
		x"0c",	--2311
		x"2f",	--2312
		x"8f",	--2313
		x"00",	--2314
		x"1d",	--2315
		x"0e",	--2316
		x"1f",	--2317
		x"0e",	--2318
		x"b0",	--2319
		x"0e",	--2320
		x"30",	--2321
		x"5e",	--2322
		x"81",	--2323
		x"3e",	--2324
		x"fc",	--2325
		x"c2",	--2326
		x"84",	--2327
		x"0f",	--2328
		x"30",	--2329
		x"3f",	--2330
		x"0f",	--2331
		x"5f",	--2332
		x"7e",	--2333
		x"8f",	--2334
		x"b0",	--2335
		x"24",	--2336
		x"30",	--2337
		x"0b",	--2338
		x"0b",	--2339
		x"0e",	--2340
		x"0e",	--2341
		x"0e",	--2342
		x"0e",	--2343
		x"0e",	--2344
		x"0f",	--2345
		x"b0",	--2346
		x"34",	--2347
		x"0f",	--2348
		x"b0",	--2349
		x"34",	--2350
		x"3b",	--2351
		x"30",	--2352
		x"0b",	--2353
		x"0a",	--2354
		x"0a",	--2355
		x"3b",	--2356
		x"07",	--2357
		x"0e",	--2358
		x"4d",	--2359
		x"7d",	--2360
		x"0f",	--2361
		x"03",	--2362
		x"0e",	--2363
		x"7d",	--2364
		x"fd",	--2365
		x"1e",	--2366
		x"0a",	--2367
		x"3f",	--2368
		x"31",	--2369
		x"b0",	--2370
		x"24",	--2371
		x"3b",	--2372
		x"3b",	--2373
		x"ef",	--2374
		x"3a",	--2375
		x"3b",	--2376
		x"30",	--2377
		x"3f",	--2378
		x"30",	--2379
		x"f5",	--2380
		x"0b",	--2381
		x"0b",	--2382
		x"0e",	--2383
		x"8e",	--2384
		x"8e",	--2385
		x"0f",	--2386
		x"b0",	--2387
		x"44",	--2388
		x"0f",	--2389
		x"b0",	--2390
		x"44",	--2391
		x"3b",	--2392
		x"30",	--2393
		x"0b",	--2394
		x"0a",	--2395
		x"0a",	--2396
		x"0b",	--2397
		x"0d",	--2398
		x"8d",	--2399
		x"8d",	--2400
		x"0f",	--2401
		x"b0",	--2402
		x"44",	--2403
		x"0f",	--2404
		x"b0",	--2405
		x"44",	--2406
		x"0c",	--2407
		x"0d",	--2408
		x"8d",	--2409
		x"8c",	--2410
		x"4d",	--2411
		x"0d",	--2412
		x"0f",	--2413
		x"b0",	--2414
		x"44",	--2415
		x"0f",	--2416
		x"b0",	--2417
		x"44",	--2418
		x"3a",	--2419
		x"3b",	--2420
		x"30",	--2421
		x"0b",	--2422
		x"0a",	--2423
		x"09",	--2424
		x"0a",	--2425
		x"0e",	--2426
		x"19",	--2427
		x"09",	--2428
		x"39",	--2429
		x"0b",	--2430
		x"0d",	--2431
		x"0d",	--2432
		x"6f",	--2433
		x"8f",	--2434
		x"b0",	--2435
		x"44",	--2436
		x"0b",	--2437
		x"0e",	--2438
		x"1b",	--2439
		x"3b",	--2440
		x"07",	--2441
		x"05",	--2442
		x"3f",	--2443
		x"20",	--2444
		x"b0",	--2445
		x"24",	--2446
		x"ef",	--2447
		x"3f",	--2448
		x"3a",	--2449
		x"b0",	--2450
		x"24",	--2451
		x"ea",	--2452
		x"39",	--2453
		x"3a",	--2454
		x"3b",	--2455
		x"30",	--2456
		x"0b",	--2457
		x"0a",	--2458
		x"09",	--2459
		x"0a",	--2460
		x"0e",	--2461
		x"17",	--2462
		x"09",	--2463
		x"39",	--2464
		x"0b",	--2465
		x"6f",	--2466
		x"8f",	--2467
		x"b0",	--2468
		x"34",	--2469
		x"0b",	--2470
		x"0e",	--2471
		x"1b",	--2472
		x"3b",	--2473
		x"07",	--2474
		x"f6",	--2475
		x"3f",	--2476
		x"20",	--2477
		x"b0",	--2478
		x"24",	--2479
		x"6f",	--2480
		x"8f",	--2481
		x"b0",	--2482
		x"34",	--2483
		x"0b",	--2484
		x"f2",	--2485
		x"39",	--2486
		x"3a",	--2487
		x"3b",	--2488
		x"30",	--2489
		x"0b",	--2490
		x"0a",	--2491
		x"09",	--2492
		x"31",	--2493
		x"ec",	--2494
		x"0b",	--2495
		x"0f",	--2496
		x"34",	--2497
		x"3b",	--2498
		x"0a",	--2499
		x"38",	--2500
		x"09",	--2501
		x"0a",	--2502
		x"0a",	--2503
		x"3e",	--2504
		x"0a",	--2505
		x"0f",	--2506
		x"b0",	--2507
		x"d8",	--2508
		x"7f",	--2509
		x"30",	--2510
		x"ca",	--2511
		x"00",	--2512
		x"19",	--2513
		x"3e",	--2514
		x"0a",	--2515
		x"0f",	--2516
		x"b0",	--2517
		x"a6",	--2518
		x"0b",	--2519
		x"3f",	--2520
		x"0a",	--2521
		x"eb",	--2522
		x"0a",	--2523
		x"1a",	--2524
		x"09",	--2525
		x"3e",	--2526
		x"0a",	--2527
		x"0f",	--2528
		x"b0",	--2529
		x"d8",	--2530
		x"7f",	--2531
		x"30",	--2532
		x"c9",	--2533
		x"00",	--2534
		x"3a",	--2535
		x"0f",	--2536
		x"0f",	--2537
		x"6f",	--2538
		x"8f",	--2539
		x"b0",	--2540
		x"24",	--2541
		x"0a",	--2542
		x"f7",	--2543
		x"31",	--2544
		x"14",	--2545
		x"39",	--2546
		x"3a",	--2547
		x"3b",	--2548
		x"30",	--2549
		x"3f",	--2550
		x"2d",	--2551
		x"b0",	--2552
		x"24",	--2553
		x"3b",	--2554
		x"1b",	--2555
		x"c5",	--2556
		x"1a",	--2557
		x"09",	--2558
		x"dd",	--2559
		x"0b",	--2560
		x"0a",	--2561
		x"09",	--2562
		x"0b",	--2563
		x"3b",	--2564
		x"39",	--2565
		x"6f",	--2566
		x"4f",	--2567
		x"0b",	--2568
		x"1a",	--2569
		x"8f",	--2570
		x"b0",	--2571
		x"24",	--2572
		x"0a",	--2573
		x"09",	--2574
		x"19",	--2575
		x"5f",	--2576
		x"01",	--2577
		x"4f",	--2578
		x"10",	--2579
		x"7f",	--2580
		x"25",	--2581
		x"f3",	--2582
		x"0a",	--2583
		x"1a",	--2584
		x"5f",	--2585
		x"01",	--2586
		x"7f",	--2587
		x"db",	--2588
		x"7f",	--2589
		x"54",	--2590
		x"ee",	--2591
		x"4f",	--2592
		x"0f",	--2593
		x"10",	--2594
		x"d6",	--2595
		x"39",	--2596
		x"3a",	--2597
		x"3b",	--2598
		x"30",	--2599
		x"09",	--2600
		x"29",	--2601
		x"1e",	--2602
		x"02",	--2603
		x"2f",	--2604
		x"b0",	--2605
		x"ec",	--2606
		x"0b",	--2607
		x"dd",	--2608
		x"09",	--2609
		x"29",	--2610
		x"2f",	--2611
		x"b0",	--2612
		x"9a",	--2613
		x"0b",	--2614
		x"d6",	--2615
		x"0f",	--2616
		x"2b",	--2617
		x"29",	--2618
		x"6f",	--2619
		x"4f",	--2620
		x"d0",	--2621
		x"19",	--2622
		x"8f",	--2623
		x"b0",	--2624
		x"24",	--2625
		x"7f",	--2626
		x"4f",	--2627
		x"fa",	--2628
		x"c8",	--2629
		x"09",	--2630
		x"29",	--2631
		x"1e",	--2632
		x"02",	--2633
		x"2f",	--2634
		x"b0",	--2635
		x"32",	--2636
		x"0b",	--2637
		x"bf",	--2638
		x"09",	--2639
		x"29",	--2640
		x"2e",	--2641
		x"0f",	--2642
		x"8f",	--2643
		x"8f",	--2644
		x"8f",	--2645
		x"8f",	--2646
		x"b0",	--2647
		x"b4",	--2648
		x"0b",	--2649
		x"b3",	--2650
		x"09",	--2651
		x"29",	--2652
		x"2f",	--2653
		x"b0",	--2654
		x"74",	--2655
		x"0b",	--2656
		x"ac",	--2657
		x"09",	--2658
		x"29",	--2659
		x"2f",	--2660
		x"b0",	--2661
		x"24",	--2662
		x"0b",	--2663
		x"a5",	--2664
		x"09",	--2665
		x"29",	--2666
		x"2f",	--2667
		x"b0",	--2668
		x"44",	--2669
		x"0b",	--2670
		x"9e",	--2671
		x"09",	--2672
		x"29",	--2673
		x"2f",	--2674
		x"b0",	--2675
		x"62",	--2676
		x"0b",	--2677
		x"97",	--2678
		x"3f",	--2679
		x"25",	--2680
		x"b0",	--2681
		x"24",	--2682
		x"92",	--2683
		x"0f",	--2684
		x"0e",	--2685
		x"1f",	--2686
		x"1c",	--2687
		x"df",	--2688
		x"85",	--2689
		x"f4",	--2690
		x"1f",	--2691
		x"1c",	--2692
		x"3f",	--2693
		x"3f",	--2694
		x"13",	--2695
		x"92",	--2696
		x"1c",	--2697
		x"1e",	--2698
		x"1c",	--2699
		x"1f",	--2700
		x"1e",	--2701
		x"0e",	--2702
		x"02",	--2703
		x"92",	--2704
		x"1e",	--2705
		x"f2",	--2706
		x"10",	--2707
		x"81",	--2708
		x"3e",	--2709
		x"3f",	--2710
		x"b1",	--2711
		x"f0",	--2712
		x"00",	--2713
		x"00",	--2714
		x"82",	--2715
		x"1c",	--2716
		x"ec",	--2717
		x"0c",	--2718
		x"0d",	--2719
		x"3e",	--2720
		x"00",	--2721
		x"3f",	--2722
		x"6e",	--2723
		x"b0",	--2724
		x"e0",	--2725
		x"3e",	--2726
		x"82",	--2727
		x"82",	--2728
		x"f2",	--2729
		x"11",	--2730
		x"80",	--2731
		x"30",	--2732
		x"1e",	--2733
		x"1c",	--2734
		x"1f",	--2735
		x"1e",	--2736
		x"0e",	--2737
		x"05",	--2738
		x"1f",	--2739
		x"1c",	--2740
		x"1f",	--2741
		x"1e",	--2742
		x"30",	--2743
		x"1d",	--2744
		x"1c",	--2745
		x"1e",	--2746
		x"1e",	--2747
		x"3f",	--2748
		x"40",	--2749
		x"0f",	--2750
		x"0f",	--2751
		x"30",	--2752
		x"1f",	--2753
		x"1e",	--2754
		x"5f",	--2755
		x"f4",	--2756
		x"1d",	--2757
		x"1e",	--2758
		x"1e",	--2759
		x"1c",	--2760
		x"0d",	--2761
		x"0b",	--2762
		x"1e",	--2763
		x"1e",	--2764
		x"3e",	--2765
		x"3f",	--2766
		x"03",	--2767
		x"82",	--2768
		x"1e",	--2769
		x"30",	--2770
		x"92",	--2771
		x"1e",	--2772
		x"30",	--2773
		x"4f",	--2774
		x"30",	--2775
		x"0b",	--2776
		x"0a",	--2777
		x"0a",	--2778
		x"0b",	--2779
		x"0c",	--2780
		x"3d",	--2781
		x"00",	--2782
		x"b0",	--2783
		x"e4",	--2784
		x"0f",	--2785
		x"07",	--2786
		x"0e",	--2787
		x"0f",	--2788
		x"b0",	--2789
		x"2a",	--2790
		x"3a",	--2791
		x"3b",	--2792
		x"30",	--2793
		x"0c",	--2794
		x"3d",	--2795
		x"00",	--2796
		x"0e",	--2797
		x"0f",	--2798
		x"b0",	--2799
		x"d0",	--2800
		x"b0",	--2801
		x"2a",	--2802
		x"0e",	--2803
		x"3f",	--2804
		x"00",	--2805
		x"3a",	--2806
		x"3b",	--2807
		x"30",	--2808
		x"0b",	--2809
		x"0a",	--2810
		x"09",	--2811
		x"08",	--2812
		x"07",	--2813
		x"06",	--2814
		x"05",	--2815
		x"04",	--2816
		x"31",	--2817
		x"fa",	--2818
		x"08",	--2819
		x"6b",	--2820
		x"6b",	--2821
		x"67",	--2822
		x"6c",	--2823
		x"6c",	--2824
		x"e9",	--2825
		x"6b",	--2826
		x"02",	--2827
		x"30",	--2828
		x"72",	--2829
		x"6c",	--2830
		x"e3",	--2831
		x"6c",	--2832
		x"bb",	--2833
		x"6b",	--2834
		x"df",	--2835
		x"91",	--2836
		x"02",	--2837
		x"00",	--2838
		x"1b",	--2839
		x"02",	--2840
		x"14",	--2841
		x"04",	--2842
		x"15",	--2843
		x"06",	--2844
		x"16",	--2845
		x"04",	--2846
		x"17",	--2847
		x"06",	--2848
		x"2c",	--2849
		x"0c",	--2850
		x"09",	--2851
		x"0c",	--2852
		x"bf",	--2853
		x"39",	--2854
		x"20",	--2855
		x"50",	--2856
		x"1c",	--2857
		x"d7",	--2858
		x"81",	--2859
		x"02",	--2860
		x"81",	--2861
		x"04",	--2862
		x"4c",	--2863
		x"7c",	--2864
		x"1f",	--2865
		x"0b",	--2866
		x"0a",	--2867
		x"0b",	--2868
		x"12",	--2869
		x"0b",	--2870
		x"0a",	--2871
		x"7c",	--2872
		x"fb",	--2873
		x"81",	--2874
		x"02",	--2875
		x"81",	--2876
		x"04",	--2877
		x"1c",	--2878
		x"0d",	--2879
		x"79",	--2880
		x"1f",	--2881
		x"04",	--2882
		x"0c",	--2883
		x"0d",	--2884
		x"79",	--2885
		x"fc",	--2886
		x"3c",	--2887
		x"3d",	--2888
		x"0c",	--2889
		x"0d",	--2890
		x"1a",	--2891
		x"0b",	--2892
		x"0c",	--2893
		x"02",	--2894
		x"0d",	--2895
		x"e5",	--2896
		x"16",	--2897
		x"02",	--2898
		x"17",	--2899
		x"04",	--2900
		x"06",	--2901
		x"07",	--2902
		x"5f",	--2903
		x"01",	--2904
		x"5f",	--2905
		x"01",	--2906
		x"28",	--2907
		x"c8",	--2908
		x"01",	--2909
		x"a8",	--2910
		x"02",	--2911
		x"0e",	--2912
		x"0f",	--2913
		x"0e",	--2914
		x"0f",	--2915
		x"88",	--2916
		x"04",	--2917
		x"88",	--2918
		x"06",	--2919
		x"f8",	--2920
		x"03",	--2921
		x"00",	--2922
		x"0f",	--2923
		x"4d",	--2924
		x"0f",	--2925
		x"31",	--2926
		x"06",	--2927
		x"34",	--2928
		x"35",	--2929
		x"36",	--2930
		x"37",	--2931
		x"38",	--2932
		x"39",	--2933
		x"3a",	--2934
		x"3b",	--2935
		x"30",	--2936
		x"2b",	--2937
		x"67",	--2938
		x"81",	--2939
		x"00",	--2940
		x"04",	--2941
		x"05",	--2942
		x"5f",	--2943
		x"01",	--2944
		x"5f",	--2945
		x"01",	--2946
		x"d8",	--2947
		x"4f",	--2948
		x"68",	--2949
		x"0e",	--2950
		x"0f",	--2951
		x"0e",	--2952
		x"0f",	--2953
		x"0f",	--2954
		x"69",	--2955
		x"c8",	--2956
		x"01",	--2957
		x"a8",	--2958
		x"02",	--2959
		x"88",	--2960
		x"04",	--2961
		x"88",	--2962
		x"06",	--2963
		x"0c",	--2964
		x"0d",	--2965
		x"3c",	--2966
		x"3d",	--2967
		x"3d",	--2968
		x"ff",	--2969
		x"05",	--2970
		x"3d",	--2971
		x"00",	--2972
		x"17",	--2973
		x"3c",	--2974
		x"15",	--2975
		x"1b",	--2976
		x"02",	--2977
		x"3b",	--2978
		x"0e",	--2979
		x"0f",	--2980
		x"0a",	--2981
		x"3b",	--2982
		x"0c",	--2983
		x"0d",	--2984
		x"3c",	--2985
		x"3d",	--2986
		x"3d",	--2987
		x"ff",	--2988
		x"f5",	--2989
		x"3c",	--2990
		x"88",	--2991
		x"04",	--2992
		x"88",	--2993
		x"06",	--2994
		x"88",	--2995
		x"02",	--2996
		x"f8",	--2997
		x"03",	--2998
		x"00",	--2999
		x"0f",	--3000
		x"b3",	--3001
		x"0c",	--3002
		x"0d",	--3003
		x"1c",	--3004
		x"0d",	--3005
		x"12",	--3006
		x"0f",	--3007
		x"0e",	--3008
		x"0a",	--3009
		x"0b",	--3010
		x"0a",	--3011
		x"0b",	--3012
		x"88",	--3013
		x"04",	--3014
		x"88",	--3015
		x"06",	--3016
		x"98",	--3017
		x"02",	--3018
		x"0f",	--3019
		x"a1",	--3020
		x"6b",	--3021
		x"9f",	--3022
		x"ad",	--3023
		x"00",	--3024
		x"9d",	--3025
		x"02",	--3026
		x"02",	--3027
		x"9d",	--3028
		x"04",	--3029
		x"04",	--3030
		x"9d",	--3031
		x"06",	--3032
		x"06",	--3033
		x"5e",	--3034
		x"01",	--3035
		x"5e",	--3036
		x"01",	--3037
		x"cd",	--3038
		x"01",	--3039
		x"0f",	--3040
		x"8c",	--3041
		x"06",	--3042
		x"07",	--3043
		x"9a",	--3044
		x"39",	--3045
		x"19",	--3046
		x"39",	--3047
		x"20",	--3048
		x"8f",	--3049
		x"3e",	--3050
		x"3c",	--3051
		x"b6",	--3052
		x"c1",	--3053
		x"0e",	--3054
		x"0f",	--3055
		x"0e",	--3056
		x"0f",	--3057
		x"97",	--3058
		x"0f",	--3059
		x"79",	--3060
		x"d8",	--3061
		x"01",	--3062
		x"a8",	--3063
		x"02",	--3064
		x"3e",	--3065
		x"3f",	--3066
		x"1e",	--3067
		x"0f",	--3068
		x"88",	--3069
		x"04",	--3070
		x"88",	--3071
		x"06",	--3072
		x"92",	--3073
		x"0c",	--3074
		x"7b",	--3075
		x"81",	--3076
		x"00",	--3077
		x"81",	--3078
		x"02",	--3079
		x"81",	--3080
		x"04",	--3081
		x"4d",	--3082
		x"7d",	--3083
		x"1f",	--3084
		x"0c",	--3085
		x"4b",	--3086
		x"0c",	--3087
		x"0d",	--3088
		x"12",	--3089
		x"0d",	--3090
		x"0c",	--3091
		x"7b",	--3092
		x"fb",	--3093
		x"81",	--3094
		x"02",	--3095
		x"81",	--3096
		x"04",	--3097
		x"1c",	--3098
		x"0d",	--3099
		x"79",	--3100
		x"1f",	--3101
		x"04",	--3102
		x"0c",	--3103
		x"0d",	--3104
		x"79",	--3105
		x"fc",	--3106
		x"3c",	--3107
		x"3d",	--3108
		x"0c",	--3109
		x"0d",	--3110
		x"1a",	--3111
		x"0b",	--3112
		x"0c",	--3113
		x"04",	--3114
		x"0d",	--3115
		x"02",	--3116
		x"0a",	--3117
		x"0b",	--3118
		x"14",	--3119
		x"02",	--3120
		x"15",	--3121
		x"04",	--3122
		x"04",	--3123
		x"05",	--3124
		x"49",	--3125
		x"0a",	--3126
		x"0b",	--3127
		x"18",	--3128
		x"6c",	--3129
		x"33",	--3130
		x"df",	--3131
		x"01",	--3132
		x"01",	--3133
		x"2f",	--3134
		x"3f",	--3135
		x"90",	--3136
		x"2c",	--3137
		x"31",	--3138
		x"e0",	--3139
		x"81",	--3140
		x"04",	--3141
		x"81",	--3142
		x"06",	--3143
		x"81",	--3144
		x"00",	--3145
		x"81",	--3146
		x"02",	--3147
		x"0e",	--3148
		x"3e",	--3149
		x"18",	--3150
		x"0f",	--3151
		x"2f",	--3152
		x"b0",	--3153
		x"ec",	--3154
		x"0e",	--3155
		x"3e",	--3156
		x"10",	--3157
		x"0f",	--3158
		x"b0",	--3159
		x"ec",	--3160
		x"0d",	--3161
		x"3d",	--3162
		x"0e",	--3163
		x"3e",	--3164
		x"10",	--3165
		x"0f",	--3166
		x"3f",	--3167
		x"18",	--3168
		x"b0",	--3169
		x"f2",	--3170
		x"b0",	--3171
		x"0e",	--3172
		x"31",	--3173
		x"20",	--3174
		x"30",	--3175
		x"31",	--3176
		x"e0",	--3177
		x"81",	--3178
		x"04",	--3179
		x"81",	--3180
		x"06",	--3181
		x"81",	--3182
		x"00",	--3183
		x"81",	--3184
		x"02",	--3185
		x"0e",	--3186
		x"3e",	--3187
		x"18",	--3188
		x"0f",	--3189
		x"2f",	--3190
		x"b0",	--3191
		x"ec",	--3192
		x"0e",	--3193
		x"3e",	--3194
		x"10",	--3195
		x"0f",	--3196
		x"b0",	--3197
		x"ec",	--3198
		x"d1",	--3199
		x"11",	--3200
		x"0d",	--3201
		x"3d",	--3202
		x"0e",	--3203
		x"3e",	--3204
		x"10",	--3205
		x"0f",	--3206
		x"3f",	--3207
		x"18",	--3208
		x"b0",	--3209
		x"f2",	--3210
		x"b0",	--3211
		x"0e",	--3212
		x"31",	--3213
		x"20",	--3214
		x"30",	--3215
		x"0b",	--3216
		x"0a",	--3217
		x"09",	--3218
		x"08",	--3219
		x"07",	--3220
		x"06",	--3221
		x"05",	--3222
		x"04",	--3223
		x"31",	--3224
		x"dc",	--3225
		x"81",	--3226
		x"04",	--3227
		x"81",	--3228
		x"06",	--3229
		x"81",	--3230
		x"00",	--3231
		x"81",	--3232
		x"02",	--3233
		x"0e",	--3234
		x"3e",	--3235
		x"18",	--3236
		x"0f",	--3237
		x"2f",	--3238
		x"b0",	--3239
		x"ec",	--3240
		x"0e",	--3241
		x"3e",	--3242
		x"10",	--3243
		x"0f",	--3244
		x"b0",	--3245
		x"ec",	--3246
		x"5f",	--3247
		x"18",	--3248
		x"6f",	--3249
		x"b6",	--3250
		x"5e",	--3251
		x"10",	--3252
		x"6e",	--3253
		x"d9",	--3254
		x"6f",	--3255
		x"ae",	--3256
		x"6e",	--3257
		x"e2",	--3258
		x"6f",	--3259
		x"ac",	--3260
		x"6e",	--3261
		x"d1",	--3262
		x"14",	--3263
		x"1c",	--3264
		x"15",	--3265
		x"1e",	--3266
		x"18",	--3267
		x"14",	--3268
		x"19",	--3269
		x"16",	--3270
		x"3c",	--3271
		x"20",	--3272
		x"0e",	--3273
		x"0f",	--3274
		x"06",	--3275
		x"07",	--3276
		x"81",	--3277
		x"20",	--3278
		x"81",	--3279
		x"22",	--3280
		x"0a",	--3281
		x"0b",	--3282
		x"81",	--3283
		x"20",	--3284
		x"08",	--3285
		x"08",	--3286
		x"09",	--3287
		x"12",	--3288
		x"05",	--3289
		x"04",	--3290
		x"b1",	--3291
		x"20",	--3292
		x"19",	--3293
		x"14",	--3294
		x"0d",	--3295
		x"0a",	--3296
		x"0b",	--3297
		x"0e",	--3298
		x"0f",	--3299
		x"1c",	--3300
		x"0d",	--3301
		x"0b",	--3302
		x"03",	--3303
		x"0b",	--3304
		x"0c",	--3305
		x"0d",	--3306
		x"0e",	--3307
		x"0f",	--3308
		x"06",	--3309
		x"07",	--3310
		x"09",	--3311
		x"e5",	--3312
		x"16",	--3313
		x"07",	--3314
		x"e2",	--3315
		x"0a",	--3316
		x"f5",	--3317
		x"f2",	--3318
		x"81",	--3319
		x"20",	--3320
		x"81",	--3321
		x"22",	--3322
		x"0c",	--3323
		x"1a",	--3324
		x"1a",	--3325
		x"1a",	--3326
		x"12",	--3327
		x"06",	--3328
		x"26",	--3329
		x"81",	--3330
		x"0a",	--3331
		x"5d",	--3332
		x"d1",	--3333
		x"11",	--3334
		x"19",	--3335
		x"83",	--3336
		x"c1",	--3337
		x"09",	--3338
		x"0c",	--3339
		x"3c",	--3340
		x"3f",	--3341
		x"00",	--3342
		x"18",	--3343
		x"1d",	--3344
		x"0a",	--3345
		x"3d",	--3346
		x"1a",	--3347
		x"20",	--3348
		x"1b",	--3349
		x"22",	--3350
		x"0c",	--3351
		x"0e",	--3352
		x"0f",	--3353
		x"0b",	--3354
		x"2a",	--3355
		x"0a",	--3356
		x"0b",	--3357
		x"3d",	--3358
		x"3f",	--3359
		x"00",	--3360
		x"f5",	--3361
		x"81",	--3362
		x"20",	--3363
		x"81",	--3364
		x"22",	--3365
		x"81",	--3366
		x"0a",	--3367
		x"0c",	--3368
		x"0d",	--3369
		x"3c",	--3370
		x"7f",	--3371
		x"0d",	--3372
		x"3c",	--3373
		x"40",	--3374
		x"44",	--3375
		x"81",	--3376
		x"0c",	--3377
		x"81",	--3378
		x"0e",	--3379
		x"f1",	--3380
		x"03",	--3381
		x"08",	--3382
		x"0f",	--3383
		x"3f",	--3384
		x"b0",	--3385
		x"0e",	--3386
		x"31",	--3387
		x"24",	--3388
		x"34",	--3389
		x"35",	--3390
		x"36",	--3391
		x"37",	--3392
		x"38",	--3393
		x"39",	--3394
		x"3a",	--3395
		x"3b",	--3396
		x"30",	--3397
		x"1e",	--3398
		x"0f",	--3399
		x"d3",	--3400
		x"3a",	--3401
		x"03",	--3402
		x"08",	--3403
		x"1e",	--3404
		x"10",	--3405
		x"1c",	--3406
		x"20",	--3407
		x"1d",	--3408
		x"22",	--3409
		x"12",	--3410
		x"0d",	--3411
		x"0c",	--3412
		x"06",	--3413
		x"07",	--3414
		x"06",	--3415
		x"37",	--3416
		x"00",	--3417
		x"81",	--3418
		x"20",	--3419
		x"81",	--3420
		x"22",	--3421
		x"12",	--3422
		x"0f",	--3423
		x"0e",	--3424
		x"1a",	--3425
		x"0f",	--3426
		x"e7",	--3427
		x"81",	--3428
		x"0a",	--3429
		x"a6",	--3430
		x"6e",	--3431
		x"36",	--3432
		x"5f",	--3433
		x"d1",	--3434
		x"11",	--3435
		x"19",	--3436
		x"20",	--3437
		x"c1",	--3438
		x"19",	--3439
		x"0f",	--3440
		x"3f",	--3441
		x"18",	--3442
		x"c5",	--3443
		x"0d",	--3444
		x"ba",	--3445
		x"0c",	--3446
		x"0d",	--3447
		x"3c",	--3448
		x"80",	--3449
		x"0d",	--3450
		x"0c",	--3451
		x"b3",	--3452
		x"0d",	--3453
		x"b1",	--3454
		x"81",	--3455
		x"20",	--3456
		x"03",	--3457
		x"81",	--3458
		x"22",	--3459
		x"ab",	--3460
		x"3e",	--3461
		x"40",	--3462
		x"0f",	--3463
		x"3e",	--3464
		x"80",	--3465
		x"3f",	--3466
		x"a4",	--3467
		x"4d",	--3468
		x"7b",	--3469
		x"4f",	--3470
		x"de",	--3471
		x"5f",	--3472
		x"d1",	--3473
		x"11",	--3474
		x"19",	--3475
		x"06",	--3476
		x"c1",	--3477
		x"11",	--3478
		x"0f",	--3479
		x"3f",	--3480
		x"10",	--3481
		x"9e",	--3482
		x"4f",	--3483
		x"f8",	--3484
		x"6f",	--3485
		x"f1",	--3486
		x"3f",	--3487
		x"90",	--3488
		x"97",	--3489
		x"0b",	--3490
		x"0a",	--3491
		x"09",	--3492
		x"08",	--3493
		x"07",	--3494
		x"31",	--3495
		x"e8",	--3496
		x"81",	--3497
		x"04",	--3498
		x"81",	--3499
		x"06",	--3500
		x"81",	--3501
		x"00",	--3502
		x"81",	--3503
		x"02",	--3504
		x"0e",	--3505
		x"3e",	--3506
		x"10",	--3507
		x"0f",	--3508
		x"2f",	--3509
		x"b0",	--3510
		x"ec",	--3511
		x"0e",	--3512
		x"3e",	--3513
		x"0f",	--3514
		x"b0",	--3515
		x"ec",	--3516
		x"5f",	--3517
		x"10",	--3518
		x"6f",	--3519
		x"5d",	--3520
		x"5e",	--3521
		x"08",	--3522
		x"6e",	--3523
		x"82",	--3524
		x"d1",	--3525
		x"09",	--3526
		x"11",	--3527
		x"6f",	--3528
		x"58",	--3529
		x"6f",	--3530
		x"56",	--3531
		x"6e",	--3532
		x"6f",	--3533
		x"6e",	--3534
		x"4c",	--3535
		x"1d",	--3536
		x"12",	--3537
		x"1d",	--3538
		x"0a",	--3539
		x"81",	--3540
		x"12",	--3541
		x"1e",	--3542
		x"14",	--3543
		x"1f",	--3544
		x"16",	--3545
		x"18",	--3546
		x"0c",	--3547
		x"19",	--3548
		x"0e",	--3549
		x"0f",	--3550
		x"1e",	--3551
		x"0e",	--3552
		x"0f",	--3553
		x"3d",	--3554
		x"81",	--3555
		x"12",	--3556
		x"37",	--3557
		x"1f",	--3558
		x"0c",	--3559
		x"3d",	--3560
		x"00",	--3561
		x"0a",	--3562
		x"0b",	--3563
		x"0b",	--3564
		x"0a",	--3565
		x"0b",	--3566
		x"0e",	--3567
		x"0f",	--3568
		x"12",	--3569
		x"0d",	--3570
		x"0c",	--3571
		x"0e",	--3572
		x"0f",	--3573
		x"37",	--3574
		x"0b",	--3575
		x"0f",	--3576
		x"f7",	--3577
		x"f2",	--3578
		x"0e",	--3579
		x"f4",	--3580
		x"ef",	--3581
		x"09",	--3582
		x"e5",	--3583
		x"0e",	--3584
		x"e3",	--3585
		x"dd",	--3586
		x"0c",	--3587
		x"0d",	--3588
		x"3c",	--3589
		x"7f",	--3590
		x"0d",	--3591
		x"3c",	--3592
		x"40",	--3593
		x"1c",	--3594
		x"81",	--3595
		x"14",	--3596
		x"81",	--3597
		x"16",	--3598
		x"0f",	--3599
		x"3f",	--3600
		x"10",	--3601
		x"b0",	--3602
		x"0e",	--3603
		x"31",	--3604
		x"18",	--3605
		x"37",	--3606
		x"38",	--3607
		x"39",	--3608
		x"3a",	--3609
		x"3b",	--3610
		x"30",	--3611
		x"e1",	--3612
		x"10",	--3613
		x"0f",	--3614
		x"3f",	--3615
		x"10",	--3616
		x"f0",	--3617
		x"4f",	--3618
		x"fa",	--3619
		x"3f",	--3620
		x"90",	--3621
		x"eb",	--3622
		x"0d",	--3623
		x"e2",	--3624
		x"0c",	--3625
		x"0d",	--3626
		x"3c",	--3627
		x"80",	--3628
		x"0d",	--3629
		x"0c",	--3630
		x"db",	--3631
		x"0d",	--3632
		x"d9",	--3633
		x"0e",	--3634
		x"02",	--3635
		x"0f",	--3636
		x"d5",	--3637
		x"3a",	--3638
		x"40",	--3639
		x"0b",	--3640
		x"3a",	--3641
		x"80",	--3642
		x"3b",	--3643
		x"ce",	--3644
		x"81",	--3645
		x"14",	--3646
		x"81",	--3647
		x"16",	--3648
		x"81",	--3649
		x"12",	--3650
		x"0f",	--3651
		x"3f",	--3652
		x"10",	--3653
		x"cb",	--3654
		x"0f",	--3655
		x"3f",	--3656
		x"c8",	--3657
		x"31",	--3658
		x"e8",	--3659
		x"81",	--3660
		x"04",	--3661
		x"81",	--3662
		x"06",	--3663
		x"81",	--3664
		x"00",	--3665
		x"81",	--3666
		x"02",	--3667
		x"0e",	--3668
		x"3e",	--3669
		x"10",	--3670
		x"0f",	--3671
		x"2f",	--3672
		x"b0",	--3673
		x"ec",	--3674
		x"0e",	--3675
		x"3e",	--3676
		x"0f",	--3677
		x"b0",	--3678
		x"ec",	--3679
		x"e1",	--3680
		x"10",	--3681
		x"0d",	--3682
		x"e1",	--3683
		x"08",	--3684
		x"0a",	--3685
		x"0e",	--3686
		x"3e",	--3687
		x"0f",	--3688
		x"3f",	--3689
		x"10",	--3690
		x"b0",	--3691
		x"10",	--3692
		x"31",	--3693
		x"18",	--3694
		x"30",	--3695
		x"3f",	--3696
		x"fb",	--3697
		x"31",	--3698
		x"e8",	--3699
		x"81",	--3700
		x"04",	--3701
		x"81",	--3702
		x"06",	--3703
		x"81",	--3704
		x"00",	--3705
		x"81",	--3706
		x"02",	--3707
		x"0e",	--3708
		x"3e",	--3709
		x"10",	--3710
		x"0f",	--3711
		x"2f",	--3712
		x"b0",	--3713
		x"ec",	--3714
		x"0e",	--3715
		x"3e",	--3716
		x"0f",	--3717
		x"b0",	--3718
		x"ec",	--3719
		x"e1",	--3720
		x"10",	--3721
		x"0d",	--3722
		x"e1",	--3723
		x"08",	--3724
		x"0a",	--3725
		x"0e",	--3726
		x"3e",	--3727
		x"0f",	--3728
		x"3f",	--3729
		x"10",	--3730
		x"b0",	--3731
		x"10",	--3732
		x"31",	--3733
		x"18",	--3734
		x"30",	--3735
		x"3f",	--3736
		x"fb",	--3737
		x"31",	--3738
		x"e8",	--3739
		x"81",	--3740
		x"04",	--3741
		x"81",	--3742
		x"06",	--3743
		x"81",	--3744
		x"00",	--3745
		x"81",	--3746
		x"02",	--3747
		x"0e",	--3748
		x"3e",	--3749
		x"10",	--3750
		x"0f",	--3751
		x"2f",	--3752
		x"b0",	--3753
		x"ec",	--3754
		x"0e",	--3755
		x"3e",	--3756
		x"0f",	--3757
		x"b0",	--3758
		x"ec",	--3759
		x"e1",	--3760
		x"10",	--3761
		x"0d",	--3762
		x"e1",	--3763
		x"08",	--3764
		x"0a",	--3765
		x"0e",	--3766
		x"3e",	--3767
		x"0f",	--3768
		x"3f",	--3769
		x"10",	--3770
		x"b0",	--3771
		x"10",	--3772
		x"31",	--3773
		x"18",	--3774
		x"30",	--3775
		x"1f",	--3776
		x"fb",	--3777
		x"0b",	--3778
		x"0a",	--3779
		x"31",	--3780
		x"f1",	--3781
		x"03",	--3782
		x"00",	--3783
		x"0d",	--3784
		x"0d",	--3785
		x"0d",	--3786
		x"0d",	--3787
		x"4c",	--3788
		x"c1",	--3789
		x"01",	--3790
		x"0e",	--3791
		x"0b",	--3792
		x"0f",	--3793
		x"09",	--3794
		x"e1",	--3795
		x"00",	--3796
		x"0f",	--3797
		x"b0",	--3798
		x"0e",	--3799
		x"31",	--3800
		x"3a",	--3801
		x"3b",	--3802
		x"30",	--3803
		x"b1",	--3804
		x"1e",	--3805
		x"02",	--3806
		x"4c",	--3807
		x"1b",	--3808
		x"0a",	--3809
		x"0b",	--3810
		x"81",	--3811
		x"04",	--3812
		x"81",	--3813
		x"06",	--3814
		x"0e",	--3815
		x"0f",	--3816
		x"b0",	--3817
		x"9c",	--3818
		x"3f",	--3819
		x"1f",	--3820
		x"e7",	--3821
		x"81",	--3822
		x"04",	--3823
		x"81",	--3824
		x"06",	--3825
		x"4e",	--3826
		x"7e",	--3827
		x"1f",	--3828
		x"0f",	--3829
		x"3e",	--3830
		x"1e",	--3831
		x"0e",	--3832
		x"81",	--3833
		x"02",	--3834
		x"d9",	--3835
		x"0e",	--3836
		x"10",	--3837
		x"0a",	--3838
		x"0b",	--3839
		x"3a",	--3840
		x"3b",	--3841
		x"1a",	--3842
		x"0b",	--3843
		x"de",	--3844
		x"91",	--3845
		x"04",	--3846
		x"04",	--3847
		x"91",	--3848
		x"06",	--3849
		x"06",	--3850
		x"7e",	--3851
		x"f8",	--3852
		x"e8",	--3853
		x"3f",	--3854
		x"00",	--3855
		x"ed",	--3856
		x"0e",	--3857
		x"3f",	--3858
		x"00",	--3859
		x"c3",	--3860
		x"31",	--3861
		x"f4",	--3862
		x"81",	--3863
		x"00",	--3864
		x"81",	--3865
		x"02",	--3866
		x"0e",	--3867
		x"2e",	--3868
		x"0f",	--3869
		x"b0",	--3870
		x"ec",	--3871
		x"5f",	--3872
		x"04",	--3873
		x"6f",	--3874
		x"28",	--3875
		x"27",	--3876
		x"6f",	--3877
		x"07",	--3878
		x"1d",	--3879
		x"06",	--3880
		x"0d",	--3881
		x"21",	--3882
		x"3d",	--3883
		x"1f",	--3884
		x"09",	--3885
		x"c1",	--3886
		x"05",	--3887
		x"26",	--3888
		x"3e",	--3889
		x"3f",	--3890
		x"ff",	--3891
		x"31",	--3892
		x"0c",	--3893
		x"30",	--3894
		x"1e",	--3895
		x"08",	--3896
		x"1f",	--3897
		x"0a",	--3898
		x"3c",	--3899
		x"1e",	--3900
		x"4c",	--3901
		x"4d",	--3902
		x"7d",	--3903
		x"1f",	--3904
		x"0f",	--3905
		x"c1",	--3906
		x"05",	--3907
		x"ef",	--3908
		x"3e",	--3909
		x"3f",	--3910
		x"1e",	--3911
		x"0f",	--3912
		x"31",	--3913
		x"0c",	--3914
		x"30",	--3915
		x"0e",	--3916
		x"0f",	--3917
		x"31",	--3918
		x"0c",	--3919
		x"30",	--3920
		x"12",	--3921
		x"0f",	--3922
		x"0e",	--3923
		x"7d",	--3924
		x"fb",	--3925
		x"eb",	--3926
		x"0e",	--3927
		x"3f",	--3928
		x"00",	--3929
		x"31",	--3930
		x"0c",	--3931
		x"30",	--3932
		x"0b",	--3933
		x"0a",	--3934
		x"09",	--3935
		x"08",	--3936
		x"31",	--3937
		x"0a",	--3938
		x"0b",	--3939
		x"c1",	--3940
		x"01",	--3941
		x"0e",	--3942
		x"0d",	--3943
		x"0b",	--3944
		x"0b",	--3945
		x"e1",	--3946
		x"00",	--3947
		x"0f",	--3948
		x"b0",	--3949
		x"0e",	--3950
		x"31",	--3951
		x"38",	--3952
		x"39",	--3953
		x"3a",	--3954
		x"3b",	--3955
		x"30",	--3956
		x"f1",	--3957
		x"03",	--3958
		x"00",	--3959
		x"b1",	--3960
		x"1e",	--3961
		x"02",	--3962
		x"81",	--3963
		x"04",	--3964
		x"81",	--3965
		x"06",	--3966
		x"0e",	--3967
		x"0f",	--3968
		x"b0",	--3969
		x"9c",	--3970
		x"3f",	--3971
		x"0f",	--3972
		x"18",	--3973
		x"e5",	--3974
		x"81",	--3975
		x"04",	--3976
		x"81",	--3977
		x"06",	--3978
		x"4e",	--3979
		x"7e",	--3980
		x"1f",	--3981
		x"06",	--3982
		x"3e",	--3983
		x"1e",	--3984
		x"0e",	--3985
		x"81",	--3986
		x"02",	--3987
		x"d7",	--3988
		x"91",	--3989
		x"04",	--3990
		x"04",	--3991
		x"91",	--3992
		x"06",	--3993
		x"06",	--3994
		x"7e",	--3995
		x"f8",	--3996
		x"f1",	--3997
		x"0e",	--3998
		x"3e",	--3999
		x"1e",	--4000
		x"1c",	--4001
		x"0d",	--4002
		x"48",	--4003
		x"78",	--4004
		x"1f",	--4005
		x"04",	--4006
		x"0c",	--4007
		x"0d",	--4008
		x"78",	--4009
		x"fc",	--4010
		x"3c",	--4011
		x"3d",	--4012
		x"0c",	--4013
		x"0d",	--4014
		x"18",	--4015
		x"09",	--4016
		x"0c",	--4017
		x"04",	--4018
		x"0d",	--4019
		x"02",	--4020
		x"08",	--4021
		x"09",	--4022
		x"7e",	--4023
		x"1f",	--4024
		x"0e",	--4025
		x"0d",	--4026
		x"0e",	--4027
		x"0d",	--4028
		x"0e",	--4029
		x"81",	--4030
		x"04",	--4031
		x"81",	--4032
		x"06",	--4033
		x"3e",	--4034
		x"1e",	--4035
		x"0e",	--4036
		x"81",	--4037
		x"02",	--4038
		x"a4",	--4039
		x"12",	--4040
		x"0b",	--4041
		x"0a",	--4042
		x"7e",	--4043
		x"fb",	--4044
		x"ec",	--4045
		x"0b",	--4046
		x"0a",	--4047
		x"09",	--4048
		x"1f",	--4049
		x"17",	--4050
		x"3e",	--4051
		x"00",	--4052
		x"2c",	--4053
		x"3a",	--4054
		x"18",	--4055
		x"0b",	--4056
		x"39",	--4057
		x"0c",	--4058
		x"0d",	--4059
		x"4f",	--4060
		x"4f",	--4061
		x"17",	--4062
		x"3c",	--4063
		x"98",	--4064
		x"6e",	--4065
		x"0f",	--4066
		x"0a",	--4067
		x"0b",	--4068
		x"0f",	--4069
		x"39",	--4070
		x"3a",	--4071
		x"3b",	--4072
		x"30",	--4073
		x"3f",	--4074
		x"00",	--4075
		x"0f",	--4076
		x"3a",	--4077
		x"0b",	--4078
		x"39",	--4079
		x"18",	--4080
		x"0c",	--4081
		x"0d",	--4082
		x"4f",	--4083
		x"4f",	--4084
		x"e9",	--4085
		x"12",	--4086
		x"0d",	--4087
		x"0c",	--4088
		x"7f",	--4089
		x"fb",	--4090
		x"e3",	--4091
		x"3a",	--4092
		x"10",	--4093
		x"0b",	--4094
		x"39",	--4095
		x"10",	--4096
		x"ef",	--4097
		x"3a",	--4098
		x"20",	--4099
		x"0b",	--4100
		x"09",	--4101
		x"ea",	--4102
		x"0b",	--4103
		x"0a",	--4104
		x"09",	--4105
		x"08",	--4106
		x"07",	--4107
		x"0d",	--4108
		x"1e",	--4109
		x"04",	--4110
		x"1f",	--4111
		x"06",	--4112
		x"5a",	--4113
		x"01",	--4114
		x"6c",	--4115
		x"6c",	--4116
		x"70",	--4117
		x"6c",	--4118
		x"6a",	--4119
		x"6c",	--4120
		x"36",	--4121
		x"0e",	--4122
		x"32",	--4123
		x"1b",	--4124
		x"02",	--4125
		x"3b",	--4126
		x"82",	--4127
		x"6d",	--4128
		x"3b",	--4129
		x"80",	--4130
		x"5e",	--4131
		x"0c",	--4132
		x"0d",	--4133
		x"3c",	--4134
		x"7f",	--4135
		x"0d",	--4136
		x"3c",	--4137
		x"40",	--4138
		x"40",	--4139
		x"3e",	--4140
		x"3f",	--4141
		x"0f",	--4142
		x"0f",	--4143
		x"4a",	--4144
		x"0d",	--4145
		x"3d",	--4146
		x"7f",	--4147
		x"12",	--4148
		x"0f",	--4149
		x"0e",	--4150
		x"12",	--4151
		x"0f",	--4152
		x"0e",	--4153
		x"12",	--4154
		x"0f",	--4155
		x"0e",	--4156
		x"12",	--4157
		x"0f",	--4158
		x"0e",	--4159
		x"12",	--4160
		x"0f",	--4161
		x"0e",	--4162
		x"12",	--4163
		x"0f",	--4164
		x"0e",	--4165
		x"12",	--4166
		x"0f",	--4167
		x"0e",	--4168
		x"3e",	--4169
		x"3f",	--4170
		x"7f",	--4171
		x"4d",	--4172
		x"05",	--4173
		x"0f",	--4174
		x"cc",	--4175
		x"4d",	--4176
		x"0e",	--4177
		x"0f",	--4178
		x"4d",	--4179
		x"0d",	--4180
		x"0d",	--4181
		x"0d",	--4182
		x"0d",	--4183
		x"0d",	--4184
		x"0d",	--4185
		x"0d",	--4186
		x"0c",	--4187
		x"3c",	--4188
		x"7f",	--4189
		x"0c",	--4190
		x"4f",	--4191
		x"0f",	--4192
		x"0f",	--4193
		x"0f",	--4194
		x"0d",	--4195
		x"0d",	--4196
		x"0f",	--4197
		x"37",	--4198
		x"38",	--4199
		x"39",	--4200
		x"3a",	--4201
		x"3b",	--4202
		x"30",	--4203
		x"0d",	--4204
		x"be",	--4205
		x"0c",	--4206
		x"0d",	--4207
		x"3c",	--4208
		x"80",	--4209
		x"0d",	--4210
		x"0c",	--4211
		x"02",	--4212
		x"0d",	--4213
		x"b8",	--4214
		x"3e",	--4215
		x"40",	--4216
		x"0f",	--4217
		x"b4",	--4218
		x"12",	--4219
		x"0f",	--4220
		x"0e",	--4221
		x"0d",	--4222
		x"3d",	--4223
		x"80",	--4224
		x"b2",	--4225
		x"7d",	--4226
		x"0e",	--4227
		x"0f",	--4228
		x"cd",	--4229
		x"0e",	--4230
		x"3f",	--4231
		x"10",	--4232
		x"3e",	--4233
		x"3f",	--4234
		x"7f",	--4235
		x"7d",	--4236
		x"c5",	--4237
		x"37",	--4238
		x"82",	--4239
		x"07",	--4240
		x"37",	--4241
		x"1a",	--4242
		x"4f",	--4243
		x"0c",	--4244
		x"0d",	--4245
		x"4b",	--4246
		x"7b",	--4247
		x"1f",	--4248
		x"05",	--4249
		x"12",	--4250
		x"0d",	--4251
		x"0c",	--4252
		x"7b",	--4253
		x"fb",	--4254
		x"18",	--4255
		x"09",	--4256
		x"77",	--4257
		x"1f",	--4258
		x"04",	--4259
		x"08",	--4260
		x"09",	--4261
		x"77",	--4262
		x"fc",	--4263
		x"38",	--4264
		x"39",	--4265
		x"08",	--4266
		x"09",	--4267
		x"1e",	--4268
		x"0f",	--4269
		x"08",	--4270
		x"04",	--4271
		x"09",	--4272
		x"02",	--4273
		x"0e",	--4274
		x"0f",	--4275
		x"08",	--4276
		x"09",	--4277
		x"08",	--4278
		x"09",	--4279
		x"0e",	--4280
		x"0f",	--4281
		x"3e",	--4282
		x"7f",	--4283
		x"0f",	--4284
		x"3e",	--4285
		x"40",	--4286
		x"26",	--4287
		x"38",	--4288
		x"3f",	--4289
		x"09",	--4290
		x"0e",	--4291
		x"0f",	--4292
		x"12",	--4293
		x"0f",	--4294
		x"0e",	--4295
		x"12",	--4296
		x"0f",	--4297
		x"0e",	--4298
		x"12",	--4299
		x"0f",	--4300
		x"0e",	--4301
		x"12",	--4302
		x"0f",	--4303
		x"0e",	--4304
		x"12",	--4305
		x"0f",	--4306
		x"0e",	--4307
		x"12",	--4308
		x"0f",	--4309
		x"0e",	--4310
		x"12",	--4311
		x"0f",	--4312
		x"0e",	--4313
		x"3e",	--4314
		x"3f",	--4315
		x"7f",	--4316
		x"5d",	--4317
		x"39",	--4318
		x"00",	--4319
		x"72",	--4320
		x"4d",	--4321
		x"70",	--4322
		x"08",	--4323
		x"09",	--4324
		x"da",	--4325
		x"0f",	--4326
		x"d8",	--4327
		x"0e",	--4328
		x"0f",	--4329
		x"3e",	--4330
		x"80",	--4331
		x"0f",	--4332
		x"0e",	--4333
		x"04",	--4334
		x"38",	--4335
		x"40",	--4336
		x"09",	--4337
		x"d0",	--4338
		x"0f",	--4339
		x"ce",	--4340
		x"f9",	--4341
		x"0b",	--4342
		x"0a",	--4343
		x"2a",	--4344
		x"5b",	--4345
		x"02",	--4346
		x"3b",	--4347
		x"7f",	--4348
		x"1d",	--4349
		x"02",	--4350
		x"12",	--4351
		x"0d",	--4352
		x"12",	--4353
		x"0d",	--4354
		x"12",	--4355
		x"0d",	--4356
		x"12",	--4357
		x"0d",	--4358
		x"12",	--4359
		x"0d",	--4360
		x"12",	--4361
		x"0d",	--4362
		x"12",	--4363
		x"0d",	--4364
		x"4d",	--4365
		x"5f",	--4366
		x"03",	--4367
		x"3f",	--4368
		x"80",	--4369
		x"0f",	--4370
		x"0f",	--4371
		x"ce",	--4372
		x"01",	--4373
		x"0d",	--4374
		x"2d",	--4375
		x"0a",	--4376
		x"51",	--4377
		x"be",	--4378
		x"82",	--4379
		x"02",	--4380
		x"0c",	--4381
		x"0d",	--4382
		x"0c",	--4383
		x"0d",	--4384
		x"0c",	--4385
		x"0d",	--4386
		x"0c",	--4387
		x"0d",	--4388
		x"0c",	--4389
		x"0d",	--4390
		x"0c",	--4391
		x"0d",	--4392
		x"0c",	--4393
		x"0d",	--4394
		x"0c",	--4395
		x"0d",	--4396
		x"fe",	--4397
		x"03",	--4398
		x"00",	--4399
		x"3d",	--4400
		x"00",	--4401
		x"0b",	--4402
		x"3f",	--4403
		x"81",	--4404
		x"0c",	--4405
		x"0d",	--4406
		x"0a",	--4407
		x"3f",	--4408
		x"3d",	--4409
		x"00",	--4410
		x"f9",	--4411
		x"8e",	--4412
		x"02",	--4413
		x"8e",	--4414
		x"04",	--4415
		x"8e",	--4416
		x"06",	--4417
		x"3a",	--4418
		x"3b",	--4419
		x"30",	--4420
		x"3d",	--4421
		x"ff",	--4422
		x"2a",	--4423
		x"3d",	--4424
		x"81",	--4425
		x"8e",	--4426
		x"02",	--4427
		x"fe",	--4428
		x"03",	--4429
		x"00",	--4430
		x"0c",	--4431
		x"0d",	--4432
		x"0c",	--4433
		x"0d",	--4434
		x"0c",	--4435
		x"0d",	--4436
		x"0c",	--4437
		x"0d",	--4438
		x"0c",	--4439
		x"0d",	--4440
		x"0c",	--4441
		x"0d",	--4442
		x"0c",	--4443
		x"0d",	--4444
		x"0c",	--4445
		x"0d",	--4446
		x"0a",	--4447
		x"0b",	--4448
		x"0a",	--4449
		x"3b",	--4450
		x"00",	--4451
		x"8e",	--4452
		x"04",	--4453
		x"8e",	--4454
		x"06",	--4455
		x"3a",	--4456
		x"3b",	--4457
		x"30",	--4458
		x"0b",	--4459
		x"ad",	--4460
		x"ee",	--4461
		x"00",	--4462
		x"3a",	--4463
		x"3b",	--4464
		x"30",	--4465
		x"0a",	--4466
		x"0c",	--4467
		x"0c",	--4468
		x"0d",	--4469
		x"0c",	--4470
		x"3d",	--4471
		x"10",	--4472
		x"0c",	--4473
		x"02",	--4474
		x"0d",	--4475
		x"08",	--4476
		x"de",	--4477
		x"00",	--4478
		x"e4",	--4479
		x"0b",	--4480
		x"f2",	--4481
		x"ee",	--4482
		x"00",	--4483
		x"e3",	--4484
		x"ce",	--4485
		x"00",	--4486
		x"dc",	--4487
		x"0b",	--4488
		x"6d",	--4489
		x"6d",	--4490
		x"12",	--4491
		x"6c",	--4492
		x"6c",	--4493
		x"0f",	--4494
		x"6d",	--4495
		x"41",	--4496
		x"6c",	--4497
		x"11",	--4498
		x"6d",	--4499
		x"0d",	--4500
		x"6c",	--4501
		x"14",	--4502
		x"5d",	--4503
		x"01",	--4504
		x"5d",	--4505
		x"01",	--4506
		x"14",	--4507
		x"4d",	--4508
		x"09",	--4509
		x"1e",	--4510
		x"0f",	--4511
		x"3b",	--4512
		x"30",	--4513
		x"6c",	--4514
		x"28",	--4515
		x"ce",	--4516
		x"01",	--4517
		x"f7",	--4518
		x"3e",	--4519
		x"0f",	--4520
		x"3b",	--4521
		x"30",	--4522
		x"cf",	--4523
		x"01",	--4524
		x"f0",	--4525
		x"3e",	--4526
		x"f8",	--4527
		x"1b",	--4528
		x"02",	--4529
		x"1c",	--4530
		x"02",	--4531
		x"0c",	--4532
		x"e6",	--4533
		x"0b",	--4534
		x"16",	--4535
		x"1b",	--4536
		x"04",	--4537
		x"1f",	--4538
		x"06",	--4539
		x"1c",	--4540
		x"04",	--4541
		x"1e",	--4542
		x"06",	--4543
		x"0e",	--4544
		x"da",	--4545
		x"0f",	--4546
		x"02",	--4547
		x"0c",	--4548
		x"d6",	--4549
		x"0f",	--4550
		x"06",	--4551
		x"0e",	--4552
		x"02",	--4553
		x"0b",	--4554
		x"02",	--4555
		x"0e",	--4556
		x"d1",	--4557
		x"4d",	--4558
		x"ce",	--4559
		x"3e",	--4560
		x"d6",	--4561
		x"6c",	--4562
		x"d7",	--4563
		x"5e",	--4564
		x"01",	--4565
		x"5f",	--4566
		x"01",	--4567
		x"0e",	--4568
		x"c5",	--4569
		x"1e",	--4570
		x"22",	--4571
		x"1e",	--4572
		x"0b",	--4573
		x"1d",	--4574
		x"20",	--4575
		x"cd",	--4576
		x"00",	--4577
		x"1d",	--4578
		x"82",	--4579
		x"20",	--4580
		x"3e",	--4581
		x"82",	--4582
		x"22",	--4583
		x"30",	--4584
		x"3f",	--4585
		x"30",	--4586
		x"0b",	--4587
		x"0a",	--4588
		x"21",	--4589
		x"81",	--4590
		x"00",	--4591
		x"1a",	--4592
		x"20",	--4593
		x"1b",	--4594
		x"22",	--4595
		x"0d",	--4596
		x"0e",	--4597
		x"3f",	--4598
		x"b4",	--4599
		x"b0",	--4600
		x"08",	--4601
		x"0f",	--4602
		x"05",	--4603
		x"0e",	--4604
		x"0e",	--4605
		x"ce",	--4606
		x"ff",	--4607
		x"04",	--4608
		x"1e",	--4609
		x"20",	--4610
		x"ce",	--4611
		x"00",	--4612
		x"21",	--4613
		x"3a",	--4614
		x"3b",	--4615
		x"30",	--4616
		x"92",	--4617
		x"02",	--4618
		x"20",	--4619
		x"b2",	--4620
		x"ff",	--4621
		x"22",	--4622
		x"0e",	--4623
		x"3e",	--4624
		x"06",	--4625
		x"1f",	--4626
		x"04",	--4627
		x"b0",	--4628
		x"d6",	--4629
		x"30",	--4630
		x"92",	--4631
		x"02",	--4632
		x"20",	--4633
		x"92",	--4634
		x"04",	--4635
		x"22",	--4636
		x"0e",	--4637
		x"3e",	--4638
		x"1f",	--4639
		x"06",	--4640
		x"b0",	--4641
		x"d6",	--4642
		x"30",	--4643
		x"0c",	--4644
		x"82",	--4645
		x"20",	--4646
		x"b2",	--4647
		x"ff",	--4648
		x"22",	--4649
		x"0e",	--4650
		x"0f",	--4651
		x"b0",	--4652
		x"d6",	--4653
		x"30",	--4654
		x"82",	--4655
		x"20",	--4656
		x"82",	--4657
		x"22",	--4658
		x"0e",	--4659
		x"0f",	--4660
		x"b0",	--4661
		x"d6",	--4662
		x"30",	--4663
		x"0b",	--4664
		x"0a",	--4665
		x"09",	--4666
		x"08",	--4667
		x"07",	--4668
		x"06",	--4669
		x"05",	--4670
		x"04",	--4671
		x"31",	--4672
		x"08",	--4673
		x"81",	--4674
		x"04",	--4675
		x"09",	--4676
		x"1f",	--4677
		x"1a",	--4678
		x"1d",	--4679
		x"1c",	--4680
		x"4c",	--4681
		x"04",	--4682
		x"84",	--4683
		x"45",	--4684
		x"4e",	--4685
		x"7e",	--4686
		x"40",	--4687
		x"11",	--4688
		x"f1",	--4689
		x"30",	--4690
		x"00",	--4691
		x"0e",	--4692
		x"8e",	--4693
		x"5e",	--4694
		x"03",	--4695
		x"7e",	--4696
		x"58",	--4697
		x"02",	--4698
		x"7e",	--4699
		x"78",	--4700
		x"c1",	--4701
		x"01",	--4702
		x"0c",	--4703
		x"2c",	--4704
		x"0f",	--4705
		x"7e",	--4706
		x"20",	--4707
		x"04",	--4708
		x"f1",	--4709
		x"30",	--4710
		x"00",	--4711
		x"04",	--4712
		x"4c",	--4713
		x"05",	--4714
		x"c1",	--4715
		x"00",	--4716
		x"0c",	--4717
		x"1c",	--4718
		x"01",	--4719
		x"0c",	--4720
		x"0a",	--4721
		x"8c",	--4722
		x"8c",	--4723
		x"8c",	--4724
		x"8c",	--4725
		x"0b",	--4726
		x"06",	--4727
		x"0c",	--4728
		x"8c",	--4729
		x"8c",	--4730
		x"8c",	--4731
		x"8c",	--4732
		x"07",	--4733
		x"0a",	--4734
		x"0b",	--4735
		x"0e",	--4736
		x"8e",	--4737
		x"c1",	--4738
		x"02",	--4739
		x"6e",	--4740
		x"02",	--4741
		x"07",	--4742
		x"01",	--4743
		x"37",	--4744
		x"4f",	--4745
		x"7f",	--4746
		x"10",	--4747
		x"3c",	--4748
		x"1d",	--4749
		x"04",	--4750
		x"3d",	--4751
		x"1d",	--4752
		x"cd",	--4753
		x"00",	--4754
		x"fc",	--4755
		x"1d",	--4756
		x"04",	--4757
		x"09",	--4758
		x"02",	--4759
		x"09",	--4760
		x"01",	--4761
		x"09",	--4762
		x"e1",	--4763
		x"02",	--4764
		x"05",	--4765
		x"09",	--4766
		x"02",	--4767
		x"09",	--4768
		x"01",	--4769
		x"09",	--4770
		x"05",	--4771
		x"07",	--4772
		x"01",	--4773
		x"05",	--4774
		x"4f",	--4775
		x"0d",	--4776
		x"f1",	--4777
		x"20",	--4778
		x"06",	--4779
		x"06",	--4780
		x"0b",	--4781
		x"0e",	--4782
		x"0f",	--4783
		x"0f",	--4784
		x"6f",	--4785
		x"8f",	--4786
		x"16",	--4787
		x"88",	--4788
		x"01",	--4789
		x"06",	--4790
		x"06",	--4791
		x"f6",	--4792
		x"0b",	--4793
		x"f1",	--4794
		x"30",	--4795
		x"06",	--4796
		x"05",	--4797
		x"05",	--4798
		x"5f",	--4799
		x"06",	--4800
		x"8f",	--4801
		x"88",	--4802
		x"1b",	--4803
		x"0f",	--4804
		x"0f",	--4805
		x"0f",	--4806
		x"f7",	--4807
		x"0a",	--4808
		x"06",	--4809
		x"0b",	--4810
		x"07",	--4811
		x"1b",	--4812
		x"0f",	--4813
		x"0f",	--4814
		x"6f",	--4815
		x"8f",	--4816
		x"16",	--4817
		x"88",	--4818
		x"06",	--4819
		x"f7",	--4820
		x"e1",	--4821
		x"02",	--4822
		x"02",	--4823
		x"4a",	--4824
		x"08",	--4825
		x"1a",	--4826
		x"04",	--4827
		x"0a",	--4828
		x"0d",	--4829
		x"3f",	--4830
		x"30",	--4831
		x"88",	--4832
		x"7a",	--4833
		x"4a",	--4834
		x"fa",	--4835
		x"44",	--4836
		x"0b",	--4837
		x"f3",	--4838
		x"37",	--4839
		x"8f",	--4840
		x"88",	--4841
		x"1b",	--4842
		x"0f",	--4843
		x"0f",	--4844
		x"6f",	--4845
		x"4f",	--4846
		x"07",	--4847
		x"07",	--4848
		x"f5",	--4849
		x"04",	--4850
		x"3f",	--4851
		x"20",	--4852
		x"88",	--4853
		x"1b",	--4854
		x"0b",	--4855
		x"fa",	--4856
		x"0f",	--4857
		x"31",	--4858
		x"34",	--4859
		x"35",	--4860
		x"36",	--4861
		x"37",	--4862
		x"38",	--4863
		x"39",	--4864
		x"3a",	--4865
		x"3b",	--4866
		x"30",	--4867
		x"0b",	--4868
		x"0a",	--4869
		x"09",	--4870
		x"08",	--4871
		x"07",	--4872
		x"06",	--4873
		x"05",	--4874
		x"04",	--4875
		x"31",	--4876
		x"b6",	--4877
		x"81",	--4878
		x"3a",	--4879
		x"06",	--4880
		x"05",	--4881
		x"81",	--4882
		x"3e",	--4883
		x"c1",	--4884
		x"2f",	--4885
		x"c1",	--4886
		x"2b",	--4887
		x"c1",	--4888
		x"2e",	--4889
		x"c1",	--4890
		x"2a",	--4891
		x"81",	--4892
		x"30",	--4893
		x"81",	--4894
		x"26",	--4895
		x"07",	--4896
		x"81",	--4897
		x"2c",	--4898
		x"0e",	--4899
		x"3e",	--4900
		x"1c",	--4901
		x"81",	--4902
		x"1c",	--4903
		x"30",	--4904
		x"82",	--4905
		x"0f",	--4906
		x"1f",	--4907
		x"81",	--4908
		x"40",	--4909
		x"07",	--4910
		x"1e",	--4911
		x"7e",	--4912
		x"25",	--4913
		x"13",	--4914
		x"81",	--4915
		x"00",	--4916
		x"81",	--4917
		x"02",	--4918
		x"81",	--4919
		x"3e",	--4920
		x"c1",	--4921
		x"2f",	--4922
		x"c1",	--4923
		x"2b",	--4924
		x"c1",	--4925
		x"2e",	--4926
		x"c1",	--4927
		x"2a",	--4928
		x"81",	--4929
		x"30",	--4930
		x"30",	--4931
		x"78",	--4932
		x"05",	--4933
		x"8e",	--4934
		x"0f",	--4935
		x"91",	--4936
		x"3c",	--4937
		x"91",	--4938
		x"2c",	--4939
		x"30",	--4940
		x"5e",	--4941
		x"7e",	--4942
		x"63",	--4943
		x"c5",	--4944
		x"7e",	--4945
		x"64",	--4946
		x"27",	--4947
		x"7e",	--4948
		x"30",	--4949
		x"94",	--4950
		x"7e",	--4951
		x"31",	--4952
		x"1a",	--4953
		x"7e",	--4954
		x"2a",	--4955
		x"77",	--4956
		x"7e",	--4957
		x"2b",	--4958
		x"0a",	--4959
		x"7e",	--4960
		x"23",	--4961
		x"42",	--4962
		x"7e",	--4963
		x"25",	--4964
		x"e0",	--4965
		x"7e",	--4966
		x"20",	--4967
		x"32",	--4968
		x"56",	--4969
		x"7e",	--4970
		x"2d",	--4971
		x"49",	--4972
		x"7e",	--4973
		x"2e",	--4974
		x"5b",	--4975
		x"7e",	--4976
		x"2b",	--4977
		x"28",	--4978
		x"47",	--4979
		x"7e",	--4980
		x"3a",	--4981
		x"8c",	--4982
		x"7e",	--4983
		x"58",	--4984
		x"21",	--4985
		x"e9",	--4986
		x"7e",	--4987
		x"6f",	--4988
		x"24",	--4989
		x"7e",	--4990
		x"70",	--4991
		x"0a",	--4992
		x"7e",	--4993
		x"69",	--4994
		x"e3",	--4995
		x"7e",	--4996
		x"6c",	--4997
		x"22",	--4998
		x"7e",	--4999
		x"64",	--5000
		x"11",	--5001
		x"dc",	--5002
		x"7e",	--5003
		x"73",	--5004
		x"98",	--5005
		x"7e",	--5006
		x"74",	--5007
		x"04",	--5008
		x"7e",	--5009
		x"70",	--5010
		x"07",	--5011
		x"b8",	--5012
		x"7e",	--5013
		x"75",	--5014
		x"d1",	--5015
		x"7e",	--5016
		x"78",	--5017
		x"d2",	--5018
		x"19",	--5019
		x"3e",	--5020
		x"18",	--5021
		x"2c",	--5022
		x"08",	--5023
		x"30",	--5024
		x"4c",	--5025
		x"b1",	--5026
		x"28",	--5027
		x"cb",	--5028
		x"f1",	--5029
		x"00",	--5030
		x"30",	--5031
		x"7c",	--5032
		x"69",	--5033
		x"59",	--5034
		x"6e",	--5035
		x"04",	--5036
		x"7e",	--5037
		x"fe",	--5038
		x"6e",	--5039
		x"01",	--5040
		x"5e",	--5041
		x"c1",	--5042
		x"00",	--5043
		x"30",	--5044
		x"7c",	--5045
		x"f1",	--5046
		x"10",	--5047
		x"00",	--5048
		x"30",	--5049
		x"7c",	--5050
		x"f1",	--5051
		x"2b",	--5052
		x"02",	--5053
		x"30",	--5054
		x"7c",	--5055
		x"f1",	--5056
		x"2b",	--5057
		x"02",	--5058
		x"02",	--5059
		x"30",	--5060
		x"7c",	--5061
		x"f1",	--5062
		x"20",	--5063
		x"02",	--5064
		x"30",	--5065
		x"7c",	--5066
		x"c1",	--5067
		x"2a",	--5068
		x"02",	--5069
		x"30",	--5070
		x"62",	--5071
		x"d1",	--5072
		x"2e",	--5073
		x"30",	--5074
		x"7c",	--5075
		x"0e",	--5076
		x"2e",	--5077
		x"2a",	--5078
		x"0a",	--5079
		x"03",	--5080
		x"81",	--5081
		x"26",	--5082
		x"0d",	--5083
		x"c1",	--5084
		x"2e",	--5085
		x"02",	--5086
		x"30",	--5087
		x"72",	--5088
		x"f1",	--5089
		x"10",	--5090
		x"00",	--5091
		x"3a",	--5092
		x"81",	--5093
		x"26",	--5094
		x"91",	--5095
		x"26",	--5096
		x"05",	--5097
		x"27",	--5098
		x"81",	--5099
		x"26",	--5100
		x"15",	--5101
		x"c1",	--5102
		x"2e",	--5103
		x"12",	--5104
		x"69",	--5105
		x"79",	--5106
		x"10",	--5107
		x"5e",	--5108
		x"01",	--5109
		x"4e",	--5110
		x"4e",	--5111
		x"0e",	--5112
		x"0e",	--5113
		x"4e",	--5114
		x"6a",	--5115
		x"7a",	--5116
		x"7f",	--5117
		x"4a",	--5118
		x"c1",	--5119
		x"00",	--5120
		x"30",	--5121
		x"7c",	--5122
		x"1a",	--5123
		x"26",	--5124
		x"0a",	--5125
		x"0c",	--5126
		x"0c",	--5127
		x"0c",	--5128
		x"0a",	--5129
		x"81",	--5130
		x"26",	--5131
		x"b1",	--5132
		x"d0",	--5133
		x"26",	--5134
		x"8e",	--5135
		x"81",	--5136
		x"26",	--5137
		x"d1",	--5138
		x"2a",	--5139
		x"30",	--5140
		x"7c",	--5141
		x"07",	--5142
		x"27",	--5143
		x"6e",	--5144
		x"c1",	--5145
		x"2e",	--5146
		x"03",	--5147
		x"c1",	--5148
		x"2a",	--5149
		x"26",	--5150
		x"c1",	--5151
		x"04",	--5152
		x"c1",	--5153
		x"05",	--5154
		x"0e",	--5155
		x"2e",	--5156
		x"03",	--5157
		x"07",	--5158
		x"27",	--5159
		x"2e",	--5160
		x"c1",	--5161
		x"2e",	--5162
		x"07",	--5163
		x"e1",	--5164
		x"01",	--5165
		x"1f",	--5166
		x"26",	--5167
		x"c1",	--5168
		x"03",	--5169
		x"06",	--5170
		x"c1",	--5171
		x"2a",	--5172
		x"03",	--5173
		x"91",	--5174
		x"26",	--5175
		x"30",	--5176
		x"0e",	--5177
		x"02",	--5178
		x"3e",	--5179
		x"98",	--5180
		x"11",	--5181
		x"04",	--5182
		x"11",	--5183
		x"04",	--5184
		x"1d",	--5185
		x"34",	--5186
		x"1f",	--5187
		x"3e",	--5188
		x"b0",	--5189
		x"70",	--5190
		x"21",	--5191
		x"81",	--5192
		x"2c",	--5193
		x"05",	--5194
		x"30",	--5195
		x"5e",	--5196
		x"07",	--5197
		x"27",	--5198
		x"29",	--5199
		x"81",	--5200
		x"1e",	--5201
		x"5e",	--5202
		x"09",	--5203
		x"01",	--5204
		x"4e",	--5205
		x"4e",	--5206
		x"4e",	--5207
		x"4e",	--5208
		x"6a",	--5209
		x"7a",	--5210
		x"f7",	--5211
		x"4a",	--5212
		x"c1",	--5213
		x"00",	--5214
		x"05",	--5215
		x"b1",	--5216
		x"10",	--5217
		x"28",	--5218
		x"53",	--5219
		x"d1",	--5220
		x"01",	--5221
		x"06",	--5222
		x"e1",	--5223
		x"00",	--5224
		x"b1",	--5225
		x"0a",	--5226
		x"28",	--5227
		x"03",	--5228
		x"b1",	--5229
		x"10",	--5230
		x"28",	--5231
		x"6b",	--5232
		x"6b",	--5233
		x"24",	--5234
		x"0c",	--5235
		x"3c",	--5236
		x"28",	--5237
		x"17",	--5238
		x"02",	--5239
		x"16",	--5240
		x"04",	--5241
		x"1b",	--5242
		x"06",	--5243
		x"81",	--5244
		x"1e",	--5245
		x"81",	--5246
		x"20",	--5247
		x"81",	--5248
		x"22",	--5249
		x"81",	--5250
		x"24",	--5251
		x"d1",	--5252
		x"2b",	--5253
		x"08",	--5254
		x"06",	--5255
		x"07",	--5256
		x"04",	--5257
		x"06",	--5258
		x"02",	--5259
		x"0b",	--5260
		x"02",	--5261
		x"c1",	--5262
		x"2b",	--5263
		x"0b",	--5264
		x"0b",	--5265
		x"0b",	--5266
		x"c1",	--5267
		x"2f",	--5268
		x"05",	--5269
		x"20",	--5270
		x"5b",	--5271
		x"07",	--5272
		x"0d",	--5273
		x"27",	--5274
		x"28",	--5275
		x"1b",	--5276
		x"02",	--5277
		x"81",	--5278
		x"1e",	--5279
		x"81",	--5280
		x"20",	--5281
		x"d1",	--5282
		x"2b",	--5283
		x"08",	--5284
		x"09",	--5285
		x"06",	--5286
		x"27",	--5287
		x"2b",	--5288
		x"81",	--5289
		x"1e",	--5290
		x"d1",	--5291
		x"2b",	--5292
		x"0b",	--5293
		x"02",	--5294
		x"c1",	--5295
		x"2b",	--5296
		x"0b",	--5297
		x"0b",	--5298
		x"0b",	--5299
		x"c1",	--5300
		x"2f",	--5301
		x"05",	--5302
		x"f1",	--5303
		x"00",	--5304
		x"12",	--5305
		x"c1",	--5306
		x"2b",	--5307
		x"0f",	--5308
		x"68",	--5309
		x"b1",	--5310
		x"10",	--5311
		x"28",	--5312
		x"03",	--5313
		x"78",	--5314
		x"40",	--5315
		x"05",	--5316
		x"b1",	--5317
		x"28",	--5318
		x"04",	--5319
		x"78",	--5320
		x"20",	--5321
		x"c1",	--5322
		x"00",	--5323
		x"68",	--5324
		x"68",	--5325
		x"30",	--5326
		x"c1",	--5327
		x"2f",	--5328
		x"2d",	--5329
		x"f1",	--5330
		x"2d",	--5331
		x"02",	--5332
		x"68",	--5333
		x"11",	--5334
		x"b1",	--5335
		x"1e",	--5336
		x"b1",	--5337
		x"20",	--5338
		x"b1",	--5339
		x"22",	--5340
		x"b1",	--5341
		x"24",	--5342
		x"91",	--5343
		x"1e",	--5344
		x"81",	--5345
		x"20",	--5346
		x"81",	--5347
		x"22",	--5348
		x"81",	--5349
		x"24",	--5350
		x"17",	--5351
		x"58",	--5352
		x"0f",	--5353
		x"1a",	--5354
		x"1e",	--5355
		x"1b",	--5356
		x"20",	--5357
		x"3a",	--5358
		x"3b",	--5359
		x"0e",	--5360
		x"0f",	--5361
		x"1e",	--5362
		x"0f",	--5363
		x"81",	--5364
		x"1e",	--5365
		x"81",	--5366
		x"20",	--5367
		x"06",	--5368
		x"1a",	--5369
		x"1e",	--5370
		x"3a",	--5371
		x"1a",	--5372
		x"81",	--5373
		x"1e",	--5374
		x"c1",	--5375
		x"1b",	--5376
		x"68",	--5377
		x"6a",	--5378
		x"16",	--5379
		x"1e",	--5380
		x"91",	--5381
		x"20",	--5382
		x"3c",	--5383
		x"18",	--5384
		x"22",	--5385
		x"14",	--5386
		x"24",	--5387
		x"07",	--5388
		x"37",	--5389
		x"1a",	--5390
		x"09",	--5391
		x"91",	--5392
		x"28",	--5393
		x"32",	--5394
		x"1b",	--5395
		x"28",	--5396
		x"8b",	--5397
		x"8b",	--5398
		x"8b",	--5399
		x"8b",	--5400
		x"81",	--5401
		x"34",	--5402
		x"81",	--5403
		x"36",	--5404
		x"81",	--5405
		x"38",	--5406
		x"11",	--5407
		x"3a",	--5408
		x"11",	--5409
		x"3a",	--5410
		x"11",	--5411
		x"3a",	--5412
		x"11",	--5413
		x"3a",	--5414
		x"0c",	--5415
		x"1d",	--5416
		x"44",	--5417
		x"0e",	--5418
		x"0f",	--5419
		x"b0",	--5420
		x"12",	--5421
		x"31",	--5422
		x"0b",	--5423
		x"3c",	--5424
		x"0a",	--5425
		x"05",	--5426
		x"7b",	--5427
		x"30",	--5428
		x"c7",	--5429
		x"00",	--5430
		x"0c",	--5431
		x"4b",	--5432
		x"d1",	--5433
		x"01",	--5434
		x"03",	--5435
		x"7a",	--5436
		x"37",	--5437
		x"02",	--5438
		x"7a",	--5439
		x"57",	--5440
		x"4a",	--5441
		x"c7",	--5442
		x"00",	--5443
		x"06",	--5444
		x"36",	--5445
		x"11",	--5446
		x"3a",	--5447
		x"11",	--5448
		x"3a",	--5449
		x"11",	--5450
		x"3a",	--5451
		x"11",	--5452
		x"3a",	--5453
		x"0c",	--5454
		x"1d",	--5455
		x"44",	--5456
		x"0e",	--5457
		x"0f",	--5458
		x"b0",	--5459
		x"ec",	--5460
		x"31",	--5461
		x"09",	--5462
		x"81",	--5463
		x"3c",	--5464
		x"08",	--5465
		x"04",	--5466
		x"37",	--5467
		x"0c",	--5468
		x"b2",	--5469
		x"0d",	--5470
		x"b0",	--5471
		x"0e",	--5472
		x"ae",	--5473
		x"0f",	--5474
		x"ac",	--5475
		x"81",	--5476
		x"1e",	--5477
		x"81",	--5478
		x"20",	--5479
		x"81",	--5480
		x"22",	--5481
		x"81",	--5482
		x"24",	--5483
		x"6c",	--5484
		x"58",	--5485
		x"3e",	--5486
		x"14",	--5487
		x"1e",	--5488
		x"17",	--5489
		x"20",	--5490
		x"08",	--5491
		x"38",	--5492
		x"1a",	--5493
		x"19",	--5494
		x"28",	--5495
		x"89",	--5496
		x"89",	--5497
		x"89",	--5498
		x"89",	--5499
		x"1c",	--5500
		x"28",	--5501
		x"0d",	--5502
		x"0e",	--5503
		x"0f",	--5504
		x"b0",	--5505
		x"16",	--5506
		x"0b",	--5507
		x"3e",	--5508
		x"0a",	--5509
		x"05",	--5510
		x"7b",	--5511
		x"30",	--5512
		x"c8",	--5513
		x"00",	--5514
		x"0c",	--5515
		x"4b",	--5516
		x"d1",	--5517
		x"01",	--5518
		x"03",	--5519
		x"7a",	--5520
		x"37",	--5521
		x"02",	--5522
		x"7a",	--5523
		x"57",	--5524
		x"4a",	--5525
		x"c8",	--5526
		x"00",	--5527
		x"06",	--5528
		x"36",	--5529
		x"1c",	--5530
		x"28",	--5531
		x"0d",	--5532
		x"0e",	--5533
		x"0f",	--5534
		x"b0",	--5535
		x"e0",	--5536
		x"04",	--5537
		x"07",	--5538
		x"38",	--5539
		x"0e",	--5540
		x"d0",	--5541
		x"0f",	--5542
		x"ce",	--5543
		x"81",	--5544
		x"1e",	--5545
		x"81",	--5546
		x"20",	--5547
		x"2c",	--5548
		x"17",	--5549
		x"1e",	--5550
		x"08",	--5551
		x"38",	--5552
		x"1a",	--5553
		x"1e",	--5554
		x"28",	--5555
		x"0f",	--5556
		x"b0",	--5557
		x"86",	--5558
		x"0d",	--5559
		x"3f",	--5560
		x"0a",	--5561
		x"05",	--5562
		x"7d",	--5563
		x"30",	--5564
		x"c8",	--5565
		x"00",	--5566
		x"0c",	--5567
		x"4d",	--5568
		x"d1",	--5569
		x"01",	--5570
		x"03",	--5571
		x"7c",	--5572
		x"37",	--5573
		x"02",	--5574
		x"7c",	--5575
		x"57",	--5576
		x"4c",	--5577
		x"c8",	--5578
		x"00",	--5579
		x"06",	--5580
		x"36",	--5581
		x"1e",	--5582
		x"28",	--5583
		x"0f",	--5584
		x"b0",	--5585
		x"6c",	--5586
		x"07",	--5587
		x"38",	--5588
		x"0f",	--5589
		x"db",	--5590
		x"81",	--5591
		x"1e",	--5592
		x"b1",	--5593
		x"0a",	--5594
		x"28",	--5595
		x"02",	--5596
		x"c1",	--5597
		x"02",	--5598
		x"c1",	--5599
		x"2e",	--5600
		x"2a",	--5601
		x"0f",	--5602
		x"3f",	--5603
		x"1c",	--5604
		x"81",	--5605
		x"42",	--5606
		x"1a",	--5607
		x"1c",	--5608
		x"8a",	--5609
		x"8a",	--5610
		x"8a",	--5611
		x"8a",	--5612
		x"81",	--5613
		x"44",	--5614
		x"81",	--5615
		x"46",	--5616
		x"0a",	--5617
		x"8a",	--5618
		x"8a",	--5619
		x"8a",	--5620
		x"8a",	--5621
		x"81",	--5622
		x"48",	--5623
		x"1c",	--5624
		x"42",	--5625
		x"1d",	--5626
		x"44",	--5627
		x"1c",	--5628
		x"46",	--5629
		x"1d",	--5630
		x"48",	--5631
		x"2c",	--5632
		x"1c",	--5633
		x"26",	--5634
		x"0e",	--5635
		x"e1",	--5636
		x"01",	--5637
		x"5e",	--5638
		x"26",	--5639
		x"4e",	--5640
		x"c1",	--5641
		x"03",	--5642
		x"06",	--5643
		x"c1",	--5644
		x"2a",	--5645
		x"03",	--5646
		x"91",	--5647
		x"26",	--5648
		x"30",	--5649
		x"11",	--5650
		x"04",	--5651
		x"11",	--5652
		x"04",	--5653
		x"1d",	--5654
		x"34",	--5655
		x"0e",	--5656
		x"1e",	--5657
		x"1f",	--5658
		x"3e",	--5659
		x"b0",	--5660
		x"70",	--5661
		x"21",	--5662
		x"81",	--5663
		x"2c",	--5664
		x"0d",	--5665
		x"7f",	--5666
		x"8f",	--5667
		x"91",	--5668
		x"3c",	--5669
		x"0e",	--5670
		x"0e",	--5671
		x"19",	--5672
		x"40",	--5673
		x"f7",	--5674
		x"81",	--5675
		x"3e",	--5676
		x"81",	--5677
		x"2c",	--5678
		x"07",	--5679
		x"0e",	--5680
		x"91",	--5681
		x"26",	--5682
		x"30",	--5683
		x"d1",	--5684
		x"2e",	--5685
		x"c1",	--5686
		x"2a",	--5687
		x"03",	--5688
		x"05",	--5689
		x"d1",	--5690
		x"2a",	--5691
		x"81",	--5692
		x"26",	--5693
		x"17",	--5694
		x"16",	--5695
		x"40",	--5696
		x"6e",	--5697
		x"4e",	--5698
		x"02",	--5699
		x"30",	--5700
		x"54",	--5701
		x"1f",	--5702
		x"2c",	--5703
		x"31",	--5704
		x"4a",	--5705
		x"34",	--5706
		x"35",	--5707
		x"36",	--5708
		x"37",	--5709
		x"38",	--5710
		x"39",	--5711
		x"3a",	--5712
		x"3b",	--5713
		x"30",	--5714
		x"0d",	--5715
		x"0f",	--5716
		x"04",	--5717
		x"3d",	--5718
		x"03",	--5719
		x"3f",	--5720
		x"1f",	--5721
		x"0e",	--5722
		x"03",	--5723
		x"5d",	--5724
		x"3e",	--5725
		x"1e",	--5726
		x"0d",	--5727
		x"b0",	--5728
		x"6c",	--5729
		x"3d",	--5730
		x"6d",	--5731
		x"02",	--5732
		x"3e",	--5733
		x"1e",	--5734
		x"5d",	--5735
		x"02",	--5736
		x"3f",	--5737
		x"1f",	--5738
		x"30",	--5739
		x"b0",	--5740
		x"a6",	--5741
		x"0f",	--5742
		x"30",	--5743
		x"0b",	--5744
		x"0a",	--5745
		x"09",	--5746
		x"79",	--5747
		x"20",	--5748
		x"0a",	--5749
		x"0b",	--5750
		x"0c",	--5751
		x"0d",	--5752
		x"0e",	--5753
		x"0f",	--5754
		x"0c",	--5755
		x"0d",	--5756
		x"0d",	--5757
		x"06",	--5758
		x"02",	--5759
		x"0c",	--5760
		x"03",	--5761
		x"0c",	--5762
		x"0d",	--5763
		x"1e",	--5764
		x"19",	--5765
		x"f2",	--5766
		x"39",	--5767
		x"3a",	--5768
		x"3b",	--5769
		x"30",	--5770
		x"b0",	--5771
		x"e0",	--5772
		x"0e",	--5773
		x"0f",	--5774
		x"30",	--5775
		x"0b",	--5776
		x"0b",	--5777
		x"0f",	--5778
		x"06",	--5779
		x"3b",	--5780
		x"03",	--5781
		x"3e",	--5782
		x"3f",	--5783
		x"1e",	--5784
		x"0f",	--5785
		x"0d",	--5786
		x"05",	--5787
		x"5b",	--5788
		x"3c",	--5789
		x"3d",	--5790
		x"1c",	--5791
		x"0d",	--5792
		x"b0",	--5793
		x"e0",	--5794
		x"6b",	--5795
		x"04",	--5796
		x"3c",	--5797
		x"3d",	--5798
		x"1c",	--5799
		x"0d",	--5800
		x"5b",	--5801
		x"04",	--5802
		x"3e",	--5803
		x"3f",	--5804
		x"1e",	--5805
		x"0f",	--5806
		x"3b",	--5807
		x"30",	--5808
		x"b0",	--5809
		x"20",	--5810
		x"0e",	--5811
		x"0f",	--5812
		x"30",	--5813
		x"7c",	--5814
		x"10",	--5815
		x"0d",	--5816
		x"0e",	--5817
		x"0f",	--5818
		x"0e",	--5819
		x"0e",	--5820
		x"02",	--5821
		x"0e",	--5822
		x"1f",	--5823
		x"1c",	--5824
		x"f8",	--5825
		x"30",	--5826
		x"b0",	--5827
		x"6c",	--5828
		x"0f",	--5829
		x"30",	--5830
		x"07",	--5831
		x"06",	--5832
		x"05",	--5833
		x"04",	--5834
		x"30",	--5835
		x"40",	--5836
		x"04",	--5837
		x"05",	--5838
		x"06",	--5839
		x"07",	--5840
		x"08",	--5841
		x"09",	--5842
		x"0a",	--5843
		x"0b",	--5844
		x"0c",	--5845
		x"0d",	--5846
		x"0e",	--5847
		x"0f",	--5848
		x"08",	--5849
		x"09",	--5850
		x"0a",	--5851
		x"0b",	--5852
		x"0b",	--5853
		x"0e",	--5854
		x"08",	--5855
		x"0a",	--5856
		x"0b",	--5857
		x"05",	--5858
		x"09",	--5859
		x"08",	--5860
		x"02",	--5861
		x"08",	--5862
		x"05",	--5863
		x"08",	--5864
		x"09",	--5865
		x"0a",	--5866
		x"0b",	--5867
		x"1c",	--5868
		x"91",	--5869
		x"00",	--5870
		x"e5",	--5871
		x"21",	--5872
		x"34",	--5873
		x"35",	--5874
		x"36",	--5875
		x"37",	--5876
		x"30",	--5877
		x"0b",	--5878
		x"0a",	--5879
		x"09",	--5880
		x"08",	--5881
		x"18",	--5882
		x"0a",	--5883
		x"19",	--5884
		x"0c",	--5885
		x"1a",	--5886
		x"0e",	--5887
		x"1b",	--5888
		x"10",	--5889
		x"b0",	--5890
		x"8e",	--5891
		x"38",	--5892
		x"39",	--5893
		x"3a",	--5894
		x"3b",	--5895
		x"30",	--5896
		x"0b",	--5897
		x"0a",	--5898
		x"09",	--5899
		x"08",	--5900
		x"18",	--5901
		x"0a",	--5902
		x"19",	--5903
		x"0c",	--5904
		x"1a",	--5905
		x"0e",	--5906
		x"1b",	--5907
		x"10",	--5908
		x"b0",	--5909
		x"8e",	--5910
		x"0c",	--5911
		x"0d",	--5912
		x"0e",	--5913
		x"0f",	--5914
		x"38",	--5915
		x"39",	--5916
		x"3a",	--5917
		x"3b",	--5918
		x"30",	--5919
		x"0b",	--5920
		x"0a",	--5921
		x"09",	--5922
		x"08",	--5923
		x"07",	--5924
		x"18",	--5925
		x"0c",	--5926
		x"19",	--5927
		x"0e",	--5928
		x"1a",	--5929
		x"10",	--5930
		x"1b",	--5931
		x"12",	--5932
		x"b0",	--5933
		x"8e",	--5934
		x"17",	--5935
		x"14",	--5936
		x"87",	--5937
		x"00",	--5938
		x"87",	--5939
		x"02",	--5940
		x"87",	--5941
		x"04",	--5942
		x"87",	--5943
		x"06",	--5944
		x"37",	--5945
		x"38",	--5946
		x"39",	--5947
		x"3a",	--5948
		x"3b",	--5949
		x"30",	--5950
		x"00",	--5951
		x"32",	--5952
		x"f0",	--5953
		x"fd",	--5954
		x"25",	--5955
		x"20",	--5956
		x"0d",	--5957
		x"00",	--5958
		x"74",	--5959
		x"70",	--5960
		x"0a",	--5961
		x"63",	--5962
		x"72",	--5963
		x"65",	--5964
		x"74",	--5965
		x"75",	--5966
		x"61",	--5967
		x"65",	--5968
		x"0d",	--5969
		x"00",	--5970
		x"25",	--5971
		x"20",	--5972
		x"45",	--5973
		x"54",	--5974
		x"52",	--5975
		x"47",	--5976
		x"54",	--5977
		x"3c",	--5978
		x"49",	--5979
		x"45",	--5980
		x"55",	--5981
		x"3e",	--5982
		x"0a",	--5983
		x"25",	--5984
		x"20",	--5985
		x"64",	--5986
		x"0a",	--5987
		x"4e",	--5988
		x"74",	--5989
		x"69",	--5990
		x"70",	--5991
		x"65",	--5992
		x"65",	--5993
		x"74",	--5994
		x"64",	--5995
		x"59",	--5996
		x"74",	--5997
		x"0a",	--5998
		x"57",	--5999
		x"69",	--6000
		x"69",	--6001
		x"67",	--6002
		x"66",	--6003
		x"72",	--6004
		x"61",	--6005
		x"6e",	--6006
		x"77",	--6007
		x"2e",	--6008
		x"69",	--6009
		x"20",	--6010
		x"69",	--6011
		x"65",	--6012
		x"0a",	--6013
		x"57",	--6014
		x"20",	--6015
		x"68",	--6016
		x"75",	--6017
		x"64",	--6018
		x"6e",	--6019
		x"74",	--6020
		x"73",	--6021
		x"65",	--6022
		x"74",	--6023
		x"61",	--6024
		x"0d",	--6025
		x"00",	--6026
		x"74",	--6027
		x"70",	--6028
		x"0a",	--6029
		x"65",	--6030
		x"72",	--6031
		x"72",	--6032
		x"20",	--6033
		x"69",	--6034
		x"73",	--6035
		x"6e",	--6036
		x"20",	--6037
		x"72",	--6038
		x"75",	--6039
		x"65",	--6040
		x"74",	--6041
		x"0a",	--6042
		x"63",	--6043
		x"72",	--6044
		x"65",	--6045
		x"74",	--6046
		x"75",	--6047
		x"61",	--6048
		x"65",	--6049
		x"0d",	--6050
		x"00",	--6051
		x"25",	--6052
		x"20",	--6053
		x"45",	--6054
		x"54",	--6055
		x"52",	--6056
		x"47",	--6057
		x"54",	--6058
		x"3c",	--6059
		x"49",	--6060
		x"45",	--6061
		x"55",	--6062
		x"3e",	--6063
		x"0a",	--6064
		x"25",	--6065
		x"20",	--6066
		x"64",	--6067
		x"0a",	--6068
		x"25",	--6069
		x"64",	--6070
		x"25",	--6071
		x"64",	--6072
		x"25",	--6073
		x"0d",	--6074
		x"00",	--6075
		x"64",	--6076
		x"25",	--6077
		x"0d",	--6078
		x"00",	--6079
		x"22",	--6080
		x"4a",	--6081
		x"50",	--6082
		x"58",	--6083
		x"60",	--6084
		x"68",	--6085
		x"3a",	--6086
		x"42",	--6087
		x"0d",	--6088
		x"3d",	--6089
		x"3d",	--6090
		x"3d",	--6091
		x"20",	--6092
		x"61",	--6093
		x"63",	--6094
		x"6c",	--6095
		x"4d",	--6096
		x"55",	--6097
		x"3d",	--6098
		x"3d",	--6099
		x"3d",	--6100
		x"0d",	--6101
		x"00",	--6102
		x"6e",	--6103
		x"65",	--6104
		x"61",	--6105
		x"74",	--6106
		x"76",	--6107
		x"20",	--6108
		x"6f",	--6109
		x"65",	--6110
		x"77",	--6111
		x"69",	--6112
		x"65",	--6113
		x"72",	--6114
		x"61",	--6115
		x"00",	--6116
		x"75",	--6117
		x"7a",	--6118
		x"72",	--6119
		x"70",	--6120
		x"6d",	--6121
		x"65",	--6122
		x"63",	--6123
		x"64",	--6124
		x"72",	--6125
		x"73",	--6126
		x"65",	--6127
		x"64",	--6128
		x"63",	--6129
		x"6e",	--6130
		x"72",	--6131
		x"6c",	--6132
		x"65",	--6133
		x"00",	--6134
		x"70",	--6135
		x"65",	--6136
		x"20",	--6137
		x"6f",	--6138
		x"66",	--6139
		x"67",	--6140
		x"72",	--6141
		x"74",	--6142
		x"6f",	--6143
		x"00",	--6144
		x"72",	--6145
		x"30",	--6146
		x"00",	--6147
		x"6f",	--6148
		x"74",	--6149
		x"6f",	--6150
		x"64",	--6151
		x"72",	--6152
		x"0d",	--6153
		x"00",	--6154
		x"20",	--6155
		x"00",	--6156
		x"63",	--6157
		x"55",	--6158
		x"0d",	--6159
		x"00",	--6160
		x"4f",	--6161
		x"4e",	--6162
		x"0a",	--6163
		x"52",	--6164
		x"47",	--6165
		x"54",	--6166
		x"0a",	--6167
		x"4c",	--6168
		x"46",	--6169
		x"0d",	--6170
		x"00",	--6171
		x"77",	--6172
		x"69",	--6173
		x"65",	--6174
		x"0d",	--6175
		x"65",	--6176
		x"72",	--6177
		x"72",	--6178
		x"20",	--6179
		x"69",	--6180
		x"73",	--6181
		x"6e",	--6182
		x"20",	--6183
		x"72",	--6184
		x"75",	--6185
		x"65",	--6186
		x"74",	--6187
		x"0a",	--6188
		x"63",	--6189
		x"72",	--6190
		x"65",	--6191
		x"74",	--6192
		x"75",	--6193
		x"61",	--6194
		x"65",	--6195
		x"0d",	--6196
		x"00",	--6197
		x"25",	--6198
		x"20",	--6199
		x"45",	--6200
		x"49",	--6201
		x"54",	--6202
		x"52",	--6203
		x"56",	--6204
		x"4c",	--6205
		x"45",	--6206
		x"0a",	--6207
		x"72",	--6208
		x"25",	--6209
		x"20",	--6210
		x"3d",	--6211
		x"64",	--6212
		x"0a",	--6213
		x"09",	--6214
		x"73",	--6215
		x"52",	--6216
		x"47",	--6217
		x"53",	--6218
		x"45",	--6219
		x"0d",	--6220
		x"00",	--6221
		x"65",	--6222
		x"64",	--6223
		x"0d",	--6224
		x"25",	--6225
		x"20",	--6226
		x"73",	--6227
		x"6e",	--6228
		x"74",	--6229
		x"61",	--6230
		x"6e",	--6231
		x"6d",	--6232
		x"65",	--6233
		x"0d",	--6234
		x"00",	--6235
		x"63",	--6236
		x"25",	--6237
		x"0d",	--6238
		x"00",	--6239
		x"63",	--6240
		x"20",	--6241
		x"6f",	--6242
		x"73",	--6243
		x"63",	--6244
		x"20",	--6245
		x"6f",	--6246
		x"6d",	--6247
		x"6e",	--6248
		x"0d",	--6249
		x"00",	--6250
		x"ee",	--6251
		x"1c",	--6252
		x"1c",	--6253
		x"1c",	--6254
		x"1c",	--6255
		x"1c",	--6256
		x"1c",	--6257
		x"1c",	--6258
		x"1c",	--6259
		x"1c",	--6260
		x"1c",	--6261
		x"1c",	--6262
		x"1c",	--6263
		x"1c",	--6264
		x"1c",	--6265
		x"1c",	--6266
		x"1c",	--6267
		x"1c",	--6268
		x"1c",	--6269
		x"1c",	--6270
		x"1c",	--6271
		x"1c",	--6272
		x"1c",	--6273
		x"1c",	--6274
		x"1c",	--6275
		x"1c",	--6276
		x"1c",	--6277
		x"1c",	--6278
		x"1c",	--6279
		x"e0",	--6280
		x"1c",	--6281
		x"1c",	--6282
		x"1c",	--6283
		x"1c",	--6284
		x"1c",	--6285
		x"1c",	--6286
		x"1c",	--6287
		x"1c",	--6288
		x"1c",	--6289
		x"1c",	--6290
		x"1c",	--6291
		x"1c",	--6292
		x"1c",	--6293
		x"1c",	--6294
		x"1c",	--6295
		x"1c",	--6296
		x"1c",	--6297
		x"1c",	--6298
		x"1c",	--6299
		x"1c",	--6300
		x"1c",	--6301
		x"1c",	--6302
		x"1c",	--6303
		x"1c",	--6304
		x"1c",	--6305
		x"1c",	--6306
		x"1c",	--6307
		x"1c",	--6308
		x"1c",	--6309
		x"1c",	--6310
		x"1c",	--6311
		x"d2",	--6312
		x"c4",	--6313
		x"b6",	--6314
		x"1c",	--6315
		x"1c",	--6316
		x"1c",	--6317
		x"1c",	--6318
		x"1c",	--6319
		x"1c",	--6320
		x"1c",	--6321
		x"9e",	--6322
		x"1c",	--6323
		x"8c",	--6324
		x"1c",	--6325
		x"1c",	--6326
		x"1c",	--6327
		x"1c",	--6328
		x"70",	--6329
		x"1c",	--6330
		x"1c",	--6331
		x"1c",	--6332
		x"62",	--6333
		x"50",	--6334
		x"30",	--6335
		x"32",	--6336
		x"34",	--6337
		x"36",	--6338
		x"38",	--6339
		x"61",	--6340
		x"63",	--6341
		x"65",	--6342
		x"00",	--6343
		x"00",	--6344
		x"00",	--6345
		x"00",	--6346
		x"00",	--6347
		x"00",	--6348
		x"02",	--6349
		x"03",	--6350
		x"03",	--6351
		x"04",	--6352
		x"04",	--6353
		x"04",	--6354
		x"04",	--6355
		x"05",	--6356
		x"05",	--6357
		x"05",	--6358
		x"05",	--6359
		x"05",	--6360
		x"05",	--6361
		x"05",	--6362
		x"05",	--6363
		x"06",	--6364
		x"06",	--6365
		x"06",	--6366
		x"06",	--6367
		x"06",	--6368
		x"06",	--6369
		x"06",	--6370
		x"06",	--6371
		x"06",	--6372
		x"06",	--6373
		x"06",	--6374
		x"06",	--6375
		x"06",	--6376
		x"06",	--6377
		x"06",	--6378
		x"06",	--6379
		x"07",	--6380
		x"07",	--6381
		x"07",	--6382
		x"07",	--6383
		x"07",	--6384
		x"07",	--6385
		x"07",	--6386
		x"07",	--6387
		x"07",	--6388
		x"07",	--6389
		x"07",	--6390
		x"07",	--6391
		x"07",	--6392
		x"07",	--6393
		x"07",	--6394
		x"07",	--6395
		x"07",	--6396
		x"07",	--6397
		x"07",	--6398
		x"07",	--6399
		x"07",	--6400
		x"07",	--6401
		x"07",	--6402
		x"07",	--6403
		x"07",	--6404
		x"07",	--6405
		x"07",	--6406
		x"07",	--6407
		x"07",	--6408
		x"07",	--6409
		x"07",	--6410
		x"07",	--6411
		x"08",	--6412
		x"08",	--6413
		x"08",	--6414
		x"08",	--6415
		x"08",	--6416
		x"08",	--6417
		x"08",	--6418
		x"08",	--6419
		x"08",	--6420
		x"08",	--6421
		x"08",	--6422
		x"08",	--6423
		x"08",	--6424
		x"08",	--6425
		x"08",	--6426
		x"08",	--6427
		x"08",	--6428
		x"08",	--6429
		x"08",	--6430
		x"08",	--6431
		x"08",	--6432
		x"08",	--6433
		x"08",	--6434
		x"08",	--6435
		x"08",	--6436
		x"08",	--6437
		x"08",	--6438
		x"08",	--6439
		x"08",	--6440
		x"08",	--6441
		x"08",	--6442
		x"08",	--6443
		x"08",	--6444
		x"08",	--6445
		x"08",	--6446
		x"08",	--6447
		x"08",	--6448
		x"08",	--6449
		x"08",	--6450
		x"08",	--6451
		x"08",	--6452
		x"08",	--6453
		x"08",	--6454
		x"08",	--6455
		x"08",	--6456
		x"08",	--6457
		x"08",	--6458
		x"08",	--6459
		x"08",	--6460
		x"08",	--6461
		x"08",	--6462
		x"08",	--6463
		x"08",	--6464
		x"08",	--6465
		x"08",	--6466
		x"08",	--6467
		x"08",	--6468
		x"08",	--6469
		x"08",	--6470
		x"08",	--6471
		x"08",	--6472
		x"08",	--6473
		x"08",	--6474
		x"08",	--6475
		x"28",	--6476
		x"75",	--6477
		x"6c",	--6478
		x"00",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"68",	--6484
		x"6c",	--6485
		x"00",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"6a",	--8176
		x"6a",	--8177
		x"6a",	--8178
		x"6a",	--8179
		x"6a",	--8180
		x"6a",	--8181
		x"6a",	--8182
		x"f8",	--8183
		x"4a",	--8184
		x"6a",	--8185
		x"6a",	--8186
		x"6a",	--8187
		x"6a",	--8188
		x"6a",	--8189
		x"6a",	--8190
		x"00");	--8191
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"05",	--5
		x"40",	--6
		x"0a",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"05",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"f2",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"03",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"05",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"d5",	--44
		x"12",	--45
		x"cf",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"ef",	--50
		x"12",	--51
		x"d4",	--52
		x"53",	--53
		x"40",	--54
		x"ef",	--55
		x"40",	--56
		x"c9",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"cf",	--61
		x"40",	--62
		x"ef",	--63
		x"40",	--64
		x"cc",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"cf",	--69
		x"40",	--70
		x"ef",	--71
		x"40",	--72
		x"cc",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"cf",	--77
		x"40",	--78
		x"ef",	--79
		x"40",	--80
		x"c4",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"cf",	--85
		x"40",	--86
		x"ef",	--87
		x"40",	--88
		x"c7",	--89
		x"40",	--90
		x"00",	--91
		x"12",	--92
		x"cf",	--93
		x"40",	--94
		x"ef",	--95
		x"40",	--96
		x"c8",	--97
		x"40",	--98
		x"00",	--99
		x"12",	--100
		x"cf",	--101
		x"40",	--102
		x"ef",	--103
		x"40",	--104
		x"c4",	--105
		x"40",	--106
		x"00",	--107
		x"12",	--108
		x"cf",	--109
		x"40",	--110
		x"ef",	--111
		x"40",	--112
		x"c5",	--113
		x"40",	--114
		x"00",	--115
		x"12",	--116
		x"cf",	--117
		x"40",	--118
		x"f0",	--119
		x"40",	--120
		x"c3",	--121
		x"40",	--122
		x"00",	--123
		x"12",	--124
		x"cf",	--125
		x"40",	--126
		x"f0",	--127
		x"40",	--128
		x"c5",	--129
		x"40",	--130
		x"00",	--131
		x"12",	--132
		x"cf",	--133
		x"43",	--134
		x"43",	--135
		x"12",	--136
		x"cf",	--137
		x"43",	--138
		x"40",	--139
		x"4e",	--140
		x"40",	--141
		x"01",	--142
		x"41",	--143
		x"50",	--144
		x"00",	--145
		x"12",	--146
		x"ce",	--147
		x"41",	--148
		x"50",	--149
		x"00",	--150
		x"12",	--151
		x"ce",	--152
		x"43",	--153
		x"40",	--154
		x"4e",	--155
		x"40",	--156
		x"01",	--157
		x"41",	--158
		x"52",	--159
		x"12",	--160
		x"ce",	--161
		x"41",	--162
		x"52",	--163
		x"12",	--164
		x"ce",	--165
		x"41",	--166
		x"52",	--167
		x"41",	--168
		x"50",	--169
		x"00",	--170
		x"12",	--171
		x"c7",	--172
		x"40",	--173
		x"01",	--174
		x"41",	--175
		x"50",	--176
		x"00",	--177
		x"12",	--178
		x"d1",	--179
		x"40",	--180
		x"01",	--181
		x"41",	--182
		x"52",	--183
		x"12",	--184
		x"d1",	--185
		x"41",	--186
		x"52",	--187
		x"41",	--188
		x"50",	--189
		x"00",	--190
		x"12",	--191
		x"c8",	--192
		x"41",	--193
		x"52",	--194
		x"41",	--195
		x"50",	--196
		x"00",	--197
		x"12",	--198
		x"c8",	--199
		x"12",	--200
		x"d0",	--201
		x"40",	--202
		x"01",	--203
		x"41",	--204
		x"53",	--205
		x"12",	--206
		x"d1",	--207
		x"41",	--208
		x"53",	--209
		x"12",	--210
		x"c4",	--211
		x"40",	--212
		x"00",	--213
		x"40",	--214
		x"11",	--215
		x"41",	--216
		x"53",	--217
		x"12",	--218
		x"d2",	--219
		x"40",	--220
		x"01",	--221
		x"41",	--222
		x"12",	--223
		x"d0",	--224
		x"41",	--225
		x"12",	--226
		x"c3",	--227
		x"12",	--228
		x"41",	--229
		x"12",	--230
		x"12",	--231
		x"12",	--232
		x"12",	--233
		x"39",	--234
		x"12",	--235
		x"b7",	--236
		x"12",	--237
		x"3a",	--238
		x"12",	--239
		x"49",	--240
		x"40",	--241
		x"00",	--242
		x"41",	--243
		x"50",	--244
		x"00",	--245
		x"41",	--246
		x"50",	--247
		x"00",	--248
		x"41",	--249
		x"50",	--250
		x"00",	--251
		x"12",	--252
		x"c6",	--253
		x"50",	--254
		x"00",	--255
		x"12",	--256
		x"41",	--257
		x"12",	--258
		x"12",	--259
		x"12",	--260
		x"12",	--261
		x"39",	--262
		x"12",	--263
		x"b7",	--264
		x"12",	--265
		x"3a",	--266
		x"12",	--267
		x"49",	--268
		x"40",	--269
		x"00",	--270
		x"41",	--271
		x"50",	--272
		x"00",	--273
		x"41",	--274
		x"50",	--275
		x"00",	--276
		x"41",	--277
		x"50",	--278
		x"00",	--279
		x"12",	--280
		x"c6",	--281
		x"50",	--282
		x"00",	--283
		x"41",	--284
		x"50",	--285
		x"00",	--286
		x"41",	--287
		x"50",	--288
		x"00",	--289
		x"12",	--290
		x"c4",	--291
		x"12",	--292
		x"c4",	--293
		x"40",	--294
		x"ff",	--295
		x"00",	--296
		x"d2",	--297
		x"43",	--298
		x"43",	--299
		x"3c",	--300
		x"43",	--301
		x"3c",	--302
		x"43",	--303
		x"3c",	--304
		x"43",	--305
		x"12",	--306
		x"d5",	--307
		x"93",	--308
		x"27",	--309
		x"12",	--310
		x"d5",	--311
		x"93",	--312
		x"20",	--313
		x"90",	--314
		x"00",	--315
		x"24",	--316
		x"90",	--317
		x"00",	--318
		x"27",	--319
		x"92",	--320
		x"20",	--321
		x"3c",	--322
		x"12",	--323
		x"f0",	--324
		x"12",	--325
		x"d4",	--326
		x"53",	--327
		x"40",	--328
		x"00",	--329
		x"51",	--330
		x"5f",	--331
		x"43",	--332
		x"00",	--333
		x"4f",	--334
		x"41",	--335
		x"00",	--336
		x"12",	--337
		x"cf",	--338
		x"43",	--339
		x"3f",	--340
		x"93",	--341
		x"27",	--342
		x"53",	--343
		x"12",	--344
		x"f0",	--345
		x"12",	--346
		x"d4",	--347
		x"53",	--348
		x"3f",	--349
		x"90",	--350
		x"00",	--351
		x"2f",	--352
		x"93",	--353
		x"02",	--354
		x"24",	--355
		x"4f",	--356
		x"11",	--357
		x"12",	--358
		x"12",	--359
		x"f0",	--360
		x"4f",	--361
		x"00",	--362
		x"12",	--363
		x"d4",	--364
		x"52",	--365
		x"41",	--366
		x"00",	--367
		x"40",	--368
		x"00",	--369
		x"51",	--370
		x"5a",	--371
		x"4f",	--372
		x"00",	--373
		x"53",	--374
		x"3f",	--375
		x"93",	--376
		x"20",	--377
		x"90",	--378
		x"00",	--379
		x"23",	--380
		x"3f",	--381
		x"93",	--382
		x"23",	--383
		x"90",	--384
		x"00",	--385
		x"24",	--386
		x"90",	--387
		x"00",	--388
		x"34",	--389
		x"90",	--390
		x"00",	--391
		x"23",	--392
		x"3c",	--393
		x"90",	--394
		x"00",	--395
		x"24",	--396
		x"90",	--397
		x"00",	--398
		x"23",	--399
		x"3c",	--400
		x"12",	--401
		x"f0",	--402
		x"12",	--403
		x"d4",	--404
		x"53",	--405
		x"12",	--406
		x"c5",	--407
		x"43",	--408
		x"3f",	--409
		x"12",	--410
		x"f0",	--411
		x"12",	--412
		x"d4",	--413
		x"53",	--414
		x"12",	--415
		x"c5",	--416
		x"43",	--417
		x"3f",	--418
		x"12",	--419
		x"f0",	--420
		x"12",	--421
		x"d4",	--422
		x"53",	--423
		x"12",	--424
		x"c5",	--425
		x"43",	--426
		x"3f",	--427
		x"12",	--428
		x"f0",	--429
		x"12",	--430
		x"d4",	--431
		x"53",	--432
		x"12",	--433
		x"c5",	--434
		x"43",	--435
		x"3f",	--436
		x"40",	--437
		x"ee",	--438
		x"12",	--439
		x"43",	--440
		x"4b",	--441
		x"42",	--442
		x"02",	--443
		x"12",	--444
		x"d0",	--445
		x"12",	--446
		x"12",	--447
		x"ee",	--448
		x"12",	--449
		x"d4",	--450
		x"52",	--451
		x"53",	--452
		x"90",	--453
		x"00",	--454
		x"23",	--455
		x"12",	--456
		x"ee",	--457
		x"12",	--458
		x"d4",	--459
		x"53",	--460
		x"41",	--461
		x"41",	--462
		x"4f",	--463
		x"02",	--464
		x"41",	--465
		x"12",	--466
		x"83",	--467
		x"4e",	--468
		x"43",	--469
		x"00",	--470
		x"93",	--471
		x"24",	--472
		x"93",	--473
		x"02",	--474
		x"24",	--475
		x"43",	--476
		x"02",	--477
		x"41",	--478
		x"4b",	--479
		x"00",	--480
		x"12",	--481
		x"cc",	--482
		x"43",	--483
		x"4f",	--484
		x"42",	--485
		x"02",	--486
		x"12",	--487
		x"d1",	--488
		x"43",	--489
		x"53",	--490
		x"41",	--491
		x"41",	--492
		x"93",	--493
		x"02",	--494
		x"24",	--495
		x"43",	--496
		x"02",	--497
		x"42",	--498
		x"02",	--499
		x"12",	--500
		x"d1",	--501
		x"43",	--502
		x"53",	--503
		x"41",	--504
		x"41",	--505
		x"43",	--506
		x"12",	--507
		x"c3",	--508
		x"43",	--509
		x"53",	--510
		x"41",	--511
		x"41",	--512
		x"43",	--513
		x"40",	--514
		x"c3",	--515
		x"12",	--516
		x"d0",	--517
		x"4f",	--518
		x"02",	--519
		x"3f",	--520
		x"4f",	--521
		x"02",	--522
		x"41",	--523
		x"12",	--524
		x"12",	--525
		x"82",	--526
		x"4f",	--527
		x"4e",	--528
		x"93",	--529
		x"38",	--530
		x"41",	--531
		x"4b",	--532
		x"00",	--533
		x"12",	--534
		x"cc",	--535
		x"4f",	--536
		x"93",	--537
		x"24",	--538
		x"41",	--539
		x"4b",	--540
		x"00",	--541
		x"4d",	--542
		x"00",	--543
		x"12",	--544
		x"cc",	--545
		x"4f",	--546
		x"41",	--547
		x"00",	--548
		x"42",	--549
		x"02",	--550
		x"12",	--551
		x"d2",	--552
		x"43",	--553
		x"52",	--554
		x"41",	--555
		x"41",	--556
		x"41",	--557
		x"40",	--558
		x"00",	--559
		x"40",	--560
		x"11",	--561
		x"3f",	--562
		x"40",	--563
		x"11",	--564
		x"3f",	--565
		x"43",	--566
		x"42",	--567
		x"02",	--568
		x"12",	--569
		x"c7",	--570
		x"43",	--571
		x"42",	--572
		x"02",	--573
		x"12",	--574
		x"c7",	--575
		x"12",	--576
		x"ee",	--577
		x"12",	--578
		x"d4",	--579
		x"53",	--580
		x"41",	--581
		x"93",	--582
		x"02",	--583
		x"24",	--584
		x"42",	--585
		x"02",	--586
		x"12",	--587
		x"c6",	--588
		x"42",	--589
		x"02",	--590
		x"12",	--591
		x"c6",	--592
		x"41",	--593
		x"43",	--594
		x"40",	--595
		x"c4",	--596
		x"12",	--597
		x"d0",	--598
		x"4f",	--599
		x"02",	--600
		x"3f",	--601
		x"4f",	--602
		x"02",	--603
		x"4e",	--604
		x"02",	--605
		x"41",	--606
		x"12",	--607
		x"12",	--608
		x"83",	--609
		x"4e",	--610
		x"90",	--611
		x"00",	--612
		x"38",	--613
		x"20",	--614
		x"41",	--615
		x"4b",	--616
		x"00",	--617
		x"12",	--618
		x"cd",	--619
		x"4f",	--620
		x"41",	--621
		x"4b",	--622
		x"00",	--623
		x"12",	--624
		x"cd",	--625
		x"4f",	--626
		x"12",	--627
		x"12",	--628
		x"12",	--629
		x"ee",	--630
		x"12",	--631
		x"d4",	--632
		x"50",	--633
		x"00",	--634
		x"4a",	--635
		x"42",	--636
		x"02",	--637
		x"12",	--638
		x"c7",	--639
		x"4b",	--640
		x"42",	--641
		x"02",	--642
		x"12",	--643
		x"c7",	--644
		x"43",	--645
		x"53",	--646
		x"41",	--647
		x"41",	--648
		x"41",	--649
		x"41",	--650
		x"4b",	--651
		x"00",	--652
		x"12",	--653
		x"cc",	--654
		x"43",	--655
		x"4f",	--656
		x"42",	--657
		x"02",	--658
		x"12",	--659
		x"d1",	--660
		x"3f",	--661
		x"12",	--662
		x"ee",	--663
		x"12",	--664
		x"d4",	--665
		x"4b",	--666
		x"00",	--667
		x"12",	--668
		x"ee",	--669
		x"12",	--670
		x"d4",	--671
		x"52",	--672
		x"43",	--673
		x"3f",	--674
		x"40",	--675
		x"ff",	--676
		x"42",	--677
		x"02",	--678
		x"12",	--679
		x"c7",	--680
		x"40",	--681
		x"00",	--682
		x"42",	--683
		x"02",	--684
		x"12",	--685
		x"c7",	--686
		x"43",	--687
		x"40",	--688
		x"00",	--689
		x"42",	--690
		x"02",	--691
		x"12",	--692
		x"d1",	--693
		x"41",	--694
		x"40",	--695
		x"00",	--696
		x"42",	--697
		x"02",	--698
		x"12",	--699
		x"c7",	--700
		x"40",	--701
		x"ff",	--702
		x"42",	--703
		x"02",	--704
		x"12",	--705
		x"c7",	--706
		x"43",	--707
		x"40",	--708
		x"00",	--709
		x"42",	--710
		x"02",	--711
		x"12",	--712
		x"d1",	--713
		x"41",	--714
		x"40",	--715
		x"ff",	--716
		x"42",	--717
		x"02",	--718
		x"12",	--719
		x"c7",	--720
		x"40",	--721
		x"ff",	--722
		x"42",	--723
		x"02",	--724
		x"12",	--725
		x"c7",	--726
		x"43",	--727
		x"40",	--728
		x"00",	--729
		x"42",	--730
		x"02",	--731
		x"12",	--732
		x"d1",	--733
		x"41",	--734
		x"40",	--735
		x"00",	--736
		x"42",	--737
		x"02",	--738
		x"12",	--739
		x"c7",	--740
		x"40",	--741
		x"00",	--742
		x"42",	--743
		x"02",	--744
		x"12",	--745
		x"c7",	--746
		x"43",	--747
		x"40",	--748
		x"00",	--749
		x"42",	--750
		x"02",	--751
		x"12",	--752
		x"d1",	--753
		x"41",	--754
		x"12",	--755
		x"ee",	--756
		x"12",	--757
		x"d4",	--758
		x"53",	--759
		x"43",	--760
		x"41",	--761
		x"40",	--762
		x"c0",	--763
		x"01",	--764
		x"40",	--765
		x"00",	--766
		x"01",	--767
		x"40",	--768
		x"02",	--769
		x"01",	--770
		x"12",	--771
		x"ee",	--772
		x"12",	--773
		x"d4",	--774
		x"43",	--775
		x"01",	--776
		x"40",	--777
		x"ee",	--778
		x"00",	--779
		x"12",	--780
		x"d4",	--781
		x"53",	--782
		x"43",	--783
		x"41",	--784
		x"12",	--785
		x"12",	--786
		x"12",	--787
		x"4f",	--788
		x"4f",	--789
		x"00",	--790
		x"12",	--791
		x"d1",	--792
		x"4e",	--793
		x"4f",	--794
		x"89",	--795
		x"00",	--796
		x"79",	--797
		x"00",	--798
		x"12",	--799
		x"dd",	--800
		x"4a",	--801
		x"00",	--802
		x"4b",	--803
		x"00",	--804
		x"4e",	--805
		x"4f",	--806
		x"49",	--807
		x"12",	--808
		x"cb",	--809
		x"43",	--810
		x"40",	--811
		x"3f",	--812
		x"12",	--813
		x"d8",	--814
		x"4e",	--815
		x"4f",	--816
		x"40",	--817
		x"66",	--818
		x"40",	--819
		x"3f",	--820
		x"12",	--821
		x"dc",	--822
		x"93",	--823
		x"24",	--824
		x"34",	--825
		x"40",	--826
		x"cc",	--827
		x"40",	--828
		x"3d",	--829
		x"4a",	--830
		x"4b",	--831
		x"12",	--832
		x"dd",	--833
		x"93",	--834
		x"34",	--835
		x"40",	--836
		x"cc",	--837
		x"40",	--838
		x"3d",	--839
		x"4a",	--840
		x"4b",	--841
		x"49",	--842
		x"00",	--843
		x"12",	--844
		x"ce",	--845
		x"41",	--846
		x"41",	--847
		x"41",	--848
		x"41",	--849
		x"40",	--850
		x"66",	--851
		x"40",	--852
		x"3f",	--853
		x"3f",	--854
		x"12",	--855
		x"12",	--856
		x"4f",	--857
		x"4c",	--858
		x"4e",	--859
		x"00",	--860
		x"4d",	--861
		x"00",	--862
		x"12",	--863
		x"00",	--864
		x"12",	--865
		x"00",	--866
		x"12",	--867
		x"00",	--868
		x"12",	--869
		x"00",	--870
		x"12",	--871
		x"00",	--872
		x"12",	--873
		x"00",	--874
		x"41",	--875
		x"00",	--876
		x"41",	--877
		x"00",	--878
		x"12",	--879
		x"ca",	--880
		x"50",	--881
		x"00",	--882
		x"4a",	--883
		x"00",	--884
		x"4b",	--885
		x"40",	--886
		x"c6",	--887
		x"12",	--888
		x"d0",	--889
		x"4f",	--890
		x"00",	--891
		x"41",	--892
		x"41",	--893
		x"41",	--894
		x"12",	--895
		x"4f",	--896
		x"4f",	--897
		x"00",	--898
		x"12",	--899
		x"d1",	--900
		x"4e",	--901
		x"00",	--902
		x"4f",	--903
		x"00",	--904
		x"43",	--905
		x"4b",	--906
		x"00",	--907
		x"4b",	--908
		x"00",	--909
		x"12",	--910
		x"d1",	--911
		x"41",	--912
		x"41",	--913
		x"12",	--914
		x"4f",	--915
		x"43",	--916
		x"40",	--917
		x"3f",	--918
		x"4f",	--919
		x"00",	--920
		x"12",	--921
		x"ce",	--922
		x"4b",	--923
		x"00",	--924
		x"12",	--925
		x"d1",	--926
		x"41",	--927
		x"41",	--928
		x"12",	--929
		x"4f",	--930
		x"4e",	--931
		x"10",	--932
		x"11",	--933
		x"10",	--934
		x"11",	--935
		x"4d",	--936
		x"12",	--937
		x"dd",	--938
		x"4e",	--939
		x"4f",	--940
		x"4b",	--941
		x"12",	--942
		x"ca",	--943
		x"41",	--944
		x"41",	--945
		x"12",	--946
		x"12",	--947
		x"43",	--948
		x"40",	--949
		x"3f",	--950
		x"4a",	--951
		x"4b",	--952
		x"42",	--953
		x"02",	--954
		x"12",	--955
		x"ce",	--956
		x"4a",	--957
		x"4b",	--958
		x"42",	--959
		x"02",	--960
		x"12",	--961
		x"ce",	--962
		x"12",	--963
		x"ef",	--964
		x"12",	--965
		x"d4",	--966
		x"53",	--967
		x"41",	--968
		x"41",	--969
		x"41",	--970
		x"4f",	--971
		x"02",	--972
		x"4e",	--973
		x"02",	--974
		x"41",	--975
		x"12",	--976
		x"12",	--977
		x"83",	--978
		x"4f",	--979
		x"4e",	--980
		x"93",	--981
		x"02",	--982
		x"24",	--983
		x"90",	--984
		x"00",	--985
		x"38",	--986
		x"20",	--987
		x"41",	--988
		x"4b",	--989
		x"00",	--990
		x"12",	--991
		x"cc",	--992
		x"4f",	--993
		x"41",	--994
		x"4b",	--995
		x"00",	--996
		x"12",	--997
		x"cc",	--998
		x"4f",	--999
		x"12",	--1000
		x"12",	--1001
		x"12",	--1002
		x"ef",	--1003
		x"12",	--1004
		x"d4",	--1005
		x"50",	--1006
		x"00",	--1007
		x"4a",	--1008
		x"43",	--1009
		x"12",	--1010
		x"de",	--1011
		x"43",	--1012
		x"40",	--1013
		x"42",	--1014
		x"12",	--1015
		x"db",	--1016
		x"4e",	--1017
		x"4f",	--1018
		x"43",	--1019
		x"40",	--1020
		x"3f",	--1021
		x"12",	--1022
		x"d8",	--1023
		x"4e",	--1024
		x"4f",	--1025
		x"42",	--1026
		x"02",	--1027
		x"12",	--1028
		x"ce",	--1029
		x"4b",	--1030
		x"43",	--1031
		x"12",	--1032
		x"de",	--1033
		x"43",	--1034
		x"40",	--1035
		x"42",	--1036
		x"12",	--1037
		x"db",	--1038
		x"4e",	--1039
		x"4f",	--1040
		x"42",	--1041
		x"02",	--1042
		x"12",	--1043
		x"ce",	--1044
		x"43",	--1045
		x"53",	--1046
		x"41",	--1047
		x"41",	--1048
		x"41",	--1049
		x"41",	--1050
		x"4b",	--1051
		x"00",	--1052
		x"12",	--1053
		x"cc",	--1054
		x"43",	--1055
		x"4f",	--1056
		x"42",	--1057
		x"02",	--1058
		x"12",	--1059
		x"d1",	--1060
		x"3f",	--1061
		x"43",	--1062
		x"40",	--1063
		x"c7",	--1064
		x"12",	--1065
		x"d0",	--1066
		x"4f",	--1067
		x"02",	--1068
		x"3f",	--1069
		x"12",	--1070
		x"ef",	--1071
		x"12",	--1072
		x"d4",	--1073
		x"40",	--1074
		x"ef",	--1075
		x"00",	--1076
		x"12",	--1077
		x"d4",	--1078
		x"4b",	--1079
		x"00",	--1080
		x"12",	--1081
		x"ef",	--1082
		x"12",	--1083
		x"d4",	--1084
		x"52",	--1085
		x"43",	--1086
		x"3f",	--1087
		x"12",	--1088
		x"12",	--1089
		x"42",	--1090
		x"02",	--1091
		x"12",	--1092
		x"d1",	--1093
		x"4e",	--1094
		x"4f",	--1095
		x"42",	--1096
		x"02",	--1097
		x"12",	--1098
		x"d1",	--1099
		x"12",	--1100
		x"12",	--1101
		x"e3",	--1102
		x"e3",	--1103
		x"53",	--1104
		x"63",	--1105
		x"12",	--1106
		x"12",	--1107
		x"12",	--1108
		x"ef",	--1109
		x"12",	--1110
		x"02",	--1111
		x"12",	--1112
		x"e4",	--1113
		x"50",	--1114
		x"00",	--1115
		x"12",	--1116
		x"02",	--1117
		x"12",	--1118
		x"ef",	--1119
		x"12",	--1120
		x"d4",	--1121
		x"52",	--1122
		x"41",	--1123
		x"41",	--1124
		x"41",	--1125
		x"4f",	--1126
		x"02",	--1127
		x"4e",	--1128
		x"02",	--1129
		x"41",	--1130
		x"4f",	--1131
		x"02",	--1132
		x"4e",	--1133
		x"02",	--1134
		x"41",	--1135
		x"12",	--1136
		x"12",	--1137
		x"12",	--1138
		x"12",	--1139
		x"83",	--1140
		x"4f",	--1141
		x"4e",	--1142
		x"43",	--1143
		x"00",	--1144
		x"93",	--1145
		x"24",	--1146
		x"93",	--1147
		x"02",	--1148
		x"24",	--1149
		x"43",	--1150
		x"02",	--1151
		x"41",	--1152
		x"4b",	--1153
		x"00",	--1154
		x"12",	--1155
		x"cc",	--1156
		x"4f",	--1157
		x"90",	--1158
		x"00",	--1159
		x"34",	--1160
		x"43",	--1161
		x"49",	--1162
		x"48",	--1163
		x"42",	--1164
		x"02",	--1165
		x"12",	--1166
		x"d1",	--1167
		x"43",	--1168
		x"53",	--1169
		x"41",	--1170
		x"41",	--1171
		x"41",	--1172
		x"41",	--1173
		x"41",	--1174
		x"93",	--1175
		x"02",	--1176
		x"24",	--1177
		x"43",	--1178
		x"02",	--1179
		x"42",	--1180
		x"02",	--1181
		x"12",	--1182
		x"d1",	--1183
		x"43",	--1184
		x"53",	--1185
		x"41",	--1186
		x"41",	--1187
		x"41",	--1188
		x"41",	--1189
		x"41",	--1190
		x"41",	--1191
		x"4b",	--1192
		x"00",	--1193
		x"12",	--1194
		x"cc",	--1195
		x"4f",	--1196
		x"90",	--1197
		x"00",	--1198
		x"3b",	--1199
		x"41",	--1200
		x"4b",	--1201
		x"00",	--1202
		x"12",	--1203
		x"cc",	--1204
		x"4f",	--1205
		x"41",	--1206
		x"4b",	--1207
		x"00",	--1208
		x"12",	--1209
		x"cc",	--1210
		x"4f",	--1211
		x"12",	--1212
		x"12",	--1213
		x"12",	--1214
		x"ef",	--1215
		x"12",	--1216
		x"d4",	--1217
		x"50",	--1218
		x"00",	--1219
		x"4a",	--1220
		x"43",	--1221
		x"12",	--1222
		x"de",	--1223
		x"43",	--1224
		x"40",	--1225
		x"42",	--1226
		x"12",	--1227
		x"db",	--1228
		x"4e",	--1229
		x"4f",	--1230
		x"42",	--1231
		x"02",	--1232
		x"12",	--1233
		x"ce",	--1234
		x"4b",	--1235
		x"43",	--1236
		x"12",	--1237
		x"de",	--1238
		x"43",	--1239
		x"40",	--1240
		x"42",	--1241
		x"12",	--1242
		x"db",	--1243
		x"4e",	--1244
		x"4f",	--1245
		x"42",	--1246
		x"02",	--1247
		x"12",	--1248
		x"ce",	--1249
		x"3f",	--1250
		x"43",	--1251
		x"12",	--1252
		x"c8",	--1253
		x"43",	--1254
		x"53",	--1255
		x"41",	--1256
		x"41",	--1257
		x"41",	--1258
		x"41",	--1259
		x"41",	--1260
		x"43",	--1261
		x"40",	--1262
		x"c8",	--1263
		x"12",	--1264
		x"d0",	--1265
		x"4f",	--1266
		x"02",	--1267
		x"3f",	--1268
		x"43",	--1269
		x"93",	--1270
		x"02",	--1271
		x"24",	--1272
		x"43",	--1273
		x"4f",	--1274
		x"02",	--1275
		x"43",	--1276
		x"41",	--1277
		x"42",	--1278
		x"00",	--1279
		x"4e",	--1280
		x"be",	--1281
		x"20",	--1282
		x"df",	--1283
		x"00",	--1284
		x"41",	--1285
		x"cf",	--1286
		x"00",	--1287
		x"41",	--1288
		x"42",	--1289
		x"02",	--1290
		x"92",	--1291
		x"2c",	--1292
		x"4e",	--1293
		x"5f",	--1294
		x"4f",	--1295
		x"ef",	--1296
		x"43",	--1297
		x"00",	--1298
		x"90",	--1299
		x"00",	--1300
		x"38",	--1301
		x"43",	--1302
		x"02",	--1303
		x"41",	--1304
		x"53",	--1305
		x"4e",	--1306
		x"02",	--1307
		x"41",	--1308
		x"40",	--1309
		x"00",	--1310
		x"00",	--1311
		x"3f",	--1312
		x"40",	--1313
		x"00",	--1314
		x"00",	--1315
		x"3f",	--1316
		x"42",	--1317
		x"00",	--1318
		x"3f",	--1319
		x"40",	--1320
		x"00",	--1321
		x"00",	--1322
		x"3f",	--1323
		x"40",	--1324
		x"00",	--1325
		x"00",	--1326
		x"3f",	--1327
		x"40",	--1328
		x"00",	--1329
		x"00",	--1330
		x"3f",	--1331
		x"40",	--1332
		x"00",	--1333
		x"00",	--1334
		x"3f",	--1335
		x"4d",	--1336
		x"00",	--1337
		x"4e",	--1338
		x"00",	--1339
		x"41",	--1340
		x"00",	--1341
		x"00",	--1342
		x"41",	--1343
		x"00",	--1344
		x"00",	--1345
		x"41",	--1346
		x"00",	--1347
		x"00",	--1348
		x"41",	--1349
		x"00",	--1350
		x"00",	--1351
		x"41",	--1352
		x"00",	--1353
		x"00",	--1354
		x"41",	--1355
		x"00",	--1356
		x"00",	--1357
		x"43",	--1358
		x"00",	--1359
		x"43",	--1360
		x"00",	--1361
		x"43",	--1362
		x"00",	--1363
		x"43",	--1364
		x"00",	--1365
		x"43",	--1366
		x"00",	--1367
		x"43",	--1368
		x"00",	--1369
		x"43",	--1370
		x"00",	--1371
		x"43",	--1372
		x"00",	--1373
		x"41",	--1374
		x"43",	--1375
		x"00",	--1376
		x"43",	--1377
		x"00",	--1378
		x"43",	--1379
		x"00",	--1380
		x"43",	--1381
		x"00",	--1382
		x"43",	--1383
		x"00",	--1384
		x"43",	--1385
		x"00",	--1386
		x"41",	--1387
		x"4d",	--1388
		x"00",	--1389
		x"4e",	--1390
		x"00",	--1391
		x"41",	--1392
		x"4d",	--1393
		x"00",	--1394
		x"4e",	--1395
		x"00",	--1396
		x"41",	--1397
		x"4d",	--1398
		x"00",	--1399
		x"4e",	--1400
		x"00",	--1401
		x"41",	--1402
		x"4d",	--1403
		x"00",	--1404
		x"4e",	--1405
		x"00",	--1406
		x"41",	--1407
		x"4d",	--1408
		x"00",	--1409
		x"4e",	--1410
		x"00",	--1411
		x"41",	--1412
		x"12",	--1413
		x"12",	--1414
		x"12",	--1415
		x"12",	--1416
		x"12",	--1417
		x"12",	--1418
		x"12",	--1419
		x"4f",	--1420
		x"4d",	--1421
		x"4e",	--1422
		x"4f",	--1423
		x"00",	--1424
		x"4f",	--1425
		x"00",	--1426
		x"4f",	--1427
		x"00",	--1428
		x"4f",	--1429
		x"00",	--1430
		x"4a",	--1431
		x"4b",	--1432
		x"46",	--1433
		x"47",	--1434
		x"12",	--1435
		x"dd",	--1436
		x"49",	--1437
		x"00",	--1438
		x"49",	--1439
		x"00",	--1440
		x"93",	--1441
		x"34",	--1442
		x"46",	--1443
		x"47",	--1444
		x"12",	--1445
		x"d8",	--1446
		x"4e",	--1447
		x"4f",	--1448
		x"4e",	--1449
		x"00",	--1450
		x"4f",	--1451
		x"00",	--1452
		x"4e",	--1453
		x"4f",	--1454
		x"4a",	--1455
		x"4b",	--1456
		x"12",	--1457
		x"dd",	--1458
		x"93",	--1459
		x"34",	--1460
		x"4a",	--1461
		x"00",	--1462
		x"4b",	--1463
		x"00",	--1464
		x"44",	--1465
		x"45",	--1466
		x"4a",	--1467
		x"4b",	--1468
		x"12",	--1469
		x"d8",	--1470
		x"4e",	--1471
		x"4f",	--1472
		x"49",	--1473
		x"00",	--1474
		x"49",	--1475
		x"00",	--1476
		x"12",	--1477
		x"d8",	--1478
		x"4e",	--1479
		x"4f",	--1480
		x"4e",	--1481
		x"00",	--1482
		x"4f",	--1483
		x"00",	--1484
		x"49",	--1485
		x"49",	--1486
		x"00",	--1487
		x"4a",	--1488
		x"4b",	--1489
		x"12",	--1490
		x"d9",	--1491
		x"4e",	--1492
		x"4f",	--1493
		x"49",	--1494
		x"00",	--1495
		x"49",	--1496
		x"00",	--1497
		x"46",	--1498
		x"47",	--1499
		x"12",	--1500
		x"d9",	--1501
		x"44",	--1502
		x"45",	--1503
		x"12",	--1504
		x"d8",	--1505
		x"4e",	--1506
		x"4f",	--1507
		x"49",	--1508
		x"00",	--1509
		x"49",	--1510
		x"00",	--1511
		x"4a",	--1512
		x"4b",	--1513
		x"12",	--1514
		x"d8",	--1515
		x"49",	--1516
		x"00",	--1517
		x"49",	--1518
		x"00",	--1519
		x"12",	--1520
		x"d9",	--1521
		x"46",	--1522
		x"47",	--1523
		x"12",	--1524
		x"d8",	--1525
		x"41",	--1526
		x"41",	--1527
		x"41",	--1528
		x"41",	--1529
		x"41",	--1530
		x"41",	--1531
		x"41",	--1532
		x"41",	--1533
		x"46",	--1534
		x"47",	--1535
		x"12",	--1536
		x"d8",	--1537
		x"4e",	--1538
		x"4f",	--1539
		x"4e",	--1540
		x"00",	--1541
		x"4f",	--1542
		x"00",	--1543
		x"4e",	--1544
		x"4f",	--1545
		x"4a",	--1546
		x"4b",	--1547
		x"12",	--1548
		x"dc",	--1549
		x"93",	--1550
		x"24",	--1551
		x"37",	--1552
		x"46",	--1553
		x"47",	--1554
		x"3f",	--1555
		x"12",	--1556
		x"12",	--1557
		x"83",	--1558
		x"4f",	--1559
		x"4e",	--1560
		x"12",	--1561
		x"f0",	--1562
		x"12",	--1563
		x"d4",	--1564
		x"53",	--1565
		x"90",	--1566
		x"00",	--1567
		x"38",	--1568
		x"41",	--1569
		x"4b",	--1570
		x"00",	--1571
		x"12",	--1572
		x"cc",	--1573
		x"4f",	--1574
		x"41",	--1575
		x"4b",	--1576
		x"00",	--1577
		x"12",	--1578
		x"cc",	--1579
		x"4f",	--1580
		x"12",	--1581
		x"12",	--1582
		x"12",	--1583
		x"f0",	--1584
		x"12",	--1585
		x"d4",	--1586
		x"50",	--1587
		x"00",	--1588
		x"4b",	--1589
		x"00",	--1590
		x"43",	--1591
		x"53",	--1592
		x"41",	--1593
		x"41",	--1594
		x"41",	--1595
		x"12",	--1596
		x"f0",	--1597
		x"12",	--1598
		x"d4",	--1599
		x"40",	--1600
		x"f0",	--1601
		x"00",	--1602
		x"12",	--1603
		x"d4",	--1604
		x"4b",	--1605
		x"00",	--1606
		x"12",	--1607
		x"f0",	--1608
		x"12",	--1609
		x"d4",	--1610
		x"52",	--1611
		x"43",	--1612
		x"3f",	--1613
		x"12",	--1614
		x"83",	--1615
		x"4e",	--1616
		x"93",	--1617
		x"24",	--1618
		x"38",	--1619
		x"12",	--1620
		x"f0",	--1621
		x"12",	--1622
		x"d4",	--1623
		x"53",	--1624
		x"41",	--1625
		x"4b",	--1626
		x"00",	--1627
		x"12",	--1628
		x"cc",	--1629
		x"12",	--1630
		x"12",	--1631
		x"12",	--1632
		x"f0",	--1633
		x"12",	--1634
		x"d4",	--1635
		x"50",	--1636
		x"00",	--1637
		x"43",	--1638
		x"53",	--1639
		x"41",	--1640
		x"41",	--1641
		x"12",	--1642
		x"f0",	--1643
		x"12",	--1644
		x"d4",	--1645
		x"40",	--1646
		x"f0",	--1647
		x"00",	--1648
		x"12",	--1649
		x"d4",	--1650
		x"4b",	--1651
		x"00",	--1652
		x"12",	--1653
		x"f0",	--1654
		x"12",	--1655
		x"d4",	--1656
		x"52",	--1657
		x"43",	--1658
		x"3f",	--1659
		x"12",	--1660
		x"12",	--1661
		x"43",	--1662
		x"00",	--1663
		x"4f",	--1664
		x"93",	--1665
		x"24",	--1666
		x"53",	--1667
		x"43",	--1668
		x"43",	--1669
		x"3c",	--1670
		x"90",	--1671
		x"00",	--1672
		x"2c",	--1673
		x"5c",	--1674
		x"5c",	--1675
		x"5c",	--1676
		x"5c",	--1677
		x"11",	--1678
		x"5d",	--1679
		x"50",	--1680
		x"ff",	--1681
		x"43",	--1682
		x"4f",	--1683
		x"93",	--1684
		x"24",	--1685
		x"90",	--1686
		x"00",	--1687
		x"24",	--1688
		x"4d",	--1689
		x"50",	--1690
		x"ff",	--1691
		x"93",	--1692
		x"23",	--1693
		x"90",	--1694
		x"00",	--1695
		x"2c",	--1696
		x"5c",	--1697
		x"4c",	--1698
		x"5b",	--1699
		x"5b",	--1700
		x"5b",	--1701
		x"11",	--1702
		x"5d",	--1703
		x"50",	--1704
		x"ff",	--1705
		x"4f",	--1706
		x"93",	--1707
		x"23",	--1708
		x"43",	--1709
		x"00",	--1710
		x"4c",	--1711
		x"41",	--1712
		x"41",	--1713
		x"41",	--1714
		x"43",	--1715
		x"3f",	--1716
		x"4d",	--1717
		x"50",	--1718
		x"ff",	--1719
		x"90",	--1720
		x"00",	--1721
		x"2c",	--1722
		x"5c",	--1723
		x"5c",	--1724
		x"5c",	--1725
		x"5c",	--1726
		x"11",	--1727
		x"5d",	--1728
		x"50",	--1729
		x"ff",	--1730
		x"43",	--1731
		x"3f",	--1732
		x"4d",	--1733
		x"50",	--1734
		x"ff",	--1735
		x"90",	--1736
		x"00",	--1737
		x"2c",	--1738
		x"5c",	--1739
		x"5c",	--1740
		x"5c",	--1741
		x"5c",	--1742
		x"11",	--1743
		x"5d",	--1744
		x"50",	--1745
		x"ff",	--1746
		x"43",	--1747
		x"3f",	--1748
		x"11",	--1749
		x"12",	--1750
		x"12",	--1751
		x"f0",	--1752
		x"12",	--1753
		x"d4",	--1754
		x"52",	--1755
		x"43",	--1756
		x"4c",	--1757
		x"41",	--1758
		x"41",	--1759
		x"41",	--1760
		x"43",	--1761
		x"3f",	--1762
		x"12",	--1763
		x"12",	--1764
		x"43",	--1765
		x"00",	--1766
		x"4f",	--1767
		x"93",	--1768
		x"24",	--1769
		x"53",	--1770
		x"43",	--1771
		x"43",	--1772
		x"3c",	--1773
		x"4b",	--1774
		x"50",	--1775
		x"ff",	--1776
		x"90",	--1777
		x"00",	--1778
		x"2c",	--1779
		x"5c",	--1780
		x"4c",	--1781
		x"5d",	--1782
		x"5d",	--1783
		x"5d",	--1784
		x"11",	--1785
		x"5b",	--1786
		x"50",	--1787
		x"ff",	--1788
		x"4f",	--1789
		x"93",	--1790
		x"24",	--1791
		x"90",	--1792
		x"00",	--1793
		x"23",	--1794
		x"43",	--1795
		x"4f",	--1796
		x"93",	--1797
		x"23",	--1798
		x"12",	--1799
		x"c2",	--1800
		x"43",	--1801
		x"4a",	--1802
		x"01",	--1803
		x"4c",	--1804
		x"01",	--1805
		x"42",	--1806
		x"01",	--1807
		x"41",	--1808
		x"43",	--1809
		x"00",	--1810
		x"41",	--1811
		x"41",	--1812
		x"41",	--1813
		x"11",	--1814
		x"12",	--1815
		x"12",	--1816
		x"f0",	--1817
		x"12",	--1818
		x"d4",	--1819
		x"52",	--1820
		x"43",	--1821
		x"41",	--1822
		x"41",	--1823
		x"41",	--1824
		x"43",	--1825
		x"3f",	--1826
		x"12",	--1827
		x"12",	--1828
		x"4e",	--1829
		x"4c",	--1830
		x"4e",	--1831
		x"00",	--1832
		x"4d",	--1833
		x"00",	--1834
		x"4c",	--1835
		x"00",	--1836
		x"4d",	--1837
		x"43",	--1838
		x"40",	--1839
		x"36",	--1840
		x"40",	--1841
		x"01",	--1842
		x"12",	--1843
		x"ed",	--1844
		x"4e",	--1845
		x"00",	--1846
		x"12",	--1847
		x"c2",	--1848
		x"43",	--1849
		x"4a",	--1850
		x"01",	--1851
		x"40",	--1852
		x"00",	--1853
		x"01",	--1854
		x"42",	--1855
		x"01",	--1856
		x"00",	--1857
		x"41",	--1858
		x"43",	--1859
		x"41",	--1860
		x"41",	--1861
		x"41",	--1862
		x"12",	--1863
		x"12",	--1864
		x"12",	--1865
		x"43",	--1866
		x"00",	--1867
		x"40",	--1868
		x"3f",	--1869
		x"00",	--1870
		x"4f",	--1871
		x"4b",	--1872
		x"00",	--1873
		x"43",	--1874
		x"12",	--1875
		x"de",	--1876
		x"43",	--1877
		x"40",	--1878
		x"3f",	--1879
		x"12",	--1880
		x"d9",	--1881
		x"4e",	--1882
		x"4f",	--1883
		x"4b",	--1884
		x"00",	--1885
		x"43",	--1886
		x"12",	--1887
		x"de",	--1888
		x"4e",	--1889
		x"4f",	--1890
		x"48",	--1891
		x"49",	--1892
		x"12",	--1893
		x"d8",	--1894
		x"12",	--1895
		x"d5",	--1896
		x"4e",	--1897
		x"00",	--1898
		x"43",	--1899
		x"00",	--1900
		x"41",	--1901
		x"41",	--1902
		x"41",	--1903
		x"41",	--1904
		x"12",	--1905
		x"12",	--1906
		x"12",	--1907
		x"4d",	--1908
		x"4e",	--1909
		x"4d",	--1910
		x"00",	--1911
		x"4e",	--1912
		x"00",	--1913
		x"4f",	--1914
		x"49",	--1915
		x"00",	--1916
		x"43",	--1917
		x"12",	--1918
		x"de",	--1919
		x"4e",	--1920
		x"4f",	--1921
		x"4a",	--1922
		x"4b",	--1923
		x"12",	--1924
		x"d9",	--1925
		x"4e",	--1926
		x"4f",	--1927
		x"49",	--1928
		x"00",	--1929
		x"43",	--1930
		x"12",	--1931
		x"de",	--1932
		x"4e",	--1933
		x"4f",	--1934
		x"4a",	--1935
		x"4b",	--1936
		x"12",	--1937
		x"d8",	--1938
		x"12",	--1939
		x"d5",	--1940
		x"4e",	--1941
		x"00",	--1942
		x"41",	--1943
		x"41",	--1944
		x"41",	--1945
		x"41",	--1946
		x"4f",	--1947
		x"4e",	--1948
		x"00",	--1949
		x"41",	--1950
		x"12",	--1951
		x"12",	--1952
		x"93",	--1953
		x"02",	--1954
		x"38",	--1955
		x"40",	--1956
		x"02",	--1957
		x"43",	--1958
		x"12",	--1959
		x"4b",	--1960
		x"ff",	--1961
		x"11",	--1962
		x"12",	--1963
		x"12",	--1964
		x"f0",	--1965
		x"12",	--1966
		x"d4",	--1967
		x"50",	--1968
		x"00",	--1969
		x"53",	--1970
		x"50",	--1971
		x"00",	--1972
		x"92",	--1973
		x"02",	--1974
		x"3b",	--1975
		x"43",	--1976
		x"41",	--1977
		x"41",	--1978
		x"41",	--1979
		x"42",	--1980
		x"02",	--1981
		x"90",	--1982
		x"00",	--1983
		x"34",	--1984
		x"4e",	--1985
		x"5f",	--1986
		x"5e",	--1987
		x"5f",	--1988
		x"50",	--1989
		x"02",	--1990
		x"40",	--1991
		x"00",	--1992
		x"00",	--1993
		x"40",	--1994
		x"cf",	--1995
		x"00",	--1996
		x"40",	--1997
		x"02",	--1998
		x"00",	--1999
		x"53",	--2000
		x"4e",	--2001
		x"02",	--2002
		x"41",	--2003
		x"12",	--2004
		x"42",	--2005
		x"02",	--2006
		x"90",	--2007
		x"00",	--2008
		x"34",	--2009
		x"4b",	--2010
		x"5c",	--2011
		x"5b",	--2012
		x"5c",	--2013
		x"50",	--2014
		x"02",	--2015
		x"4f",	--2016
		x"00",	--2017
		x"4e",	--2018
		x"00",	--2019
		x"4d",	--2020
		x"00",	--2021
		x"53",	--2022
		x"4b",	--2023
		x"02",	--2024
		x"43",	--2025
		x"41",	--2026
		x"41",	--2027
		x"43",	--2028
		x"3f",	--2029
		x"12",	--2030
		x"50",	--2031
		x"ff",	--2032
		x"42",	--2033
		x"02",	--2034
		x"93",	--2035
		x"38",	--2036
		x"92",	--2037
		x"02",	--2038
		x"24",	--2039
		x"40",	--2040
		x"02",	--2041
		x"43",	--2042
		x"3c",	--2043
		x"50",	--2044
		x"00",	--2045
		x"9f",	--2046
		x"ff",	--2047
		x"24",	--2048
		x"53",	--2049
		x"9b",	--2050
		x"23",	--2051
		x"12",	--2052
		x"f0",	--2053
		x"12",	--2054
		x"d4",	--2055
		x"53",	--2056
		x"43",	--2057
		x"50",	--2058
		x"00",	--2059
		x"41",	--2060
		x"41",	--2061
		x"43",	--2062
		x"4e",	--2063
		x"00",	--2064
		x"4e",	--2065
		x"93",	--2066
		x"24",	--2067
		x"53",	--2068
		x"43",	--2069
		x"3c",	--2070
		x"4e",	--2071
		x"93",	--2072
		x"24",	--2073
		x"53",	--2074
		x"92",	--2075
		x"34",	--2076
		x"90",	--2077
		x"00",	--2078
		x"23",	--2079
		x"43",	--2080
		x"ff",	--2081
		x"4f",	--2082
		x"5d",	--2083
		x"51",	--2084
		x"4e",	--2085
		x"00",	--2086
		x"53",	--2087
		x"4e",	--2088
		x"93",	--2089
		x"23",	--2090
		x"4c",	--2091
		x"5e",	--2092
		x"5e",	--2093
		x"5c",	--2094
		x"50",	--2095
		x"02",	--2096
		x"41",	--2097
		x"12",	--2098
		x"00",	--2099
		x"50",	--2100
		x"00",	--2101
		x"41",	--2102
		x"41",	--2103
		x"43",	--2104
		x"3f",	--2105
		x"4e",	--2106
		x"00",	--2107
		x"43",	--2108
		x"41",	--2109
		x"5e",	--2110
		x"5f",	--2111
		x"4e",	--2112
		x"41",	--2113
		x"12",	--2114
		x"12",	--2115
		x"5e",	--2116
		x"5f",	--2117
		x"4e",	--2118
		x"43",	--2119
		x"4c",	--2120
		x"4d",	--2121
		x"5e",	--2122
		x"6f",	--2123
		x"4e",	--2124
		x"4f",	--2125
		x"5a",	--2126
		x"6b",	--2127
		x"5a",	--2128
		x"6b",	--2129
		x"40",	--2130
		x"00",	--2131
		x"43",	--2132
		x"5a",	--2133
		x"6b",	--2134
		x"12",	--2135
		x"ec",	--2136
		x"4e",	--2137
		x"41",	--2138
		x"41",	--2139
		x"41",	--2140
		x"d0",	--2141
		x"02",	--2142
		x"01",	--2143
		x"40",	--2144
		x"0b",	--2145
		x"01",	--2146
		x"43",	--2147
		x"41",	--2148
		x"12",	--2149
		x"4f",	--2150
		x"42",	--2151
		x"02",	--2152
		x"90",	--2153
		x"00",	--2154
		x"34",	--2155
		x"4f",	--2156
		x"5c",	--2157
		x"4c",	--2158
		x"5d",	--2159
		x"5d",	--2160
		x"5d",	--2161
		x"8c",	--2162
		x"50",	--2163
		x"03",	--2164
		x"43",	--2165
		x"00",	--2166
		x"43",	--2167
		x"00",	--2168
		x"43",	--2169
		x"00",	--2170
		x"4b",	--2171
		x"00",	--2172
		x"4e",	--2173
		x"00",	--2174
		x"4f",	--2175
		x"53",	--2176
		x"4e",	--2177
		x"02",	--2178
		x"41",	--2179
		x"41",	--2180
		x"43",	--2181
		x"3f",	--2182
		x"5f",	--2183
		x"4f",	--2184
		x"5c",	--2185
		x"5c",	--2186
		x"5c",	--2187
		x"8f",	--2188
		x"50",	--2189
		x"03",	--2190
		x"43",	--2191
		x"00",	--2192
		x"4e",	--2193
		x"00",	--2194
		x"43",	--2195
		x"00",	--2196
		x"4d",	--2197
		x"00",	--2198
		x"43",	--2199
		x"00",	--2200
		x"43",	--2201
		x"41",	--2202
		x"5f",	--2203
		x"4f",	--2204
		x"5e",	--2205
		x"5e",	--2206
		x"5e",	--2207
		x"8f",	--2208
		x"43",	--2209
		x"03",	--2210
		x"43",	--2211
		x"41",	--2212
		x"12",	--2213
		x"12",	--2214
		x"12",	--2215
		x"12",	--2216
		x"12",	--2217
		x"12",	--2218
		x"12",	--2219
		x"12",	--2220
		x"12",	--2221
		x"93",	--2222
		x"02",	--2223
		x"38",	--2224
		x"40",	--2225
		x"03",	--2226
		x"4a",	--2227
		x"53",	--2228
		x"4a",	--2229
		x"52",	--2230
		x"4a",	--2231
		x"50",	--2232
		x"00",	--2233
		x"43",	--2234
		x"3c",	--2235
		x"53",	--2236
		x"4f",	--2237
		x"00",	--2238
		x"53",	--2239
		x"50",	--2240
		x"00",	--2241
		x"50",	--2242
		x"00",	--2243
		x"50",	--2244
		x"00",	--2245
		x"50",	--2246
		x"00",	--2247
		x"92",	--2248
		x"02",	--2249
		x"34",	--2250
		x"93",	--2251
		x"00",	--2252
		x"27",	--2253
		x"4b",	--2254
		x"9b",	--2255
		x"00",	--2256
		x"2b",	--2257
		x"43",	--2258
		x"00",	--2259
		x"4b",	--2260
		x"00",	--2261
		x"12",	--2262
		x"00",	--2263
		x"93",	--2264
		x"00",	--2265
		x"27",	--2266
		x"47",	--2267
		x"53",	--2268
		x"4f",	--2269
		x"00",	--2270
		x"98",	--2271
		x"2b",	--2272
		x"43",	--2273
		x"00",	--2274
		x"3f",	--2275
		x"f0",	--2276
		x"ff",	--2277
		x"01",	--2278
		x"41",	--2279
		x"41",	--2280
		x"41",	--2281
		x"41",	--2282
		x"41",	--2283
		x"41",	--2284
		x"41",	--2285
		x"41",	--2286
		x"41",	--2287
		x"13",	--2288
		x"4e",	--2289
		x"00",	--2290
		x"43",	--2291
		x"41",	--2292
		x"4f",	--2293
		x"4f",	--2294
		x"4f",	--2295
		x"00",	--2296
		x"41",	--2297
		x"43",	--2298
		x"00",	--2299
		x"41",	--2300
		x"4e",	--2301
		x"00",	--2302
		x"40",	--2303
		x"d1",	--2304
		x"12",	--2305
		x"d0",	--2306
		x"4f",	--2307
		x"02",	--2308
		x"43",	--2309
		x"41",	--2310
		x"4d",	--2311
		x"4f",	--2312
		x"4e",	--2313
		x"00",	--2314
		x"43",	--2315
		x"4c",	--2316
		x"42",	--2317
		x"02",	--2318
		x"12",	--2319
		x"d1",	--2320
		x"41",	--2321
		x"42",	--2322
		x"00",	--2323
		x"f2",	--2324
		x"23",	--2325
		x"4f",	--2326
		x"00",	--2327
		x"43",	--2328
		x"41",	--2329
		x"f0",	--2330
		x"00",	--2331
		x"4f",	--2332
		x"f1",	--2333
		x"11",	--2334
		x"12",	--2335
		x"d2",	--2336
		x"41",	--2337
		x"12",	--2338
		x"4f",	--2339
		x"4f",	--2340
		x"11",	--2341
		x"11",	--2342
		x"11",	--2343
		x"11",	--2344
		x"4e",	--2345
		x"12",	--2346
		x"d2",	--2347
		x"4b",	--2348
		x"12",	--2349
		x"d2",	--2350
		x"41",	--2351
		x"41",	--2352
		x"12",	--2353
		x"12",	--2354
		x"4f",	--2355
		x"40",	--2356
		x"00",	--2357
		x"4a",	--2358
		x"4b",	--2359
		x"f0",	--2360
		x"00",	--2361
		x"24",	--2362
		x"11",	--2363
		x"53",	--2364
		x"23",	--2365
		x"f3",	--2366
		x"24",	--2367
		x"40",	--2368
		x"00",	--2369
		x"12",	--2370
		x"d2",	--2371
		x"53",	--2372
		x"93",	--2373
		x"23",	--2374
		x"41",	--2375
		x"41",	--2376
		x"41",	--2377
		x"40",	--2378
		x"00",	--2379
		x"3f",	--2380
		x"12",	--2381
		x"4f",	--2382
		x"4f",	--2383
		x"10",	--2384
		x"11",	--2385
		x"4e",	--2386
		x"12",	--2387
		x"d2",	--2388
		x"4b",	--2389
		x"12",	--2390
		x"d2",	--2391
		x"41",	--2392
		x"41",	--2393
		x"12",	--2394
		x"12",	--2395
		x"4e",	--2396
		x"4f",	--2397
		x"4f",	--2398
		x"10",	--2399
		x"11",	--2400
		x"4d",	--2401
		x"12",	--2402
		x"d2",	--2403
		x"4b",	--2404
		x"12",	--2405
		x"d2",	--2406
		x"4b",	--2407
		x"4a",	--2408
		x"10",	--2409
		x"10",	--2410
		x"ec",	--2411
		x"ec",	--2412
		x"4d",	--2413
		x"12",	--2414
		x"d2",	--2415
		x"4a",	--2416
		x"12",	--2417
		x"d2",	--2418
		x"41",	--2419
		x"41",	--2420
		x"41",	--2421
		x"12",	--2422
		x"12",	--2423
		x"12",	--2424
		x"4f",	--2425
		x"93",	--2426
		x"24",	--2427
		x"4e",	--2428
		x"53",	--2429
		x"43",	--2430
		x"4a",	--2431
		x"5b",	--2432
		x"4d",	--2433
		x"11",	--2434
		x"12",	--2435
		x"d2",	--2436
		x"99",	--2437
		x"24",	--2438
		x"53",	--2439
		x"b0",	--2440
		x"00",	--2441
		x"20",	--2442
		x"40",	--2443
		x"00",	--2444
		x"12",	--2445
		x"d2",	--2446
		x"3f",	--2447
		x"40",	--2448
		x"00",	--2449
		x"12",	--2450
		x"d2",	--2451
		x"3f",	--2452
		x"41",	--2453
		x"41",	--2454
		x"41",	--2455
		x"41",	--2456
		x"12",	--2457
		x"12",	--2458
		x"12",	--2459
		x"4f",	--2460
		x"93",	--2461
		x"24",	--2462
		x"4e",	--2463
		x"53",	--2464
		x"43",	--2465
		x"4a",	--2466
		x"11",	--2467
		x"12",	--2468
		x"d2",	--2469
		x"99",	--2470
		x"24",	--2471
		x"53",	--2472
		x"b0",	--2473
		x"00",	--2474
		x"23",	--2475
		x"40",	--2476
		x"00",	--2477
		x"12",	--2478
		x"d2",	--2479
		x"4a",	--2480
		x"11",	--2481
		x"12",	--2482
		x"d2",	--2483
		x"99",	--2484
		x"23",	--2485
		x"41",	--2486
		x"41",	--2487
		x"41",	--2488
		x"41",	--2489
		x"12",	--2490
		x"12",	--2491
		x"12",	--2492
		x"50",	--2493
		x"ff",	--2494
		x"4f",	--2495
		x"93",	--2496
		x"38",	--2497
		x"90",	--2498
		x"00",	--2499
		x"38",	--2500
		x"43",	--2501
		x"41",	--2502
		x"59",	--2503
		x"40",	--2504
		x"00",	--2505
		x"4b",	--2506
		x"12",	--2507
		x"ec",	--2508
		x"50",	--2509
		x"00",	--2510
		x"4f",	--2511
		x"00",	--2512
		x"53",	--2513
		x"40",	--2514
		x"00",	--2515
		x"4b",	--2516
		x"12",	--2517
		x"ec",	--2518
		x"4f",	--2519
		x"90",	--2520
		x"00",	--2521
		x"37",	--2522
		x"49",	--2523
		x"53",	--2524
		x"51",	--2525
		x"40",	--2526
		x"00",	--2527
		x"4b",	--2528
		x"12",	--2529
		x"ec",	--2530
		x"50",	--2531
		x"00",	--2532
		x"4f",	--2533
		x"00",	--2534
		x"53",	--2535
		x"41",	--2536
		x"5a",	--2537
		x"4f",	--2538
		x"11",	--2539
		x"12",	--2540
		x"d2",	--2541
		x"93",	--2542
		x"23",	--2543
		x"50",	--2544
		x"00",	--2545
		x"41",	--2546
		x"41",	--2547
		x"41",	--2548
		x"41",	--2549
		x"40",	--2550
		x"00",	--2551
		x"12",	--2552
		x"d2",	--2553
		x"e3",	--2554
		x"53",	--2555
		x"3f",	--2556
		x"43",	--2557
		x"43",	--2558
		x"3f",	--2559
		x"12",	--2560
		x"12",	--2561
		x"12",	--2562
		x"41",	--2563
		x"52",	--2564
		x"4b",	--2565
		x"49",	--2566
		x"93",	--2567
		x"20",	--2568
		x"3c",	--2569
		x"11",	--2570
		x"12",	--2571
		x"d2",	--2572
		x"49",	--2573
		x"4a",	--2574
		x"53",	--2575
		x"4a",	--2576
		x"00",	--2577
		x"93",	--2578
		x"24",	--2579
		x"90",	--2580
		x"00",	--2581
		x"23",	--2582
		x"49",	--2583
		x"53",	--2584
		x"49",	--2585
		x"00",	--2586
		x"50",	--2587
		x"ff",	--2588
		x"90",	--2589
		x"00",	--2590
		x"2f",	--2591
		x"4f",	--2592
		x"5f",	--2593
		x"4f",	--2594
		x"f0",	--2595
		x"41",	--2596
		x"41",	--2597
		x"41",	--2598
		x"41",	--2599
		x"4b",	--2600
		x"52",	--2601
		x"4b",	--2602
		x"00",	--2603
		x"4b",	--2604
		x"12",	--2605
		x"d2",	--2606
		x"49",	--2607
		x"3f",	--2608
		x"4b",	--2609
		x"53",	--2610
		x"4b",	--2611
		x"12",	--2612
		x"d2",	--2613
		x"49",	--2614
		x"3f",	--2615
		x"4b",	--2616
		x"53",	--2617
		x"4f",	--2618
		x"49",	--2619
		x"93",	--2620
		x"27",	--2621
		x"53",	--2622
		x"11",	--2623
		x"12",	--2624
		x"d2",	--2625
		x"49",	--2626
		x"93",	--2627
		x"23",	--2628
		x"3f",	--2629
		x"4b",	--2630
		x"52",	--2631
		x"4b",	--2632
		x"00",	--2633
		x"4b",	--2634
		x"12",	--2635
		x"d3",	--2636
		x"49",	--2637
		x"3f",	--2638
		x"4b",	--2639
		x"53",	--2640
		x"4b",	--2641
		x"4e",	--2642
		x"10",	--2643
		x"11",	--2644
		x"10",	--2645
		x"11",	--2646
		x"12",	--2647
		x"d2",	--2648
		x"49",	--2649
		x"3f",	--2650
		x"4b",	--2651
		x"53",	--2652
		x"4b",	--2653
		x"12",	--2654
		x"d3",	--2655
		x"49",	--2656
		x"3f",	--2657
		x"4b",	--2658
		x"53",	--2659
		x"4b",	--2660
		x"12",	--2661
		x"d2",	--2662
		x"49",	--2663
		x"3f",	--2664
		x"4b",	--2665
		x"53",	--2666
		x"4b",	--2667
		x"12",	--2668
		x"d2",	--2669
		x"49",	--2670
		x"3f",	--2671
		x"4b",	--2672
		x"53",	--2673
		x"4b",	--2674
		x"12",	--2675
		x"d2",	--2676
		x"49",	--2677
		x"3f",	--2678
		x"40",	--2679
		x"00",	--2680
		x"12",	--2681
		x"d2",	--2682
		x"3f",	--2683
		x"12",	--2684
		x"12",	--2685
		x"42",	--2686
		x"02",	--2687
		x"42",	--2688
		x"00",	--2689
		x"04",	--2690
		x"42",	--2691
		x"02",	--2692
		x"90",	--2693
		x"00",	--2694
		x"34",	--2695
		x"53",	--2696
		x"02",	--2697
		x"42",	--2698
		x"02",	--2699
		x"42",	--2700
		x"02",	--2701
		x"9f",	--2702
		x"20",	--2703
		x"53",	--2704
		x"02",	--2705
		x"40",	--2706
		x"00",	--2707
		x"00",	--2708
		x"41",	--2709
		x"41",	--2710
		x"c0",	--2711
		x"00",	--2712
		x"00",	--2713
		x"13",	--2714
		x"43",	--2715
		x"02",	--2716
		x"3f",	--2717
		x"4e",	--2718
		x"4f",	--2719
		x"40",	--2720
		x"36",	--2721
		x"40",	--2722
		x"01",	--2723
		x"12",	--2724
		x"ec",	--2725
		x"53",	--2726
		x"4e",	--2727
		x"00",	--2728
		x"40",	--2729
		x"00",	--2730
		x"00",	--2731
		x"41",	--2732
		x"42",	--2733
		x"02",	--2734
		x"42",	--2735
		x"02",	--2736
		x"9f",	--2737
		x"38",	--2738
		x"42",	--2739
		x"02",	--2740
		x"82",	--2741
		x"02",	--2742
		x"41",	--2743
		x"42",	--2744
		x"02",	--2745
		x"42",	--2746
		x"02",	--2747
		x"40",	--2748
		x"00",	--2749
		x"8d",	--2750
		x"8e",	--2751
		x"41",	--2752
		x"42",	--2753
		x"02",	--2754
		x"4f",	--2755
		x"04",	--2756
		x"42",	--2757
		x"02",	--2758
		x"42",	--2759
		x"02",	--2760
		x"9e",	--2761
		x"24",	--2762
		x"42",	--2763
		x"02",	--2764
		x"90",	--2765
		x"00",	--2766
		x"38",	--2767
		x"43",	--2768
		x"02",	--2769
		x"41",	--2770
		x"53",	--2771
		x"02",	--2772
		x"41",	--2773
		x"43",	--2774
		x"41",	--2775
		x"12",	--2776
		x"12",	--2777
		x"4e",	--2778
		x"4f",	--2779
		x"43",	--2780
		x"40",	--2781
		x"4f",	--2782
		x"12",	--2783
		x"dc",	--2784
		x"93",	--2785
		x"34",	--2786
		x"4a",	--2787
		x"4b",	--2788
		x"12",	--2789
		x"de",	--2790
		x"41",	--2791
		x"41",	--2792
		x"41",	--2793
		x"43",	--2794
		x"40",	--2795
		x"4f",	--2796
		x"4a",	--2797
		x"4b",	--2798
		x"12",	--2799
		x"d8",	--2800
		x"12",	--2801
		x"de",	--2802
		x"53",	--2803
		x"60",	--2804
		x"80",	--2805
		x"41",	--2806
		x"41",	--2807
		x"41",	--2808
		x"12",	--2809
		x"12",	--2810
		x"12",	--2811
		x"12",	--2812
		x"12",	--2813
		x"12",	--2814
		x"12",	--2815
		x"12",	--2816
		x"50",	--2817
		x"ff",	--2818
		x"4d",	--2819
		x"4f",	--2820
		x"93",	--2821
		x"28",	--2822
		x"4e",	--2823
		x"93",	--2824
		x"28",	--2825
		x"92",	--2826
		x"20",	--2827
		x"40",	--2828
		x"d8",	--2829
		x"92",	--2830
		x"24",	--2831
		x"93",	--2832
		x"24",	--2833
		x"93",	--2834
		x"24",	--2835
		x"4f",	--2836
		x"00",	--2837
		x"00",	--2838
		x"4e",	--2839
		x"00",	--2840
		x"4f",	--2841
		x"00",	--2842
		x"4f",	--2843
		x"00",	--2844
		x"4e",	--2845
		x"00",	--2846
		x"4e",	--2847
		x"00",	--2848
		x"41",	--2849
		x"8b",	--2850
		x"4c",	--2851
		x"93",	--2852
		x"38",	--2853
		x"90",	--2854
		x"00",	--2855
		x"34",	--2856
		x"93",	--2857
		x"38",	--2858
		x"46",	--2859
		x"00",	--2860
		x"47",	--2861
		x"00",	--2862
		x"49",	--2863
		x"f0",	--2864
		x"00",	--2865
		x"24",	--2866
		x"46",	--2867
		x"47",	--2868
		x"c3",	--2869
		x"10",	--2870
		x"10",	--2871
		x"53",	--2872
		x"23",	--2873
		x"4a",	--2874
		x"00",	--2875
		x"4b",	--2876
		x"00",	--2877
		x"43",	--2878
		x"43",	--2879
		x"f0",	--2880
		x"00",	--2881
		x"24",	--2882
		x"5c",	--2883
		x"6d",	--2884
		x"53",	--2885
		x"23",	--2886
		x"53",	--2887
		x"63",	--2888
		x"f6",	--2889
		x"f7",	--2890
		x"43",	--2891
		x"43",	--2892
		x"93",	--2893
		x"20",	--2894
		x"93",	--2895
		x"24",	--2896
		x"41",	--2897
		x"00",	--2898
		x"41",	--2899
		x"00",	--2900
		x"da",	--2901
		x"db",	--2902
		x"4f",	--2903
		x"00",	--2904
		x"9e",	--2905
		x"00",	--2906
		x"20",	--2907
		x"4f",	--2908
		x"00",	--2909
		x"41",	--2910
		x"00",	--2911
		x"46",	--2912
		x"47",	--2913
		x"54",	--2914
		x"65",	--2915
		x"4e",	--2916
		x"00",	--2917
		x"4f",	--2918
		x"00",	--2919
		x"40",	--2920
		x"00",	--2921
		x"00",	--2922
		x"93",	--2923
		x"38",	--2924
		x"48",	--2925
		x"50",	--2926
		x"00",	--2927
		x"41",	--2928
		x"41",	--2929
		x"41",	--2930
		x"41",	--2931
		x"41",	--2932
		x"41",	--2933
		x"41",	--2934
		x"41",	--2935
		x"41",	--2936
		x"91",	--2937
		x"38",	--2938
		x"4b",	--2939
		x"00",	--2940
		x"43",	--2941
		x"43",	--2942
		x"4f",	--2943
		x"00",	--2944
		x"9e",	--2945
		x"00",	--2946
		x"27",	--2947
		x"93",	--2948
		x"24",	--2949
		x"46",	--2950
		x"47",	--2951
		x"84",	--2952
		x"75",	--2953
		x"93",	--2954
		x"38",	--2955
		x"43",	--2956
		x"00",	--2957
		x"41",	--2958
		x"00",	--2959
		x"4e",	--2960
		x"00",	--2961
		x"4f",	--2962
		x"00",	--2963
		x"4e",	--2964
		x"4f",	--2965
		x"53",	--2966
		x"63",	--2967
		x"90",	--2968
		x"3f",	--2969
		x"28",	--2970
		x"90",	--2971
		x"40",	--2972
		x"2c",	--2973
		x"93",	--2974
		x"2c",	--2975
		x"48",	--2976
		x"00",	--2977
		x"53",	--2978
		x"5e",	--2979
		x"6f",	--2980
		x"4b",	--2981
		x"53",	--2982
		x"4e",	--2983
		x"4f",	--2984
		x"53",	--2985
		x"63",	--2986
		x"90",	--2987
		x"3f",	--2988
		x"2b",	--2989
		x"24",	--2990
		x"4e",	--2991
		x"00",	--2992
		x"4f",	--2993
		x"00",	--2994
		x"4a",	--2995
		x"00",	--2996
		x"40",	--2997
		x"00",	--2998
		x"00",	--2999
		x"93",	--3000
		x"37",	--3001
		x"4e",	--3002
		x"4f",	--3003
		x"f3",	--3004
		x"f3",	--3005
		x"c3",	--3006
		x"10",	--3007
		x"10",	--3008
		x"4c",	--3009
		x"4d",	--3010
		x"de",	--3011
		x"df",	--3012
		x"4a",	--3013
		x"00",	--3014
		x"4b",	--3015
		x"00",	--3016
		x"53",	--3017
		x"00",	--3018
		x"48",	--3019
		x"3f",	--3020
		x"93",	--3021
		x"23",	--3022
		x"4f",	--3023
		x"00",	--3024
		x"4f",	--3025
		x"00",	--3026
		x"00",	--3027
		x"4f",	--3028
		x"00",	--3029
		x"00",	--3030
		x"4f",	--3031
		x"00",	--3032
		x"00",	--3033
		x"4e",	--3034
		x"00",	--3035
		x"ff",	--3036
		x"00",	--3037
		x"4e",	--3038
		x"00",	--3039
		x"4d",	--3040
		x"3f",	--3041
		x"43",	--3042
		x"43",	--3043
		x"3f",	--3044
		x"e3",	--3045
		x"53",	--3046
		x"90",	--3047
		x"00",	--3048
		x"37",	--3049
		x"3f",	--3050
		x"93",	--3051
		x"2b",	--3052
		x"3f",	--3053
		x"44",	--3054
		x"45",	--3055
		x"86",	--3056
		x"77",	--3057
		x"3f",	--3058
		x"4e",	--3059
		x"3f",	--3060
		x"43",	--3061
		x"00",	--3062
		x"41",	--3063
		x"00",	--3064
		x"e3",	--3065
		x"e3",	--3066
		x"53",	--3067
		x"63",	--3068
		x"4e",	--3069
		x"00",	--3070
		x"4f",	--3071
		x"00",	--3072
		x"3f",	--3073
		x"93",	--3074
		x"27",	--3075
		x"59",	--3076
		x"00",	--3077
		x"44",	--3078
		x"00",	--3079
		x"45",	--3080
		x"00",	--3081
		x"49",	--3082
		x"f0",	--3083
		x"00",	--3084
		x"24",	--3085
		x"4d",	--3086
		x"44",	--3087
		x"45",	--3088
		x"c3",	--3089
		x"10",	--3090
		x"10",	--3091
		x"53",	--3092
		x"23",	--3093
		x"4c",	--3094
		x"00",	--3095
		x"4d",	--3096
		x"00",	--3097
		x"43",	--3098
		x"43",	--3099
		x"f0",	--3100
		x"00",	--3101
		x"24",	--3102
		x"5c",	--3103
		x"6d",	--3104
		x"53",	--3105
		x"23",	--3106
		x"53",	--3107
		x"63",	--3108
		x"f4",	--3109
		x"f5",	--3110
		x"43",	--3111
		x"43",	--3112
		x"93",	--3113
		x"20",	--3114
		x"93",	--3115
		x"20",	--3116
		x"43",	--3117
		x"43",	--3118
		x"41",	--3119
		x"00",	--3120
		x"41",	--3121
		x"00",	--3122
		x"da",	--3123
		x"db",	--3124
		x"3f",	--3125
		x"43",	--3126
		x"43",	--3127
		x"3f",	--3128
		x"92",	--3129
		x"23",	--3130
		x"9e",	--3131
		x"00",	--3132
		x"00",	--3133
		x"27",	--3134
		x"40",	--3135
		x"f1",	--3136
		x"3f",	--3137
		x"50",	--3138
		x"ff",	--3139
		x"4e",	--3140
		x"00",	--3141
		x"4f",	--3142
		x"00",	--3143
		x"4c",	--3144
		x"00",	--3145
		x"4d",	--3146
		x"00",	--3147
		x"41",	--3148
		x"50",	--3149
		x"00",	--3150
		x"41",	--3151
		x"52",	--3152
		x"12",	--3153
		x"e1",	--3154
		x"41",	--3155
		x"50",	--3156
		x"00",	--3157
		x"41",	--3158
		x"12",	--3159
		x"e1",	--3160
		x"41",	--3161
		x"52",	--3162
		x"41",	--3163
		x"50",	--3164
		x"00",	--3165
		x"41",	--3166
		x"50",	--3167
		x"00",	--3168
		x"12",	--3169
		x"d5",	--3170
		x"12",	--3171
		x"e0",	--3172
		x"50",	--3173
		x"00",	--3174
		x"41",	--3175
		x"50",	--3176
		x"ff",	--3177
		x"4e",	--3178
		x"00",	--3179
		x"4f",	--3180
		x"00",	--3181
		x"4c",	--3182
		x"00",	--3183
		x"4d",	--3184
		x"00",	--3185
		x"41",	--3186
		x"50",	--3187
		x"00",	--3188
		x"41",	--3189
		x"52",	--3190
		x"12",	--3191
		x"e1",	--3192
		x"41",	--3193
		x"50",	--3194
		x"00",	--3195
		x"41",	--3196
		x"12",	--3197
		x"e1",	--3198
		x"e3",	--3199
		x"00",	--3200
		x"41",	--3201
		x"52",	--3202
		x"41",	--3203
		x"50",	--3204
		x"00",	--3205
		x"41",	--3206
		x"50",	--3207
		x"00",	--3208
		x"12",	--3209
		x"d5",	--3210
		x"12",	--3211
		x"e0",	--3212
		x"50",	--3213
		x"00",	--3214
		x"41",	--3215
		x"12",	--3216
		x"12",	--3217
		x"12",	--3218
		x"12",	--3219
		x"12",	--3220
		x"12",	--3221
		x"12",	--3222
		x"12",	--3223
		x"50",	--3224
		x"ff",	--3225
		x"4e",	--3226
		x"00",	--3227
		x"4f",	--3228
		x"00",	--3229
		x"4c",	--3230
		x"00",	--3231
		x"4d",	--3232
		x"00",	--3233
		x"41",	--3234
		x"50",	--3235
		x"00",	--3236
		x"41",	--3237
		x"52",	--3238
		x"12",	--3239
		x"e1",	--3240
		x"41",	--3241
		x"50",	--3242
		x"00",	--3243
		x"41",	--3244
		x"12",	--3245
		x"e1",	--3246
		x"41",	--3247
		x"00",	--3248
		x"93",	--3249
		x"28",	--3250
		x"41",	--3251
		x"00",	--3252
		x"93",	--3253
		x"28",	--3254
		x"92",	--3255
		x"24",	--3256
		x"92",	--3257
		x"24",	--3258
		x"93",	--3259
		x"24",	--3260
		x"93",	--3261
		x"24",	--3262
		x"41",	--3263
		x"00",	--3264
		x"41",	--3265
		x"00",	--3266
		x"41",	--3267
		x"00",	--3268
		x"41",	--3269
		x"00",	--3270
		x"40",	--3271
		x"00",	--3272
		x"43",	--3273
		x"43",	--3274
		x"43",	--3275
		x"43",	--3276
		x"43",	--3277
		x"00",	--3278
		x"43",	--3279
		x"00",	--3280
		x"43",	--3281
		x"43",	--3282
		x"4c",	--3283
		x"00",	--3284
		x"3c",	--3285
		x"58",	--3286
		x"69",	--3287
		x"c3",	--3288
		x"10",	--3289
		x"10",	--3290
		x"53",	--3291
		x"00",	--3292
		x"24",	--3293
		x"b3",	--3294
		x"24",	--3295
		x"58",	--3296
		x"69",	--3297
		x"56",	--3298
		x"67",	--3299
		x"43",	--3300
		x"43",	--3301
		x"99",	--3302
		x"28",	--3303
		x"24",	--3304
		x"43",	--3305
		x"43",	--3306
		x"5c",	--3307
		x"6d",	--3308
		x"56",	--3309
		x"67",	--3310
		x"93",	--3311
		x"37",	--3312
		x"d3",	--3313
		x"d3",	--3314
		x"3f",	--3315
		x"98",	--3316
		x"2b",	--3317
		x"3f",	--3318
		x"4a",	--3319
		x"00",	--3320
		x"4b",	--3321
		x"00",	--3322
		x"4f",	--3323
		x"41",	--3324
		x"00",	--3325
		x"51",	--3326
		x"00",	--3327
		x"4a",	--3328
		x"53",	--3329
		x"46",	--3330
		x"00",	--3331
		x"43",	--3332
		x"91",	--3333
		x"00",	--3334
		x"00",	--3335
		x"24",	--3336
		x"4d",	--3337
		x"00",	--3338
		x"93",	--3339
		x"38",	--3340
		x"90",	--3341
		x"40",	--3342
		x"2c",	--3343
		x"41",	--3344
		x"00",	--3345
		x"53",	--3346
		x"41",	--3347
		x"00",	--3348
		x"41",	--3349
		x"00",	--3350
		x"4d",	--3351
		x"5e",	--3352
		x"6f",	--3353
		x"93",	--3354
		x"38",	--3355
		x"5a",	--3356
		x"6b",	--3357
		x"53",	--3358
		x"90",	--3359
		x"40",	--3360
		x"2b",	--3361
		x"4a",	--3362
		x"00",	--3363
		x"4b",	--3364
		x"00",	--3365
		x"4c",	--3366
		x"00",	--3367
		x"4e",	--3368
		x"4f",	--3369
		x"f0",	--3370
		x"00",	--3371
		x"f3",	--3372
		x"90",	--3373
		x"00",	--3374
		x"24",	--3375
		x"4e",	--3376
		x"00",	--3377
		x"4f",	--3378
		x"00",	--3379
		x"40",	--3380
		x"00",	--3381
		x"00",	--3382
		x"41",	--3383
		x"52",	--3384
		x"12",	--3385
		x"e0",	--3386
		x"50",	--3387
		x"00",	--3388
		x"41",	--3389
		x"41",	--3390
		x"41",	--3391
		x"41",	--3392
		x"41",	--3393
		x"41",	--3394
		x"41",	--3395
		x"41",	--3396
		x"41",	--3397
		x"d3",	--3398
		x"d3",	--3399
		x"3f",	--3400
		x"50",	--3401
		x"00",	--3402
		x"4a",	--3403
		x"b3",	--3404
		x"24",	--3405
		x"41",	--3406
		x"00",	--3407
		x"41",	--3408
		x"00",	--3409
		x"c3",	--3410
		x"10",	--3411
		x"10",	--3412
		x"4c",	--3413
		x"4d",	--3414
		x"d3",	--3415
		x"d0",	--3416
		x"80",	--3417
		x"46",	--3418
		x"00",	--3419
		x"47",	--3420
		x"00",	--3421
		x"c3",	--3422
		x"10",	--3423
		x"10",	--3424
		x"53",	--3425
		x"93",	--3426
		x"3b",	--3427
		x"48",	--3428
		x"00",	--3429
		x"3f",	--3430
		x"93",	--3431
		x"24",	--3432
		x"43",	--3433
		x"91",	--3434
		x"00",	--3435
		x"00",	--3436
		x"24",	--3437
		x"4f",	--3438
		x"00",	--3439
		x"41",	--3440
		x"50",	--3441
		x"00",	--3442
		x"3f",	--3443
		x"93",	--3444
		x"23",	--3445
		x"4e",	--3446
		x"4f",	--3447
		x"f0",	--3448
		x"00",	--3449
		x"f3",	--3450
		x"93",	--3451
		x"23",	--3452
		x"93",	--3453
		x"23",	--3454
		x"93",	--3455
		x"00",	--3456
		x"20",	--3457
		x"93",	--3458
		x"00",	--3459
		x"27",	--3460
		x"50",	--3461
		x"00",	--3462
		x"63",	--3463
		x"f0",	--3464
		x"ff",	--3465
		x"f3",	--3466
		x"3f",	--3467
		x"43",	--3468
		x"3f",	--3469
		x"43",	--3470
		x"3f",	--3471
		x"43",	--3472
		x"91",	--3473
		x"00",	--3474
		x"00",	--3475
		x"24",	--3476
		x"4f",	--3477
		x"00",	--3478
		x"41",	--3479
		x"50",	--3480
		x"00",	--3481
		x"3f",	--3482
		x"43",	--3483
		x"3f",	--3484
		x"93",	--3485
		x"23",	--3486
		x"40",	--3487
		x"f1",	--3488
		x"3f",	--3489
		x"12",	--3490
		x"12",	--3491
		x"12",	--3492
		x"12",	--3493
		x"12",	--3494
		x"50",	--3495
		x"ff",	--3496
		x"4e",	--3497
		x"00",	--3498
		x"4f",	--3499
		x"00",	--3500
		x"4c",	--3501
		x"00",	--3502
		x"4d",	--3503
		x"00",	--3504
		x"41",	--3505
		x"50",	--3506
		x"00",	--3507
		x"41",	--3508
		x"52",	--3509
		x"12",	--3510
		x"e1",	--3511
		x"41",	--3512
		x"52",	--3513
		x"41",	--3514
		x"12",	--3515
		x"e1",	--3516
		x"41",	--3517
		x"00",	--3518
		x"93",	--3519
		x"28",	--3520
		x"41",	--3521
		x"00",	--3522
		x"93",	--3523
		x"28",	--3524
		x"e1",	--3525
		x"00",	--3526
		x"00",	--3527
		x"92",	--3528
		x"24",	--3529
		x"93",	--3530
		x"24",	--3531
		x"92",	--3532
		x"24",	--3533
		x"93",	--3534
		x"24",	--3535
		x"41",	--3536
		x"00",	--3537
		x"81",	--3538
		x"00",	--3539
		x"4d",	--3540
		x"00",	--3541
		x"41",	--3542
		x"00",	--3543
		x"41",	--3544
		x"00",	--3545
		x"41",	--3546
		x"00",	--3547
		x"41",	--3548
		x"00",	--3549
		x"99",	--3550
		x"2c",	--3551
		x"5e",	--3552
		x"6f",	--3553
		x"53",	--3554
		x"4d",	--3555
		x"00",	--3556
		x"40",	--3557
		x"00",	--3558
		x"43",	--3559
		x"40",	--3560
		x"40",	--3561
		x"43",	--3562
		x"43",	--3563
		x"3c",	--3564
		x"dc",	--3565
		x"dd",	--3566
		x"88",	--3567
		x"79",	--3568
		x"c3",	--3569
		x"10",	--3570
		x"10",	--3571
		x"5e",	--3572
		x"6f",	--3573
		x"53",	--3574
		x"24",	--3575
		x"99",	--3576
		x"2b",	--3577
		x"23",	--3578
		x"98",	--3579
		x"2b",	--3580
		x"3f",	--3581
		x"9f",	--3582
		x"2b",	--3583
		x"98",	--3584
		x"2f",	--3585
		x"3f",	--3586
		x"4a",	--3587
		x"4b",	--3588
		x"f0",	--3589
		x"00",	--3590
		x"f3",	--3591
		x"90",	--3592
		x"00",	--3593
		x"24",	--3594
		x"4a",	--3595
		x"00",	--3596
		x"4b",	--3597
		x"00",	--3598
		x"41",	--3599
		x"50",	--3600
		x"00",	--3601
		x"12",	--3602
		x"e0",	--3603
		x"50",	--3604
		x"00",	--3605
		x"41",	--3606
		x"41",	--3607
		x"41",	--3608
		x"41",	--3609
		x"41",	--3610
		x"41",	--3611
		x"42",	--3612
		x"00",	--3613
		x"41",	--3614
		x"50",	--3615
		x"00",	--3616
		x"3f",	--3617
		x"9e",	--3618
		x"23",	--3619
		x"40",	--3620
		x"f1",	--3621
		x"3f",	--3622
		x"93",	--3623
		x"23",	--3624
		x"4a",	--3625
		x"4b",	--3626
		x"f0",	--3627
		x"00",	--3628
		x"f3",	--3629
		x"93",	--3630
		x"23",	--3631
		x"93",	--3632
		x"23",	--3633
		x"93",	--3634
		x"20",	--3635
		x"93",	--3636
		x"27",	--3637
		x"50",	--3638
		x"00",	--3639
		x"63",	--3640
		x"f0",	--3641
		x"ff",	--3642
		x"f3",	--3643
		x"3f",	--3644
		x"43",	--3645
		x"00",	--3646
		x"43",	--3647
		x"00",	--3648
		x"43",	--3649
		x"00",	--3650
		x"41",	--3651
		x"50",	--3652
		x"00",	--3653
		x"3f",	--3654
		x"41",	--3655
		x"52",	--3656
		x"3f",	--3657
		x"50",	--3658
		x"ff",	--3659
		x"4e",	--3660
		x"00",	--3661
		x"4f",	--3662
		x"00",	--3663
		x"4c",	--3664
		x"00",	--3665
		x"4d",	--3666
		x"00",	--3667
		x"41",	--3668
		x"50",	--3669
		x"00",	--3670
		x"41",	--3671
		x"52",	--3672
		x"12",	--3673
		x"e1",	--3674
		x"41",	--3675
		x"52",	--3676
		x"41",	--3677
		x"12",	--3678
		x"e1",	--3679
		x"93",	--3680
		x"00",	--3681
		x"28",	--3682
		x"93",	--3683
		x"00",	--3684
		x"28",	--3685
		x"41",	--3686
		x"52",	--3687
		x"41",	--3688
		x"50",	--3689
		x"00",	--3690
		x"12",	--3691
		x"e3",	--3692
		x"50",	--3693
		x"00",	--3694
		x"41",	--3695
		x"43",	--3696
		x"3f",	--3697
		x"50",	--3698
		x"ff",	--3699
		x"4e",	--3700
		x"00",	--3701
		x"4f",	--3702
		x"00",	--3703
		x"4c",	--3704
		x"00",	--3705
		x"4d",	--3706
		x"00",	--3707
		x"41",	--3708
		x"50",	--3709
		x"00",	--3710
		x"41",	--3711
		x"52",	--3712
		x"12",	--3713
		x"e1",	--3714
		x"41",	--3715
		x"52",	--3716
		x"41",	--3717
		x"12",	--3718
		x"e1",	--3719
		x"93",	--3720
		x"00",	--3721
		x"28",	--3722
		x"93",	--3723
		x"00",	--3724
		x"28",	--3725
		x"41",	--3726
		x"52",	--3727
		x"41",	--3728
		x"50",	--3729
		x"00",	--3730
		x"12",	--3731
		x"e3",	--3732
		x"50",	--3733
		x"00",	--3734
		x"41",	--3735
		x"43",	--3736
		x"3f",	--3737
		x"50",	--3738
		x"ff",	--3739
		x"4e",	--3740
		x"00",	--3741
		x"4f",	--3742
		x"00",	--3743
		x"4c",	--3744
		x"00",	--3745
		x"4d",	--3746
		x"00",	--3747
		x"41",	--3748
		x"50",	--3749
		x"00",	--3750
		x"41",	--3751
		x"52",	--3752
		x"12",	--3753
		x"e1",	--3754
		x"41",	--3755
		x"52",	--3756
		x"41",	--3757
		x"12",	--3758
		x"e1",	--3759
		x"93",	--3760
		x"00",	--3761
		x"28",	--3762
		x"93",	--3763
		x"00",	--3764
		x"28",	--3765
		x"41",	--3766
		x"52",	--3767
		x"41",	--3768
		x"50",	--3769
		x"00",	--3770
		x"12",	--3771
		x"e3",	--3772
		x"50",	--3773
		x"00",	--3774
		x"41",	--3775
		x"43",	--3776
		x"3f",	--3777
		x"12",	--3778
		x"12",	--3779
		x"82",	--3780
		x"40",	--3781
		x"00",	--3782
		x"00",	--3783
		x"4f",	--3784
		x"5d",	--3785
		x"43",	--3786
		x"6d",	--3787
		x"4d",	--3788
		x"4d",	--3789
		x"00",	--3790
		x"93",	--3791
		x"20",	--3792
		x"93",	--3793
		x"20",	--3794
		x"43",	--3795
		x"00",	--3796
		x"41",	--3797
		x"12",	--3798
		x"e0",	--3799
		x"52",	--3800
		x"41",	--3801
		x"41",	--3802
		x"41",	--3803
		x"40",	--3804
		x"00",	--3805
		x"00",	--3806
		x"93",	--3807
		x"20",	--3808
		x"4e",	--3809
		x"4f",	--3810
		x"4a",	--3811
		x"00",	--3812
		x"4b",	--3813
		x"00",	--3814
		x"4a",	--3815
		x"4b",	--3816
		x"12",	--3817
		x"df",	--3818
		x"53",	--3819
		x"93",	--3820
		x"3b",	--3821
		x"4a",	--3822
		x"00",	--3823
		x"4b",	--3824
		x"00",	--3825
		x"4f",	--3826
		x"f0",	--3827
		x"00",	--3828
		x"20",	--3829
		x"40",	--3830
		x"00",	--3831
		x"8f",	--3832
		x"4e",	--3833
		x"00",	--3834
		x"3f",	--3835
		x"93",	--3836
		x"24",	--3837
		x"4e",	--3838
		x"4f",	--3839
		x"e3",	--3840
		x"e3",	--3841
		x"53",	--3842
		x"63",	--3843
		x"3f",	--3844
		x"51",	--3845
		x"00",	--3846
		x"00",	--3847
		x"61",	--3848
		x"00",	--3849
		x"00",	--3850
		x"53",	--3851
		x"23",	--3852
		x"3f",	--3853
		x"90",	--3854
		x"80",	--3855
		x"23",	--3856
		x"43",	--3857
		x"40",	--3858
		x"cf",	--3859
		x"3f",	--3860
		x"50",	--3861
		x"ff",	--3862
		x"4e",	--3863
		x"00",	--3864
		x"4f",	--3865
		x"00",	--3866
		x"41",	--3867
		x"52",	--3868
		x"41",	--3869
		x"12",	--3870
		x"e1",	--3871
		x"41",	--3872
		x"00",	--3873
		x"93",	--3874
		x"24",	--3875
		x"28",	--3876
		x"92",	--3877
		x"24",	--3878
		x"41",	--3879
		x"00",	--3880
		x"93",	--3881
		x"38",	--3882
		x"90",	--3883
		x"00",	--3884
		x"38",	--3885
		x"93",	--3886
		x"00",	--3887
		x"20",	--3888
		x"43",	--3889
		x"40",	--3890
		x"7f",	--3891
		x"50",	--3892
		x"00",	--3893
		x"41",	--3894
		x"41",	--3895
		x"00",	--3896
		x"41",	--3897
		x"00",	--3898
		x"40",	--3899
		x"00",	--3900
		x"8d",	--3901
		x"4c",	--3902
		x"f0",	--3903
		x"00",	--3904
		x"20",	--3905
		x"93",	--3906
		x"00",	--3907
		x"27",	--3908
		x"e3",	--3909
		x"e3",	--3910
		x"53",	--3911
		x"63",	--3912
		x"50",	--3913
		x"00",	--3914
		x"41",	--3915
		x"43",	--3916
		x"43",	--3917
		x"50",	--3918
		x"00",	--3919
		x"41",	--3920
		x"c3",	--3921
		x"10",	--3922
		x"10",	--3923
		x"53",	--3924
		x"23",	--3925
		x"3f",	--3926
		x"43",	--3927
		x"40",	--3928
		x"80",	--3929
		x"50",	--3930
		x"00",	--3931
		x"41",	--3932
		x"12",	--3933
		x"12",	--3934
		x"12",	--3935
		x"12",	--3936
		x"82",	--3937
		x"4e",	--3938
		x"4f",	--3939
		x"43",	--3940
		x"00",	--3941
		x"93",	--3942
		x"20",	--3943
		x"93",	--3944
		x"20",	--3945
		x"43",	--3946
		x"00",	--3947
		x"41",	--3948
		x"12",	--3949
		x"e0",	--3950
		x"52",	--3951
		x"41",	--3952
		x"41",	--3953
		x"41",	--3954
		x"41",	--3955
		x"41",	--3956
		x"40",	--3957
		x"00",	--3958
		x"00",	--3959
		x"40",	--3960
		x"00",	--3961
		x"00",	--3962
		x"4a",	--3963
		x"00",	--3964
		x"4b",	--3965
		x"00",	--3966
		x"4a",	--3967
		x"4b",	--3968
		x"12",	--3969
		x"df",	--3970
		x"53",	--3971
		x"93",	--3972
		x"38",	--3973
		x"27",	--3974
		x"4a",	--3975
		x"00",	--3976
		x"4b",	--3977
		x"00",	--3978
		x"4f",	--3979
		x"f0",	--3980
		x"00",	--3981
		x"20",	--3982
		x"40",	--3983
		x"00",	--3984
		x"8f",	--3985
		x"4e",	--3986
		x"00",	--3987
		x"3f",	--3988
		x"51",	--3989
		x"00",	--3990
		x"00",	--3991
		x"61",	--3992
		x"00",	--3993
		x"00",	--3994
		x"53",	--3995
		x"23",	--3996
		x"3f",	--3997
		x"4f",	--3998
		x"e3",	--3999
		x"53",	--4000
		x"43",	--4001
		x"43",	--4002
		x"4e",	--4003
		x"f0",	--4004
		x"00",	--4005
		x"24",	--4006
		x"5c",	--4007
		x"6d",	--4008
		x"53",	--4009
		x"23",	--4010
		x"53",	--4011
		x"63",	--4012
		x"fa",	--4013
		x"fb",	--4014
		x"43",	--4015
		x"43",	--4016
		x"93",	--4017
		x"20",	--4018
		x"93",	--4019
		x"20",	--4020
		x"43",	--4021
		x"43",	--4022
		x"f0",	--4023
		x"00",	--4024
		x"20",	--4025
		x"48",	--4026
		x"49",	--4027
		x"da",	--4028
		x"db",	--4029
		x"4d",	--4030
		x"00",	--4031
		x"4e",	--4032
		x"00",	--4033
		x"40",	--4034
		x"00",	--4035
		x"8f",	--4036
		x"4e",	--4037
		x"00",	--4038
		x"3f",	--4039
		x"c3",	--4040
		x"10",	--4041
		x"10",	--4042
		x"53",	--4043
		x"23",	--4044
		x"3f",	--4045
		x"12",	--4046
		x"12",	--4047
		x"12",	--4048
		x"93",	--4049
		x"2c",	--4050
		x"90",	--4051
		x"01",	--4052
		x"28",	--4053
		x"40",	--4054
		x"00",	--4055
		x"43",	--4056
		x"42",	--4057
		x"4e",	--4058
		x"4f",	--4059
		x"49",	--4060
		x"93",	--4061
		x"20",	--4062
		x"50",	--4063
		x"f1",	--4064
		x"4c",	--4065
		x"43",	--4066
		x"8e",	--4067
		x"7f",	--4068
		x"4a",	--4069
		x"41",	--4070
		x"41",	--4071
		x"41",	--4072
		x"41",	--4073
		x"90",	--4074
		x"01",	--4075
		x"28",	--4076
		x"42",	--4077
		x"43",	--4078
		x"40",	--4079
		x"00",	--4080
		x"4e",	--4081
		x"4f",	--4082
		x"49",	--4083
		x"93",	--4084
		x"27",	--4085
		x"c3",	--4086
		x"10",	--4087
		x"10",	--4088
		x"53",	--4089
		x"23",	--4090
		x"3f",	--4091
		x"40",	--4092
		x"00",	--4093
		x"43",	--4094
		x"40",	--4095
		x"00",	--4096
		x"3f",	--4097
		x"40",	--4098
		x"00",	--4099
		x"43",	--4100
		x"43",	--4101
		x"3f",	--4102
		x"12",	--4103
		x"12",	--4104
		x"12",	--4105
		x"12",	--4106
		x"12",	--4107
		x"4f",	--4108
		x"4f",	--4109
		x"00",	--4110
		x"4f",	--4111
		x"00",	--4112
		x"4d",	--4113
		x"00",	--4114
		x"4d",	--4115
		x"93",	--4116
		x"28",	--4117
		x"92",	--4118
		x"24",	--4119
		x"93",	--4120
		x"24",	--4121
		x"93",	--4122
		x"24",	--4123
		x"4d",	--4124
		x"00",	--4125
		x"90",	--4126
		x"ff",	--4127
		x"38",	--4128
		x"90",	--4129
		x"00",	--4130
		x"34",	--4131
		x"4e",	--4132
		x"4f",	--4133
		x"f0",	--4134
		x"00",	--4135
		x"f3",	--4136
		x"90",	--4137
		x"00",	--4138
		x"24",	--4139
		x"50",	--4140
		x"00",	--4141
		x"63",	--4142
		x"93",	--4143
		x"38",	--4144
		x"4b",	--4145
		x"50",	--4146
		x"00",	--4147
		x"c3",	--4148
		x"10",	--4149
		x"10",	--4150
		x"c3",	--4151
		x"10",	--4152
		x"10",	--4153
		x"c3",	--4154
		x"10",	--4155
		x"10",	--4156
		x"c3",	--4157
		x"10",	--4158
		x"10",	--4159
		x"c3",	--4160
		x"10",	--4161
		x"10",	--4162
		x"c3",	--4163
		x"10",	--4164
		x"10",	--4165
		x"c3",	--4166
		x"10",	--4167
		x"10",	--4168
		x"f3",	--4169
		x"f0",	--4170
		x"00",	--4171
		x"4d",	--4172
		x"3c",	--4173
		x"93",	--4174
		x"23",	--4175
		x"43",	--4176
		x"43",	--4177
		x"43",	--4178
		x"4d",	--4179
		x"5d",	--4180
		x"5d",	--4181
		x"5d",	--4182
		x"5d",	--4183
		x"5d",	--4184
		x"5d",	--4185
		x"5d",	--4186
		x"4f",	--4187
		x"f0",	--4188
		x"00",	--4189
		x"dd",	--4190
		x"4a",	--4191
		x"11",	--4192
		x"43",	--4193
		x"10",	--4194
		x"4c",	--4195
		x"df",	--4196
		x"4d",	--4197
		x"41",	--4198
		x"41",	--4199
		x"41",	--4200
		x"41",	--4201
		x"41",	--4202
		x"41",	--4203
		x"93",	--4204
		x"23",	--4205
		x"4e",	--4206
		x"4f",	--4207
		x"f0",	--4208
		x"00",	--4209
		x"f3",	--4210
		x"93",	--4211
		x"20",	--4212
		x"93",	--4213
		x"27",	--4214
		x"50",	--4215
		x"00",	--4216
		x"63",	--4217
		x"3f",	--4218
		x"c3",	--4219
		x"10",	--4220
		x"10",	--4221
		x"4b",	--4222
		x"50",	--4223
		x"00",	--4224
		x"3f",	--4225
		x"43",	--4226
		x"43",	--4227
		x"43",	--4228
		x"3f",	--4229
		x"d3",	--4230
		x"d0",	--4231
		x"00",	--4232
		x"f3",	--4233
		x"f0",	--4234
		x"00",	--4235
		x"43",	--4236
		x"3f",	--4237
		x"40",	--4238
		x"ff",	--4239
		x"8b",	--4240
		x"90",	--4241
		x"00",	--4242
		x"34",	--4243
		x"4e",	--4244
		x"4f",	--4245
		x"47",	--4246
		x"f0",	--4247
		x"00",	--4248
		x"24",	--4249
		x"c3",	--4250
		x"10",	--4251
		x"10",	--4252
		x"53",	--4253
		x"23",	--4254
		x"43",	--4255
		x"43",	--4256
		x"f0",	--4257
		x"00",	--4258
		x"24",	--4259
		x"58",	--4260
		x"69",	--4261
		x"53",	--4262
		x"23",	--4263
		x"53",	--4264
		x"63",	--4265
		x"fe",	--4266
		x"ff",	--4267
		x"43",	--4268
		x"43",	--4269
		x"93",	--4270
		x"20",	--4271
		x"93",	--4272
		x"20",	--4273
		x"43",	--4274
		x"43",	--4275
		x"4e",	--4276
		x"4f",	--4277
		x"dc",	--4278
		x"dd",	--4279
		x"48",	--4280
		x"49",	--4281
		x"f0",	--4282
		x"00",	--4283
		x"f3",	--4284
		x"90",	--4285
		x"00",	--4286
		x"24",	--4287
		x"50",	--4288
		x"00",	--4289
		x"63",	--4290
		x"48",	--4291
		x"49",	--4292
		x"c3",	--4293
		x"10",	--4294
		x"10",	--4295
		x"c3",	--4296
		x"10",	--4297
		x"10",	--4298
		x"c3",	--4299
		x"10",	--4300
		x"10",	--4301
		x"c3",	--4302
		x"10",	--4303
		x"10",	--4304
		x"c3",	--4305
		x"10",	--4306
		x"10",	--4307
		x"c3",	--4308
		x"10",	--4309
		x"10",	--4310
		x"c3",	--4311
		x"10",	--4312
		x"10",	--4313
		x"f3",	--4314
		x"f0",	--4315
		x"00",	--4316
		x"43",	--4317
		x"90",	--4318
		x"40",	--4319
		x"2f",	--4320
		x"43",	--4321
		x"3f",	--4322
		x"43",	--4323
		x"43",	--4324
		x"3f",	--4325
		x"93",	--4326
		x"23",	--4327
		x"48",	--4328
		x"49",	--4329
		x"f0",	--4330
		x"00",	--4331
		x"f3",	--4332
		x"93",	--4333
		x"24",	--4334
		x"50",	--4335
		x"00",	--4336
		x"63",	--4337
		x"3f",	--4338
		x"93",	--4339
		x"27",	--4340
		x"3f",	--4341
		x"12",	--4342
		x"12",	--4343
		x"4f",	--4344
		x"4f",	--4345
		x"00",	--4346
		x"f0",	--4347
		x"00",	--4348
		x"4f",	--4349
		x"00",	--4350
		x"c3",	--4351
		x"10",	--4352
		x"c3",	--4353
		x"10",	--4354
		x"c3",	--4355
		x"10",	--4356
		x"c3",	--4357
		x"10",	--4358
		x"c3",	--4359
		x"10",	--4360
		x"c3",	--4361
		x"10",	--4362
		x"c3",	--4363
		x"10",	--4364
		x"4d",	--4365
		x"4f",	--4366
		x"00",	--4367
		x"b0",	--4368
		x"00",	--4369
		x"43",	--4370
		x"6f",	--4371
		x"4f",	--4372
		x"00",	--4373
		x"93",	--4374
		x"20",	--4375
		x"93",	--4376
		x"24",	--4377
		x"40",	--4378
		x"ff",	--4379
		x"00",	--4380
		x"4a",	--4381
		x"4b",	--4382
		x"5c",	--4383
		x"6d",	--4384
		x"5c",	--4385
		x"6d",	--4386
		x"5c",	--4387
		x"6d",	--4388
		x"5c",	--4389
		x"6d",	--4390
		x"5c",	--4391
		x"6d",	--4392
		x"5c",	--4393
		x"6d",	--4394
		x"5c",	--4395
		x"6d",	--4396
		x"40",	--4397
		x"00",	--4398
		x"00",	--4399
		x"90",	--4400
		x"40",	--4401
		x"2c",	--4402
		x"40",	--4403
		x"ff",	--4404
		x"5c",	--4405
		x"6d",	--4406
		x"4f",	--4407
		x"53",	--4408
		x"90",	--4409
		x"40",	--4410
		x"2b",	--4411
		x"4a",	--4412
		x"00",	--4413
		x"4c",	--4414
		x"00",	--4415
		x"4d",	--4416
		x"00",	--4417
		x"41",	--4418
		x"41",	--4419
		x"41",	--4420
		x"90",	--4421
		x"00",	--4422
		x"24",	--4423
		x"50",	--4424
		x"ff",	--4425
		x"4d",	--4426
		x"00",	--4427
		x"40",	--4428
		x"00",	--4429
		x"00",	--4430
		x"4a",	--4431
		x"4b",	--4432
		x"5c",	--4433
		x"6d",	--4434
		x"5c",	--4435
		x"6d",	--4436
		x"5c",	--4437
		x"6d",	--4438
		x"5c",	--4439
		x"6d",	--4440
		x"5c",	--4441
		x"6d",	--4442
		x"5c",	--4443
		x"6d",	--4444
		x"5c",	--4445
		x"6d",	--4446
		x"4c",	--4447
		x"4d",	--4448
		x"d3",	--4449
		x"d0",	--4450
		x"40",	--4451
		x"4a",	--4452
		x"00",	--4453
		x"4b",	--4454
		x"00",	--4455
		x"41",	--4456
		x"41",	--4457
		x"41",	--4458
		x"93",	--4459
		x"23",	--4460
		x"43",	--4461
		x"00",	--4462
		x"41",	--4463
		x"41",	--4464
		x"41",	--4465
		x"93",	--4466
		x"24",	--4467
		x"4a",	--4468
		x"4b",	--4469
		x"f3",	--4470
		x"f0",	--4471
		x"00",	--4472
		x"93",	--4473
		x"20",	--4474
		x"93",	--4475
		x"24",	--4476
		x"43",	--4477
		x"00",	--4478
		x"3f",	--4479
		x"93",	--4480
		x"23",	--4481
		x"42",	--4482
		x"00",	--4483
		x"3f",	--4484
		x"43",	--4485
		x"00",	--4486
		x"3f",	--4487
		x"12",	--4488
		x"4f",	--4489
		x"93",	--4490
		x"28",	--4491
		x"4e",	--4492
		x"93",	--4493
		x"28",	--4494
		x"92",	--4495
		x"24",	--4496
		x"92",	--4497
		x"24",	--4498
		x"93",	--4499
		x"24",	--4500
		x"93",	--4501
		x"24",	--4502
		x"4f",	--4503
		x"00",	--4504
		x"9e",	--4505
		x"00",	--4506
		x"24",	--4507
		x"93",	--4508
		x"20",	--4509
		x"43",	--4510
		x"4e",	--4511
		x"41",	--4512
		x"41",	--4513
		x"93",	--4514
		x"24",	--4515
		x"93",	--4516
		x"00",	--4517
		x"23",	--4518
		x"43",	--4519
		x"4e",	--4520
		x"41",	--4521
		x"41",	--4522
		x"93",	--4523
		x"00",	--4524
		x"27",	--4525
		x"43",	--4526
		x"3f",	--4527
		x"4f",	--4528
		x"00",	--4529
		x"4e",	--4530
		x"00",	--4531
		x"9b",	--4532
		x"3b",	--4533
		x"9c",	--4534
		x"38",	--4535
		x"4f",	--4536
		x"00",	--4537
		x"4f",	--4538
		x"00",	--4539
		x"4e",	--4540
		x"00",	--4541
		x"4e",	--4542
		x"00",	--4543
		x"9f",	--4544
		x"2b",	--4545
		x"9e",	--4546
		x"28",	--4547
		x"9b",	--4548
		x"2b",	--4549
		x"9e",	--4550
		x"28",	--4551
		x"9f",	--4552
		x"28",	--4553
		x"9c",	--4554
		x"28",	--4555
		x"43",	--4556
		x"3f",	--4557
		x"93",	--4558
		x"23",	--4559
		x"43",	--4560
		x"3f",	--4561
		x"92",	--4562
		x"23",	--4563
		x"4e",	--4564
		x"00",	--4565
		x"4f",	--4566
		x"00",	--4567
		x"8f",	--4568
		x"3f",	--4569
		x"42",	--4570
		x"02",	--4571
		x"93",	--4572
		x"38",	--4573
		x"42",	--4574
		x"02",	--4575
		x"4f",	--4576
		x"00",	--4577
		x"53",	--4578
		x"4d",	--4579
		x"02",	--4580
		x"53",	--4581
		x"4e",	--4582
		x"02",	--4583
		x"41",	--4584
		x"43",	--4585
		x"41",	--4586
		x"12",	--4587
		x"12",	--4588
		x"83",	--4589
		x"4e",	--4590
		x"00",	--4591
		x"42",	--4592
		x"02",	--4593
		x"42",	--4594
		x"02",	--4595
		x"4e",	--4596
		x"4f",	--4597
		x"40",	--4598
		x"e3",	--4599
		x"12",	--4600
		x"e6",	--4601
		x"9b",	--4602
		x"38",	--4603
		x"4a",	--4604
		x"5b",	--4605
		x"43",	--4606
		x"ff",	--4607
		x"3c",	--4608
		x"42",	--4609
		x"02",	--4610
		x"43",	--4611
		x"00",	--4612
		x"53",	--4613
		x"41",	--4614
		x"41",	--4615
		x"41",	--4616
		x"41",	--4617
		x"00",	--4618
		x"02",	--4619
		x"40",	--4620
		x"7f",	--4621
		x"02",	--4622
		x"41",	--4623
		x"50",	--4624
		x"00",	--4625
		x"41",	--4626
		x"00",	--4627
		x"12",	--4628
		x"e3",	--4629
		x"41",	--4630
		x"41",	--4631
		x"00",	--4632
		x"02",	--4633
		x"41",	--4634
		x"00",	--4635
		x"02",	--4636
		x"41",	--4637
		x"52",	--4638
		x"41",	--4639
		x"00",	--4640
		x"12",	--4641
		x"e3",	--4642
		x"41",	--4643
		x"4e",	--4644
		x"4f",	--4645
		x"02",	--4646
		x"40",	--4647
		x"7f",	--4648
		x"02",	--4649
		x"4d",	--4650
		x"4c",	--4651
		x"12",	--4652
		x"e3",	--4653
		x"41",	--4654
		x"4f",	--4655
		x"02",	--4656
		x"4e",	--4657
		x"02",	--4658
		x"4c",	--4659
		x"4d",	--4660
		x"12",	--4661
		x"e3",	--4662
		x"41",	--4663
		x"12",	--4664
		x"12",	--4665
		x"12",	--4666
		x"12",	--4667
		x"12",	--4668
		x"12",	--4669
		x"12",	--4670
		x"12",	--4671
		x"82",	--4672
		x"4f",	--4673
		x"4e",	--4674
		x"00",	--4675
		x"4d",	--4676
		x"41",	--4677
		x"00",	--4678
		x"41",	--4679
		x"00",	--4680
		x"4d",	--4681
		x"4d",	--4682
		x"10",	--4683
		x"44",	--4684
		x"4f",	--4685
		x"b0",	--4686
		x"00",	--4687
		x"24",	--4688
		x"40",	--4689
		x"00",	--4690
		x"00",	--4691
		x"4f",	--4692
		x"10",	--4693
		x"f3",	--4694
		x"24",	--4695
		x"40",	--4696
		x"00",	--4697
		x"3c",	--4698
		x"40",	--4699
		x"00",	--4700
		x"4e",	--4701
		x"00",	--4702
		x"41",	--4703
		x"53",	--4704
		x"3c",	--4705
		x"f0",	--4706
		x"00",	--4707
		x"24",	--4708
		x"40",	--4709
		x"00",	--4710
		x"00",	--4711
		x"3c",	--4712
		x"93",	--4713
		x"24",	--4714
		x"4d",	--4715
		x"00",	--4716
		x"41",	--4717
		x"53",	--4718
		x"3c",	--4719
		x"41",	--4720
		x"4c",	--4721
		x"10",	--4722
		x"11",	--4723
		x"10",	--4724
		x"11",	--4725
		x"4c",	--4726
		x"41",	--4727
		x"41",	--4728
		x"10",	--4729
		x"11",	--4730
		x"10",	--4731
		x"11",	--4732
		x"4c",	--4733
		x"86",	--4734
		x"77",	--4735
		x"4f",	--4736
		x"10",	--4737
		x"4e",	--4738
		x"00",	--4739
		x"f2",	--4740
		x"24",	--4741
		x"45",	--4742
		x"3c",	--4743
		x"43",	--4744
		x"4f",	--4745
		x"b0",	--4746
		x"00",	--4747
		x"20",	--4748
		x"41",	--4749
		x"00",	--4750
		x"53",	--4751
		x"53",	--4752
		x"93",	--4753
		x"00",	--4754
		x"23",	--4755
		x"81",	--4756
		x"00",	--4757
		x"9a",	--4758
		x"28",	--4759
		x"8a",	--4760
		x"3c",	--4761
		x"43",	--4762
		x"b3",	--4763
		x"00",	--4764
		x"24",	--4765
		x"95",	--4766
		x"28",	--4767
		x"85",	--4768
		x"3c",	--4769
		x"43",	--4770
		x"4d",	--4771
		x"9d",	--4772
		x"2c",	--4773
		x"47",	--4774
		x"93",	--4775
		x"38",	--4776
		x"40",	--4777
		x"00",	--4778
		x"00",	--4779
		x"43",	--4780
		x"43",	--4781
		x"3c",	--4782
		x"41",	--4783
		x"56",	--4784
		x"4f",	--4785
		x"11",	--4786
		x"53",	--4787
		x"12",	--4788
		x"3c",	--4789
		x"43",	--4790
		x"9a",	--4791
		x"3b",	--4792
		x"4a",	--4793
		x"40",	--4794
		x"00",	--4795
		x"00",	--4796
		x"8b",	--4797
		x"3c",	--4798
		x"41",	--4799
		x"00",	--4800
		x"11",	--4801
		x"12",	--4802
		x"53",	--4803
		x"45",	--4804
		x"5b",	--4805
		x"99",	--4806
		x"2b",	--4807
		x"3c",	--4808
		x"43",	--4809
		x"43",	--4810
		x"3c",	--4811
		x"53",	--4812
		x"41",	--4813
		x"56",	--4814
		x"4f",	--4815
		x"11",	--4816
		x"53",	--4817
		x"12",	--4818
		x"9a",	--4819
		x"3b",	--4820
		x"b3",	--4821
		x"00",	--4822
		x"24",	--4823
		x"44",	--4824
		x"3c",	--4825
		x"41",	--4826
		x"00",	--4827
		x"8b",	--4828
		x"3c",	--4829
		x"40",	--4830
		x"00",	--4831
		x"12",	--4832
		x"53",	--4833
		x"93",	--4834
		x"23",	--4835
		x"44",	--4836
		x"54",	--4837
		x"3f",	--4838
		x"53",	--4839
		x"11",	--4840
		x"12",	--4841
		x"53",	--4842
		x"4a",	--4843
		x"5b",	--4844
		x"4f",	--4845
		x"93",	--4846
		x"24",	--4847
		x"93",	--4848
		x"23",	--4849
		x"3c",	--4850
		x"40",	--4851
		x"00",	--4852
		x"12",	--4853
		x"53",	--4854
		x"99",	--4855
		x"2b",	--4856
		x"4b",	--4857
		x"52",	--4858
		x"41",	--4859
		x"41",	--4860
		x"41",	--4861
		x"41",	--4862
		x"41",	--4863
		x"41",	--4864
		x"41",	--4865
		x"41",	--4866
		x"41",	--4867
		x"12",	--4868
		x"12",	--4869
		x"12",	--4870
		x"12",	--4871
		x"12",	--4872
		x"12",	--4873
		x"12",	--4874
		x"12",	--4875
		x"50",	--4876
		x"ff",	--4877
		x"4f",	--4878
		x"00",	--4879
		x"4e",	--4880
		x"4d",	--4881
		x"4e",	--4882
		x"00",	--4883
		x"43",	--4884
		x"00",	--4885
		x"43",	--4886
		x"00",	--4887
		x"43",	--4888
		x"00",	--4889
		x"43",	--4890
		x"00",	--4891
		x"43",	--4892
		x"00",	--4893
		x"43",	--4894
		x"00",	--4895
		x"43",	--4896
		x"43",	--4897
		x"00",	--4898
		x"41",	--4899
		x"50",	--4900
		x"00",	--4901
		x"4e",	--4902
		x"00",	--4903
		x"40",	--4904
		x"ec",	--4905
		x"46",	--4906
		x"53",	--4907
		x"4f",	--4908
		x"00",	--4909
		x"93",	--4910
		x"20",	--4911
		x"90",	--4912
		x"00",	--4913
		x"20",	--4914
		x"43",	--4915
		x"00",	--4916
		x"43",	--4917
		x"00",	--4918
		x"46",	--4919
		x"00",	--4920
		x"43",	--4921
		x"00",	--4922
		x"43",	--4923
		x"00",	--4924
		x"43",	--4925
		x"00",	--4926
		x"43",	--4927
		x"00",	--4928
		x"43",	--4929
		x"00",	--4930
		x"40",	--4931
		x"ec",	--4932
		x"47",	--4933
		x"11",	--4934
		x"4e",	--4935
		x"12",	--4936
		x"00",	--4937
		x"53",	--4938
		x"00",	--4939
		x"40",	--4940
		x"ec",	--4941
		x"90",	--4942
		x"00",	--4943
		x"24",	--4944
		x"90",	--4945
		x"00",	--4946
		x"34",	--4947
		x"90",	--4948
		x"00",	--4949
		x"24",	--4950
		x"90",	--4951
		x"00",	--4952
		x"34",	--4953
		x"90",	--4954
		x"00",	--4955
		x"24",	--4956
		x"90",	--4957
		x"00",	--4958
		x"34",	--4959
		x"90",	--4960
		x"00",	--4961
		x"24",	--4962
		x"90",	--4963
		x"00",	--4964
		x"27",	--4965
		x"90",	--4966
		x"00",	--4967
		x"20",	--4968
		x"3c",	--4969
		x"90",	--4970
		x"00",	--4971
		x"24",	--4972
		x"90",	--4973
		x"00",	--4974
		x"24",	--4975
		x"90",	--4976
		x"00",	--4977
		x"20",	--4978
		x"3c",	--4979
		x"90",	--4980
		x"00",	--4981
		x"38",	--4982
		x"90",	--4983
		x"00",	--4984
		x"20",	--4985
		x"3c",	--4986
		x"90",	--4987
		x"00",	--4988
		x"24",	--4989
		x"90",	--4990
		x"00",	--4991
		x"34",	--4992
		x"90",	--4993
		x"00",	--4994
		x"24",	--4995
		x"90",	--4996
		x"00",	--4997
		x"24",	--4998
		x"90",	--4999
		x"00",	--5000
		x"20",	--5001
		x"3c",	--5002
		x"90",	--5003
		x"00",	--5004
		x"24",	--5005
		x"90",	--5006
		x"00",	--5007
		x"34",	--5008
		x"90",	--5009
		x"00",	--5010
		x"20",	--5011
		x"3c",	--5012
		x"90",	--5013
		x"00",	--5014
		x"24",	--5015
		x"90",	--5016
		x"00",	--5017
		x"24",	--5018
		x"41",	--5019
		x"00",	--5020
		x"41",	--5021
		x"00",	--5022
		x"89",	--5023
		x"40",	--5024
		x"ec",	--5025
		x"42",	--5026
		x"00",	--5027
		x"3c",	--5028
		x"d2",	--5029
		x"00",	--5030
		x"40",	--5031
		x"ec",	--5032
		x"41",	--5033
		x"f3",	--5034
		x"41",	--5035
		x"24",	--5036
		x"f0",	--5037
		x"ff",	--5038
		x"d3",	--5039
		x"3c",	--5040
		x"d3",	--5041
		x"4e",	--5042
		x"00",	--5043
		x"40",	--5044
		x"ec",	--5045
		x"d0",	--5046
		x"00",	--5047
		x"00",	--5048
		x"40",	--5049
		x"ec",	--5050
		x"40",	--5051
		x"00",	--5052
		x"00",	--5053
		x"40",	--5054
		x"ec",	--5055
		x"90",	--5056
		x"00",	--5057
		x"00",	--5058
		x"20",	--5059
		x"40",	--5060
		x"ec",	--5061
		x"40",	--5062
		x"00",	--5063
		x"00",	--5064
		x"40",	--5065
		x"ec",	--5066
		x"93",	--5067
		x"00",	--5068
		x"24",	--5069
		x"40",	--5070
		x"ec",	--5071
		x"43",	--5072
		x"00",	--5073
		x"40",	--5074
		x"ec",	--5075
		x"45",	--5076
		x"53",	--5077
		x"45",	--5078
		x"93",	--5079
		x"38",	--5080
		x"4a",	--5081
		x"00",	--5082
		x"3c",	--5083
		x"93",	--5084
		x"00",	--5085
		x"24",	--5086
		x"40",	--5087
		x"ec",	--5088
		x"d0",	--5089
		x"00",	--5090
		x"00",	--5091
		x"e3",	--5092
		x"4a",	--5093
		x"00",	--5094
		x"53",	--5095
		x"00",	--5096
		x"4e",	--5097
		x"3c",	--5098
		x"93",	--5099
		x"00",	--5100
		x"20",	--5101
		x"93",	--5102
		x"00",	--5103
		x"20",	--5104
		x"41",	--5105
		x"f0",	--5106
		x"00",	--5107
		x"43",	--5108
		x"24",	--5109
		x"43",	--5110
		x"4e",	--5111
		x"11",	--5112
		x"43",	--5113
		x"10",	--5114
		x"41",	--5115
		x"f0",	--5116
		x"00",	--5117
		x"de",	--5118
		x"4a",	--5119
		x"00",	--5120
		x"40",	--5121
		x"ec",	--5122
		x"41",	--5123
		x"00",	--5124
		x"5a",	--5125
		x"4a",	--5126
		x"5c",	--5127
		x"5c",	--5128
		x"5c",	--5129
		x"4a",	--5130
		x"00",	--5131
		x"50",	--5132
		x"ff",	--5133
		x"00",	--5134
		x"11",	--5135
		x"5e",	--5136
		x"00",	--5137
		x"43",	--5138
		x"00",	--5139
		x"40",	--5140
		x"ec",	--5141
		x"45",	--5142
		x"53",	--5143
		x"45",	--5144
		x"93",	--5145
		x"00",	--5146
		x"20",	--5147
		x"93",	--5148
		x"00",	--5149
		x"27",	--5150
		x"4e",	--5151
		x"00",	--5152
		x"43",	--5153
		x"00",	--5154
		x"41",	--5155
		x"52",	--5156
		x"3c",	--5157
		x"45",	--5158
		x"53",	--5159
		x"45",	--5160
		x"93",	--5161
		x"00",	--5162
		x"24",	--5163
		x"d2",	--5164
		x"00",	--5165
		x"41",	--5166
		x"00",	--5167
		x"4f",	--5168
		x"00",	--5169
		x"3c",	--5170
		x"93",	--5171
		x"00",	--5172
		x"24",	--5173
		x"41",	--5174
		x"00",	--5175
		x"00",	--5176
		x"93",	--5177
		x"20",	--5178
		x"40",	--5179
		x"f2",	--5180
		x"12",	--5181
		x"00",	--5182
		x"12",	--5183
		x"00",	--5184
		x"41",	--5185
		x"00",	--5186
		x"41",	--5187
		x"00",	--5188
		x"12",	--5189
		x"e4",	--5190
		x"52",	--5191
		x"5f",	--5192
		x"00",	--5193
		x"47",	--5194
		x"40",	--5195
		x"ec",	--5196
		x"45",	--5197
		x"53",	--5198
		x"45",	--5199
		x"49",	--5200
		x"00",	--5201
		x"43",	--5202
		x"93",	--5203
		x"20",	--5204
		x"43",	--5205
		x"5e",	--5206
		x"5e",	--5207
		x"5e",	--5208
		x"41",	--5209
		x"f0",	--5210
		x"ff",	--5211
		x"de",	--5212
		x"4a",	--5213
		x"00",	--5214
		x"47",	--5215
		x"40",	--5216
		x"00",	--5217
		x"00",	--5218
		x"3c",	--5219
		x"d3",	--5220
		x"00",	--5221
		x"3c",	--5222
		x"d2",	--5223
		x"00",	--5224
		x"40",	--5225
		x"00",	--5226
		x"00",	--5227
		x"3c",	--5228
		x"40",	--5229
		x"00",	--5230
		x"00",	--5231
		x"41",	--5232
		x"b3",	--5233
		x"24",	--5234
		x"45",	--5235
		x"52",	--5236
		x"45",	--5237
		x"45",	--5238
		x"00",	--5239
		x"45",	--5240
		x"00",	--5241
		x"45",	--5242
		x"00",	--5243
		x"48",	--5244
		x"00",	--5245
		x"47",	--5246
		x"00",	--5247
		x"46",	--5248
		x"00",	--5249
		x"4b",	--5250
		x"00",	--5251
		x"43",	--5252
		x"00",	--5253
		x"93",	--5254
		x"20",	--5255
		x"93",	--5256
		x"20",	--5257
		x"93",	--5258
		x"20",	--5259
		x"93",	--5260
		x"24",	--5261
		x"43",	--5262
		x"00",	--5263
		x"5b",	--5264
		x"43",	--5265
		x"6b",	--5266
		x"4b",	--5267
		x"00",	--5268
		x"4c",	--5269
		x"3c",	--5270
		x"f3",	--5271
		x"45",	--5272
		x"24",	--5273
		x"52",	--5274
		x"45",	--5275
		x"45",	--5276
		x"00",	--5277
		x"48",	--5278
		x"00",	--5279
		x"4b",	--5280
		x"00",	--5281
		x"43",	--5282
		x"00",	--5283
		x"93",	--5284
		x"20",	--5285
		x"3c",	--5286
		x"53",	--5287
		x"45",	--5288
		x"4b",	--5289
		x"00",	--5290
		x"43",	--5291
		x"00",	--5292
		x"93",	--5293
		x"24",	--5294
		x"43",	--5295
		x"00",	--5296
		x"5b",	--5297
		x"43",	--5298
		x"6b",	--5299
		x"4b",	--5300
		x"00",	--5301
		x"47",	--5302
		x"b2",	--5303
		x"00",	--5304
		x"24",	--5305
		x"93",	--5306
		x"00",	--5307
		x"20",	--5308
		x"41",	--5309
		x"90",	--5310
		x"00",	--5311
		x"00",	--5312
		x"20",	--5313
		x"d0",	--5314
		x"00",	--5315
		x"3c",	--5316
		x"92",	--5317
		x"00",	--5318
		x"20",	--5319
		x"d0",	--5320
		x"00",	--5321
		x"48",	--5322
		x"00",	--5323
		x"41",	--5324
		x"b2",	--5325
		x"24",	--5326
		x"93",	--5327
		x"00",	--5328
		x"24",	--5329
		x"40",	--5330
		x"00",	--5331
		x"00",	--5332
		x"b3",	--5333
		x"24",	--5334
		x"e3",	--5335
		x"00",	--5336
		x"e3",	--5337
		x"00",	--5338
		x"e3",	--5339
		x"00",	--5340
		x"e3",	--5341
		x"00",	--5342
		x"53",	--5343
		x"00",	--5344
		x"63",	--5345
		x"00",	--5346
		x"63",	--5347
		x"00",	--5348
		x"63",	--5349
		x"00",	--5350
		x"3c",	--5351
		x"b3",	--5352
		x"24",	--5353
		x"41",	--5354
		x"00",	--5355
		x"41",	--5356
		x"00",	--5357
		x"e3",	--5358
		x"e3",	--5359
		x"4a",	--5360
		x"4b",	--5361
		x"53",	--5362
		x"63",	--5363
		x"4e",	--5364
		x"00",	--5365
		x"4f",	--5366
		x"00",	--5367
		x"3c",	--5368
		x"41",	--5369
		x"00",	--5370
		x"e3",	--5371
		x"53",	--5372
		x"4a",	--5373
		x"00",	--5374
		x"43",	--5375
		x"00",	--5376
		x"b3",	--5377
		x"24",	--5378
		x"41",	--5379
		x"00",	--5380
		x"41",	--5381
		x"00",	--5382
		x"00",	--5383
		x"41",	--5384
		x"00",	--5385
		x"41",	--5386
		x"00",	--5387
		x"41",	--5388
		x"50",	--5389
		x"00",	--5390
		x"46",	--5391
		x"41",	--5392
		x"00",	--5393
		x"00",	--5394
		x"41",	--5395
		x"00",	--5396
		x"10",	--5397
		x"11",	--5398
		x"10",	--5399
		x"11",	--5400
		x"4b",	--5401
		x"00",	--5402
		x"4b",	--5403
		x"00",	--5404
		x"4b",	--5405
		x"00",	--5406
		x"12",	--5407
		x"00",	--5408
		x"12",	--5409
		x"00",	--5410
		x"12",	--5411
		x"00",	--5412
		x"12",	--5413
		x"00",	--5414
		x"49",	--5415
		x"41",	--5416
		x"00",	--5417
		x"48",	--5418
		x"44",	--5419
		x"12",	--5420
		x"ee",	--5421
		x"52",	--5422
		x"4c",	--5423
		x"90",	--5424
		x"00",	--5425
		x"34",	--5426
		x"50",	--5427
		x"00",	--5428
		x"4b",	--5429
		x"00",	--5430
		x"3c",	--5431
		x"4c",	--5432
		x"b3",	--5433
		x"00",	--5434
		x"24",	--5435
		x"40",	--5436
		x"00",	--5437
		x"3c",	--5438
		x"40",	--5439
		x"00",	--5440
		x"5b",	--5441
		x"4a",	--5442
		x"00",	--5443
		x"47",	--5444
		x"53",	--5445
		x"12",	--5446
		x"00",	--5447
		x"12",	--5448
		x"00",	--5449
		x"12",	--5450
		x"00",	--5451
		x"12",	--5452
		x"00",	--5453
		x"49",	--5454
		x"41",	--5455
		x"00",	--5456
		x"48",	--5457
		x"44",	--5458
		x"12",	--5459
		x"ed",	--5460
		x"52",	--5461
		x"4c",	--5462
		x"4d",	--5463
		x"00",	--5464
		x"4e",	--5465
		x"4f",	--5466
		x"53",	--5467
		x"93",	--5468
		x"23",	--5469
		x"93",	--5470
		x"23",	--5471
		x"93",	--5472
		x"23",	--5473
		x"93",	--5474
		x"23",	--5475
		x"43",	--5476
		x"00",	--5477
		x"43",	--5478
		x"00",	--5479
		x"43",	--5480
		x"00",	--5481
		x"43",	--5482
		x"00",	--5483
		x"3c",	--5484
		x"b3",	--5485
		x"24",	--5486
		x"41",	--5487
		x"00",	--5488
		x"41",	--5489
		x"00",	--5490
		x"41",	--5491
		x"50",	--5492
		x"00",	--5493
		x"41",	--5494
		x"00",	--5495
		x"10",	--5496
		x"11",	--5497
		x"10",	--5498
		x"11",	--5499
		x"41",	--5500
		x"00",	--5501
		x"49",	--5502
		x"44",	--5503
		x"47",	--5504
		x"12",	--5505
		x"ed",	--5506
		x"4e",	--5507
		x"90",	--5508
		x"00",	--5509
		x"34",	--5510
		x"50",	--5511
		x"00",	--5512
		x"4b",	--5513
		x"00",	--5514
		x"3c",	--5515
		x"4e",	--5516
		x"b3",	--5517
		x"00",	--5518
		x"24",	--5519
		x"40",	--5520
		x"00",	--5521
		x"3c",	--5522
		x"40",	--5523
		x"00",	--5524
		x"5b",	--5525
		x"4a",	--5526
		x"00",	--5527
		x"48",	--5528
		x"53",	--5529
		x"41",	--5530
		x"00",	--5531
		x"49",	--5532
		x"44",	--5533
		x"47",	--5534
		x"12",	--5535
		x"ec",	--5536
		x"4e",	--5537
		x"4f",	--5538
		x"53",	--5539
		x"93",	--5540
		x"23",	--5541
		x"93",	--5542
		x"23",	--5543
		x"43",	--5544
		x"00",	--5545
		x"43",	--5546
		x"00",	--5547
		x"3c",	--5548
		x"41",	--5549
		x"00",	--5550
		x"41",	--5551
		x"50",	--5552
		x"00",	--5553
		x"41",	--5554
		x"00",	--5555
		x"47",	--5556
		x"12",	--5557
		x"ed",	--5558
		x"4f",	--5559
		x"90",	--5560
		x"00",	--5561
		x"34",	--5562
		x"50",	--5563
		x"00",	--5564
		x"4d",	--5565
		x"00",	--5566
		x"3c",	--5567
		x"4f",	--5568
		x"b3",	--5569
		x"00",	--5570
		x"24",	--5571
		x"40",	--5572
		x"00",	--5573
		x"3c",	--5574
		x"40",	--5575
		x"00",	--5576
		x"5d",	--5577
		x"4c",	--5578
		x"00",	--5579
		x"48",	--5580
		x"53",	--5581
		x"41",	--5582
		x"00",	--5583
		x"47",	--5584
		x"12",	--5585
		x"ed",	--5586
		x"4f",	--5587
		x"53",	--5588
		x"93",	--5589
		x"23",	--5590
		x"43",	--5591
		x"00",	--5592
		x"90",	--5593
		x"00",	--5594
		x"00",	--5595
		x"24",	--5596
		x"43",	--5597
		x"00",	--5598
		x"93",	--5599
		x"00",	--5600
		x"24",	--5601
		x"41",	--5602
		x"50",	--5603
		x"00",	--5604
		x"4f",	--5605
		x"00",	--5606
		x"41",	--5607
		x"00",	--5608
		x"10",	--5609
		x"11",	--5610
		x"10",	--5611
		x"11",	--5612
		x"4a",	--5613
		x"00",	--5614
		x"46",	--5615
		x"00",	--5616
		x"46",	--5617
		x"10",	--5618
		x"11",	--5619
		x"10",	--5620
		x"11",	--5621
		x"4a",	--5622
		x"00",	--5623
		x"41",	--5624
		x"00",	--5625
		x"41",	--5626
		x"00",	--5627
		x"81",	--5628
		x"00",	--5629
		x"71",	--5630
		x"00",	--5631
		x"83",	--5632
		x"91",	--5633
		x"00",	--5634
		x"2c",	--5635
		x"d3",	--5636
		x"00",	--5637
		x"41",	--5638
		x"00",	--5639
		x"8c",	--5640
		x"4e",	--5641
		x"00",	--5642
		x"3c",	--5643
		x"93",	--5644
		x"00",	--5645
		x"24",	--5646
		x"41",	--5647
		x"00",	--5648
		x"00",	--5649
		x"12",	--5650
		x"00",	--5651
		x"12",	--5652
		x"00",	--5653
		x"41",	--5654
		x"00",	--5655
		x"46",	--5656
		x"53",	--5657
		x"41",	--5658
		x"00",	--5659
		x"12",	--5660
		x"e4",	--5661
		x"52",	--5662
		x"5f",	--5663
		x"00",	--5664
		x"3c",	--5665
		x"49",	--5666
		x"11",	--5667
		x"12",	--5668
		x"00",	--5669
		x"49",	--5670
		x"58",	--5671
		x"91",	--5672
		x"00",	--5673
		x"2b",	--5674
		x"49",	--5675
		x"00",	--5676
		x"4e",	--5677
		x"00",	--5678
		x"43",	--5679
		x"3c",	--5680
		x"41",	--5681
		x"00",	--5682
		x"00",	--5683
		x"43",	--5684
		x"00",	--5685
		x"43",	--5686
		x"00",	--5687
		x"3c",	--5688
		x"4e",	--5689
		x"43",	--5690
		x"00",	--5691
		x"43",	--5692
		x"00",	--5693
		x"43",	--5694
		x"41",	--5695
		x"00",	--5696
		x"46",	--5697
		x"93",	--5698
		x"24",	--5699
		x"40",	--5700
		x"e6",	--5701
		x"41",	--5702
		x"00",	--5703
		x"50",	--5704
		x"00",	--5705
		x"41",	--5706
		x"41",	--5707
		x"41",	--5708
		x"41",	--5709
		x"41",	--5710
		x"41",	--5711
		x"41",	--5712
		x"41",	--5713
		x"41",	--5714
		x"43",	--5715
		x"93",	--5716
		x"34",	--5717
		x"40",	--5718
		x"00",	--5719
		x"e3",	--5720
		x"53",	--5721
		x"93",	--5722
		x"34",	--5723
		x"e3",	--5724
		x"e3",	--5725
		x"53",	--5726
		x"12",	--5727
		x"12",	--5728
		x"ed",	--5729
		x"41",	--5730
		x"b3",	--5731
		x"24",	--5732
		x"e3",	--5733
		x"53",	--5734
		x"b3",	--5735
		x"24",	--5736
		x"e3",	--5737
		x"53",	--5738
		x"41",	--5739
		x"12",	--5740
		x"ec",	--5741
		x"4e",	--5742
		x"41",	--5743
		x"12",	--5744
		x"12",	--5745
		x"12",	--5746
		x"40",	--5747
		x"00",	--5748
		x"4c",	--5749
		x"4d",	--5750
		x"43",	--5751
		x"43",	--5752
		x"5e",	--5753
		x"6f",	--5754
		x"6c",	--5755
		x"6d",	--5756
		x"9b",	--5757
		x"28",	--5758
		x"20",	--5759
		x"9a",	--5760
		x"28",	--5761
		x"8a",	--5762
		x"7b",	--5763
		x"d3",	--5764
		x"83",	--5765
		x"23",	--5766
		x"41",	--5767
		x"41",	--5768
		x"41",	--5769
		x"41",	--5770
		x"12",	--5771
		x"ec",	--5772
		x"4c",	--5773
		x"4d",	--5774
		x"41",	--5775
		x"12",	--5776
		x"43",	--5777
		x"93",	--5778
		x"34",	--5779
		x"40",	--5780
		x"00",	--5781
		x"e3",	--5782
		x"e3",	--5783
		x"53",	--5784
		x"63",	--5785
		x"93",	--5786
		x"34",	--5787
		x"e3",	--5788
		x"e3",	--5789
		x"e3",	--5790
		x"53",	--5791
		x"63",	--5792
		x"12",	--5793
		x"ec",	--5794
		x"b3",	--5795
		x"24",	--5796
		x"e3",	--5797
		x"e3",	--5798
		x"53",	--5799
		x"63",	--5800
		x"b3",	--5801
		x"24",	--5802
		x"e3",	--5803
		x"e3",	--5804
		x"53",	--5805
		x"63",	--5806
		x"41",	--5807
		x"41",	--5808
		x"12",	--5809
		x"ed",	--5810
		x"4c",	--5811
		x"4d",	--5812
		x"41",	--5813
		x"40",	--5814
		x"00",	--5815
		x"4e",	--5816
		x"43",	--5817
		x"5f",	--5818
		x"6e",	--5819
		x"9d",	--5820
		x"28",	--5821
		x"8d",	--5822
		x"d3",	--5823
		x"83",	--5824
		x"23",	--5825
		x"41",	--5826
		x"12",	--5827
		x"ed",	--5828
		x"4e",	--5829
		x"41",	--5830
		x"12",	--5831
		x"12",	--5832
		x"12",	--5833
		x"12",	--5834
		x"12",	--5835
		x"00",	--5836
		x"48",	--5837
		x"49",	--5838
		x"4a",	--5839
		x"4b",	--5840
		x"43",	--5841
		x"43",	--5842
		x"43",	--5843
		x"43",	--5844
		x"5c",	--5845
		x"6d",	--5846
		x"6e",	--5847
		x"6f",	--5848
		x"68",	--5849
		x"69",	--5850
		x"6a",	--5851
		x"6b",	--5852
		x"97",	--5853
		x"28",	--5854
		x"20",	--5855
		x"96",	--5856
		x"28",	--5857
		x"20",	--5858
		x"95",	--5859
		x"28",	--5860
		x"20",	--5861
		x"94",	--5862
		x"28",	--5863
		x"84",	--5864
		x"75",	--5865
		x"76",	--5866
		x"77",	--5867
		x"d3",	--5868
		x"83",	--5869
		x"00",	--5870
		x"23",	--5871
		x"53",	--5872
		x"41",	--5873
		x"41",	--5874
		x"41",	--5875
		x"41",	--5876
		x"41",	--5877
		x"12",	--5878
		x"12",	--5879
		x"12",	--5880
		x"12",	--5881
		x"41",	--5882
		x"00",	--5883
		x"41",	--5884
		x"00",	--5885
		x"41",	--5886
		x"00",	--5887
		x"41",	--5888
		x"00",	--5889
		x"12",	--5890
		x"ed",	--5891
		x"41",	--5892
		x"41",	--5893
		x"41",	--5894
		x"41",	--5895
		x"41",	--5896
		x"12",	--5897
		x"12",	--5898
		x"12",	--5899
		x"12",	--5900
		x"41",	--5901
		x"00",	--5902
		x"41",	--5903
		x"00",	--5904
		x"41",	--5905
		x"00",	--5906
		x"41",	--5907
		x"00",	--5908
		x"12",	--5909
		x"ed",	--5910
		x"48",	--5911
		x"49",	--5912
		x"4a",	--5913
		x"4b",	--5914
		x"41",	--5915
		x"41",	--5916
		x"41",	--5917
		x"41",	--5918
		x"41",	--5919
		x"12",	--5920
		x"12",	--5921
		x"12",	--5922
		x"12",	--5923
		x"12",	--5924
		x"41",	--5925
		x"00",	--5926
		x"41",	--5927
		x"00",	--5928
		x"41",	--5929
		x"00",	--5930
		x"41",	--5931
		x"00",	--5932
		x"12",	--5933
		x"ed",	--5934
		x"41",	--5935
		x"00",	--5936
		x"48",	--5937
		x"00",	--5938
		x"49",	--5939
		x"00",	--5940
		x"4a",	--5941
		x"00",	--5942
		x"4b",	--5943
		x"00",	--5944
		x"41",	--5945
		x"41",	--5946
		x"41",	--5947
		x"41",	--5948
		x"41",	--5949
		x"41",	--5950
		x"13",	--5951
		x"d0",	--5952
		x"00",	--5953
		x"3f",	--5954
		x"64",	--5955
		x"00",	--5956
		x"0a",	--5957
		x"53",	--5958
		x"6f",	--5959
		x"0d",	--5960
		x"00",	--5961
		x"6f",	--5962
		x"72",	--5963
		x"63",	--5964
		x"20",	--5965
		x"73",	--5966
		x"67",	--5967
		x"3a",	--5968
		x"0a",	--5969
		x"09",	--5970
		x"63",	--5971
		x"4c",	--5972
		x"46",	--5973
		x"20",	--5974
		x"49",	--5975
		x"48",	--5976
		x"20",	--5977
		x"54",	--5978
		x"4d",	--5979
		x"4f",	--5980
		x"54",	--5981
		x"0d",	--5982
		x"00",	--5983
		x"64",	--5984
		x"25",	--5985
		x"0d",	--5986
		x"00",	--5987
		x"6f",	--5988
		x"20",	--5989
		x"6d",	--5990
		x"6c",	--5991
		x"6d",	--5992
		x"6e",	--5993
		x"65",	--5994
		x"20",	--5995
		x"65",	--5996
		x"0d",	--5997
		x"00",	--5998
		x"61",	--5999
		x"74",	--6000
		x"6e",	--6001
		x"20",	--6002
		x"6f",	--6003
		x"20",	--6004
		x"20",	--6005
		x"65",	--6006
		x"20",	--6007
		x"62",	--6008
		x"6e",	--6009
		x"66",	--6010
		x"6c",	--6011
		x"0d",	--6012
		x"00",	--6013
		x"65",	--6014
		x"73",	--6015
		x"6f",	--6016
		x"6c",	--6017
		x"20",	--6018
		x"6f",	--6019
		x"20",	--6020
		x"65",	--6021
		x"20",	--6022
		x"68",	--6023
		x"74",	--6024
		x"0a",	--6025
		x"53",	--6026
		x"6f",	--6027
		x"0d",	--6028
		x"00",	--6029
		x"72",	--6030
		x"6f",	--6031
		x"3a",	--6032
		x"6d",	--6033
		x"73",	--6034
		x"69",	--6035
		x"67",	--6036
		x"61",	--6037
		x"67",	--6038
		x"6d",	--6039
		x"6e",	--6040
		x"0d",	--6041
		x"00",	--6042
		x"6f",	--6043
		x"72",	--6044
		x"63",	--6045
		x"20",	--6046
		x"73",	--6047
		x"67",	--6048
		x"3a",	--6049
		x"0a",	--6050
		x"09",	--6051
		x"73",	--6052
		x"4c",	--6053
		x"46",	--6054
		x"20",	--6055
		x"49",	--6056
		x"48",	--6057
		x"20",	--6058
		x"54",	--6059
		x"4d",	--6060
		x"4f",	--6061
		x"54",	--6062
		x"0d",	--6063
		x"00",	--6064
		x"64",	--6065
		x"25",	--6066
		x"0d",	--6067
		x"00",	--6068
		x"6c",	--6069
		x"20",	--6070
		x"6c",	--6071
		x"00",	--6072
		x"73",	--6073
		x"0a",	--6074
		x"25",	--6075
		x"20",	--6076
		x"64",	--6077
		x"0a",	--6078
		x"00",	--6079
		x"ca",	--6080
		x"ca",	--6081
		x"ca",	--6082
		x"ca",	--6083
		x"ca",	--6084
		x"ca",	--6085
		x"ca",	--6086
		x"ca",	--6087
		x"0a",	--6088
		x"3d",	--6089
		x"3d",	--6090
		x"3d",	--6091
		x"4d",	--6092
		x"72",	--6093
		x"65",	--6094
		x"20",	--6095
		x"43",	--6096
		x"20",	--6097
		x"3d",	--6098
		x"3d",	--6099
		x"3d",	--6100
		x"0a",	--6101
		x"69",	--6102
		x"74",	--6103
		x"72",	--6104
		x"63",	--6105
		x"69",	--6106
		x"65",	--6107
		x"6d",	--6108
		x"64",	--6109
		x"00",	--6110
		x"72",	--6111
		x"74",	--6112
		x"00",	--6113
		x"65",	--6114
		x"64",	--6115
		x"62",	--6116
		x"7a",	--6117
		x"65",	--6118
		x"00",	--6119
		x"77",	--6120
		x"00",	--6121
		x"6e",	--6122
		x"6f",	--6123
		x"65",	--6124
		x"00",	--6125
		x"70",	--6126
		x"65",	--6127
		x"20",	--6128
		x"6f",	--6129
		x"74",	--6130
		x"6f",	--6131
		x"6c",	--6132
		x"72",	--6133
		x"73",	--6134
		x"65",	--6135
		x"64",	--6136
		x"63",	--6137
		x"6e",	--6138
		x"69",	--6139
		x"75",	--6140
		x"61",	--6141
		x"69",	--6142
		x"6e",	--6143
		x"73",	--6144
		x"66",	--6145
		x"35",	--6146
		x"62",	--6147
		x"6f",	--6148
		x"6c",	--6149
		x"61",	--6150
		x"65",	--6151
		x"00",	--6152
		x"0a",	--6153
		x"08",	--6154
		x"08",	--6155
		x"25",	--6156
		x"00",	--6157
		x"50",	--6158
		x"0a",	--6159
		x"44",	--6160
		x"57",	--6161
		x"0d",	--6162
		x"00",	--6163
		x"49",	--6164
		x"48",	--6165
		x"0d",	--6166
		x"00",	--6167
		x"45",	--6168
		x"54",	--6169
		x"0a",	--6170
		x"00",	--6171
		x"72",	--6172
		x"74",	--6173
		x"0a",	--6174
		x"00",	--6175
		x"72",	--6176
		x"6f",	--6177
		x"3a",	--6178
		x"6d",	--6179
		x"73",	--6180
		x"69",	--6181
		x"67",	--6182
		x"61",	--6183
		x"67",	--6184
		x"6d",	--6185
		x"6e",	--6186
		x"0d",	--6187
		x"00",	--6188
		x"6f",	--6189
		x"72",	--6190
		x"63",	--6191
		x"20",	--6192
		x"73",	--6193
		x"67",	--6194
		x"3a",	--6195
		x"0a",	--6196
		x"09",	--6197
		x"73",	--6198
		x"52",	--6199
		x"47",	--6200
		x"53",	--6201
		x"45",	--6202
		x"20",	--6203
		x"41",	--6204
		x"55",	--6205
		x"0d",	--6206
		x"00",	--6207
		x"3d",	--6208
		x"64",	--6209
		x"76",	--6210
		x"25",	--6211
		x"0d",	--6212
		x"00",	--6213
		x"25",	--6214
		x"20",	--6215
		x"45",	--6216
		x"49",	--6217
		x"54",	--6218
		x"52",	--6219
		x"0a",	--6220
		x"72",	--6221
		x"61",	--6222
		x"0a",	--6223
		x"00",	--6224
		x"63",	--6225
		x"69",	--6226
		x"20",	--6227
		x"6f",	--6228
		x"20",	--6229
		x"20",	--6230
		x"75",	--6231
		x"62",	--6232
		x"72",	--6233
		x"0a",	--6234
		x"25",	--6235
		x"20",	--6236
		x"73",	--6237
		x"0a",	--6238
		x"25",	--6239
		x"3a",	--6240
		x"6e",	--6241
		x"20",	--6242
		x"75",	--6243
		x"68",	--6244
		x"63",	--6245
		x"6d",	--6246
		x"61",	--6247
		x"64",	--6248
		x"0a",	--6249
		x"00",	--6250
		x"d4",	--6251
		x"d4",	--6252
		x"d4",	--6253
		x"d4",	--6254
		x"d4",	--6255
		x"d4",	--6256
		x"d4",	--6257
		x"d4",	--6258
		x"d4",	--6259
		x"d4",	--6260
		x"d4",	--6261
		x"d4",	--6262
		x"d4",	--6263
		x"d4",	--6264
		x"d4",	--6265
		x"d4",	--6266
		x"d4",	--6267
		x"d4",	--6268
		x"d4",	--6269
		x"d4",	--6270
		x"d4",	--6271
		x"d4",	--6272
		x"d4",	--6273
		x"d4",	--6274
		x"d4",	--6275
		x"d4",	--6276
		x"d4",	--6277
		x"d4",	--6278
		x"d4",	--6279
		x"d4",	--6280
		x"d4",	--6281
		x"d4",	--6282
		x"d4",	--6283
		x"d4",	--6284
		x"d4",	--6285
		x"d4",	--6286
		x"d4",	--6287
		x"d4",	--6288
		x"d4",	--6289
		x"d4",	--6290
		x"d4",	--6291
		x"d4",	--6292
		x"d4",	--6293
		x"d4",	--6294
		x"d4",	--6295
		x"d4",	--6296
		x"d4",	--6297
		x"d4",	--6298
		x"d4",	--6299
		x"d4",	--6300
		x"d4",	--6301
		x"d4",	--6302
		x"d4",	--6303
		x"d4",	--6304
		x"d4",	--6305
		x"d4",	--6306
		x"d4",	--6307
		x"d4",	--6308
		x"d4",	--6309
		x"d4",	--6310
		x"d4",	--6311
		x"d4",	--6312
		x"d4",	--6313
		x"d4",	--6314
		x"d4",	--6315
		x"d4",	--6316
		x"d4",	--6317
		x"d4",	--6318
		x"d4",	--6319
		x"d4",	--6320
		x"d4",	--6321
		x"d4",	--6322
		x"d4",	--6323
		x"d4",	--6324
		x"d4",	--6325
		x"d4",	--6326
		x"d4",	--6327
		x"d4",	--6328
		x"d4",	--6329
		x"d4",	--6330
		x"d4",	--6331
		x"d4",	--6332
		x"d4",	--6333
		x"d4",	--6334
		x"31",	--6335
		x"33",	--6336
		x"35",	--6337
		x"37",	--6338
		x"39",	--6339
		x"62",	--6340
		x"64",	--6341
		x"66",	--6342
		x"00",	--6343
		x"00",	--6344
		x"00",	--6345
		x"00",	--6346
		x"00",	--6347
		x"01",	--6348
		x"02",	--6349
		x"03",	--6350
		x"03",	--6351
		x"04",	--6352
		x"04",	--6353
		x"04",	--6354
		x"04",	--6355
		x"05",	--6356
		x"05",	--6357
		x"05",	--6358
		x"05",	--6359
		x"05",	--6360
		x"05",	--6361
		x"05",	--6362
		x"05",	--6363
		x"06",	--6364
		x"06",	--6365
		x"06",	--6366
		x"06",	--6367
		x"06",	--6368
		x"06",	--6369
		x"06",	--6370
		x"06",	--6371
		x"06",	--6372
		x"06",	--6373
		x"06",	--6374
		x"06",	--6375
		x"06",	--6376
		x"06",	--6377
		x"06",	--6378
		x"06",	--6379
		x"07",	--6380
		x"07",	--6381
		x"07",	--6382
		x"07",	--6383
		x"07",	--6384
		x"07",	--6385
		x"07",	--6386
		x"07",	--6387
		x"07",	--6388
		x"07",	--6389
		x"07",	--6390
		x"07",	--6391
		x"07",	--6392
		x"07",	--6393
		x"07",	--6394
		x"07",	--6395
		x"07",	--6396
		x"07",	--6397
		x"07",	--6398
		x"07",	--6399
		x"07",	--6400
		x"07",	--6401
		x"07",	--6402
		x"07",	--6403
		x"07",	--6404
		x"07",	--6405
		x"07",	--6406
		x"07",	--6407
		x"07",	--6408
		x"07",	--6409
		x"07",	--6410
		x"07",	--6411
		x"08",	--6412
		x"08",	--6413
		x"08",	--6414
		x"08",	--6415
		x"08",	--6416
		x"08",	--6417
		x"08",	--6418
		x"08",	--6419
		x"08",	--6420
		x"08",	--6421
		x"08",	--6422
		x"08",	--6423
		x"08",	--6424
		x"08",	--6425
		x"08",	--6426
		x"08",	--6427
		x"08",	--6428
		x"08",	--6429
		x"08",	--6430
		x"08",	--6431
		x"08",	--6432
		x"08",	--6433
		x"08",	--6434
		x"08",	--6435
		x"08",	--6436
		x"08",	--6437
		x"08",	--6438
		x"08",	--6439
		x"08",	--6440
		x"08",	--6441
		x"08",	--6442
		x"08",	--6443
		x"08",	--6444
		x"08",	--6445
		x"08",	--6446
		x"08",	--6447
		x"08",	--6448
		x"08",	--6449
		x"08",	--6450
		x"08",	--6451
		x"08",	--6452
		x"08",	--6453
		x"08",	--6454
		x"08",	--6455
		x"08",	--6456
		x"08",	--6457
		x"08",	--6458
		x"08",	--6459
		x"08",	--6460
		x"08",	--6461
		x"08",	--6462
		x"08",	--6463
		x"08",	--6464
		x"08",	--6465
		x"08",	--6466
		x"08",	--6467
		x"08",	--6468
		x"08",	--6469
		x"08",	--6470
		x"08",	--6471
		x"08",	--6472
		x"08",	--6473
		x"08",	--6474
		x"08",	--6475
		x"6e",	--6476
		x"6c",	--6477
		x"29",	--6478
		x"00",	--6479
		x"ff",	--6480
		x"ff",	--6481
		x"ff",	--6482
		x"ff",	--6483
		x"65",	--6484
		x"70",	--6485
		x"00",	--6486
		x"ff",	--6487
		x"ff",	--6488
		x"ff",	--6489
		x"ff",	--6490
		x"ff",	--6491
		x"ff",	--6492
		x"ff",	--6493
		x"ff",	--6494
		x"ff",	--6495
		x"ff",	--6496
		x"ff",	--6497
		x"ff",	--6498
		x"ff",	--6499
		x"ff",	--6500
		x"ff",	--6501
		x"ff",	--6502
		x"ff",	--6503
		x"ff",	--6504
		x"ff",	--6505
		x"ff",	--6506
		x"ff",	--6507
		x"ff",	--6508
		x"ff",	--6509
		x"ff",	--6510
		x"ff",	--6511
		x"ff",	--6512
		x"ff",	--6513
		x"ff",	--6514
		x"ff",	--6515
		x"ff",	--6516
		x"ff",	--6517
		x"ff",	--6518
		x"ff",	--6519
		x"ff",	--6520
		x"ff",	--6521
		x"ff",	--6522
		x"ff",	--6523
		x"ff",	--6524
		x"ff",	--6525
		x"ff",	--6526
		x"ff",	--6527
		x"ff",	--6528
		x"ff",	--6529
		x"ff",	--6530
		x"ff",	--6531
		x"ff",	--6532
		x"ff",	--6533
		x"ff",	--6534
		x"ff",	--6535
		x"ff",	--6536
		x"ff",	--6537
		x"ff",	--6538
		x"ff",	--6539
		x"ff",	--6540
		x"ff",	--6541
		x"ff",	--6542
		x"ff",	--6543
		x"ff",	--6544
		x"ff",	--6545
		x"ff",	--6546
		x"ff",	--6547
		x"ff",	--6548
		x"ff",	--6549
		x"ff",	--6550
		x"ff",	--6551
		x"ff",	--6552
		x"ff",	--6553
		x"ff",	--6554
		x"ff",	--6555
		x"ff",	--6556
		x"ff",	--6557
		x"ff",	--6558
		x"ff",	--6559
		x"ff",	--6560
		x"ff",	--6561
		x"ff",	--6562
		x"ff",	--6563
		x"ff",	--6564
		x"ff",	--6565
		x"ff",	--6566
		x"ff",	--6567
		x"ff",	--6568
		x"ff",	--6569
		x"ff",	--6570
		x"ff",	--6571
		x"ff",	--6572
		x"ff",	--6573
		x"ff",	--6574
		x"ff",	--6575
		x"ff",	--6576
		x"ff",	--6577
		x"ff",	--6578
		x"ff",	--6579
		x"ff",	--6580
		x"ff",	--6581
		x"ff",	--6582
		x"ff",	--6583
		x"ff",	--6584
		x"ff",	--6585
		x"ff",	--6586
		x"ff",	--6587
		x"ff",	--6588
		x"ff",	--6589
		x"ff",	--6590
		x"ff",	--6591
		x"ff",	--6592
		x"ff",	--6593
		x"ff",	--6594
		x"ff",	--6595
		x"ff",	--6596
		x"ff",	--6597
		x"ff",	--6598
		x"ff",	--6599
		x"ff",	--6600
		x"ff",	--6601
		x"ff",	--6602
		x"ff",	--6603
		x"ff",	--6604
		x"ff",	--6605
		x"ff",	--6606
		x"ff",	--6607
		x"ff",	--6608
		x"ff",	--6609
		x"ff",	--6610
		x"ff",	--6611
		x"ff",	--6612
		x"ff",	--6613
		x"ff",	--6614
		x"ff",	--6615
		x"ff",	--6616
		x"ff",	--6617
		x"ff",	--6618
		x"ff",	--6619
		x"ff",	--6620
		x"ff",	--6621
		x"ff",	--6622
		x"ff",	--6623
		x"ff",	--6624
		x"ff",	--6625
		x"ff",	--6626
		x"ff",	--6627
		x"ff",	--6628
		x"ff",	--6629
		x"ff",	--6630
		x"ff",	--6631
		x"ff",	--6632
		x"ff",	--6633
		x"ff",	--6634
		x"ff",	--6635
		x"ff",	--6636
		x"ff",	--6637
		x"ff",	--6638
		x"ff",	--6639
		x"ff",	--6640
		x"ff",	--6641
		x"ff",	--6642
		x"ff",	--6643
		x"ff",	--6644
		x"ff",	--6645
		x"ff",	--6646
		x"ff",	--6647
		x"ff",	--6648
		x"ff",	--6649
		x"ff",	--6650
		x"ff",	--6651
		x"ff",	--6652
		x"ff",	--6653
		x"ff",	--6654
		x"ff",	--6655
		x"ff",	--6656
		x"ff",	--6657
		x"ff",	--6658
		x"ff",	--6659
		x"ff",	--6660
		x"ff",	--6661
		x"ff",	--6662
		x"ff",	--6663
		x"ff",	--6664
		x"ff",	--6665
		x"ff",	--6666
		x"ff",	--6667
		x"ff",	--6668
		x"ff",	--6669
		x"ff",	--6670
		x"ff",	--6671
		x"ff",	--6672
		x"ff",	--6673
		x"ff",	--6674
		x"ff",	--6675
		x"ff",	--6676
		x"ff",	--6677
		x"ff",	--6678
		x"ff",	--6679
		x"ff",	--6680
		x"ff",	--6681
		x"ff",	--6682
		x"ff",	--6683
		x"ff",	--6684
		x"ff",	--6685
		x"ff",	--6686
		x"ff",	--6687
		x"ff",	--6688
		x"ff",	--6689
		x"ff",	--6690
		x"ff",	--6691
		x"ff",	--6692
		x"ff",	--6693
		x"ff",	--6694
		x"ff",	--6695
		x"ff",	--6696
		x"ff",	--6697
		x"ff",	--6698
		x"ff",	--6699
		x"ff",	--6700
		x"ff",	--6701
		x"ff",	--6702
		x"ff",	--6703
		x"ff",	--6704
		x"ff",	--6705
		x"ff",	--6706
		x"ff",	--6707
		x"ff",	--6708
		x"ff",	--6709
		x"ff",	--6710
		x"ff",	--6711
		x"ff",	--6712
		x"ff",	--6713
		x"ff",	--6714
		x"ff",	--6715
		x"ff",	--6716
		x"ff",	--6717
		x"ff",	--6718
		x"ff",	--6719
		x"ff",	--6720
		x"ff",	--6721
		x"ff",	--6722
		x"ff",	--6723
		x"ff",	--6724
		x"ff",	--6725
		x"ff",	--6726
		x"ff",	--6727
		x"ff",	--6728
		x"ff",	--6729
		x"ff",	--6730
		x"ff",	--6731
		x"ff",	--6732
		x"ff",	--6733
		x"ff",	--6734
		x"ff",	--6735
		x"ff",	--6736
		x"ff",	--6737
		x"ff",	--6738
		x"ff",	--6739
		x"ff",	--6740
		x"ff",	--6741
		x"ff",	--6742
		x"ff",	--6743
		x"ff",	--6744
		x"ff",	--6745
		x"ff",	--6746
		x"ff",	--6747
		x"ff",	--6748
		x"ff",	--6749
		x"ff",	--6750
		x"ff",	--6751
		x"ff",	--6752
		x"ff",	--6753
		x"ff",	--6754
		x"ff",	--6755
		x"ff",	--6756
		x"ff",	--6757
		x"ff",	--6758
		x"ff",	--6759
		x"ff",	--6760
		x"ff",	--6761
		x"ff",	--6762
		x"ff",	--6763
		x"ff",	--6764
		x"ff",	--6765
		x"ff",	--6766
		x"ff",	--6767
		x"ff",	--6768
		x"ff",	--6769
		x"ff",	--6770
		x"ff",	--6771
		x"ff",	--6772
		x"ff",	--6773
		x"ff",	--6774
		x"ff",	--6775
		x"ff",	--6776
		x"ff",	--6777
		x"ff",	--6778
		x"ff",	--6779
		x"ff",	--6780
		x"ff",	--6781
		x"ff",	--6782
		x"ff",	--6783
		x"ff",	--6784
		x"ff",	--6785
		x"ff",	--6786
		x"ff",	--6787
		x"ff",	--6788
		x"ff",	--6789
		x"ff",	--6790
		x"ff",	--6791
		x"ff",	--6792
		x"ff",	--6793
		x"ff",	--6794
		x"ff",	--6795
		x"ff",	--6796
		x"ff",	--6797
		x"ff",	--6798
		x"ff",	--6799
		x"ff",	--6800
		x"ff",	--6801
		x"ff",	--6802
		x"ff",	--6803
		x"ff",	--6804
		x"ff",	--6805
		x"ff",	--6806
		x"ff",	--6807
		x"ff",	--6808
		x"ff",	--6809
		x"ff",	--6810
		x"ff",	--6811
		x"ff",	--6812
		x"ff",	--6813
		x"ff",	--6814
		x"ff",	--6815
		x"ff",	--6816
		x"ff",	--6817
		x"ff",	--6818
		x"ff",	--6819
		x"ff",	--6820
		x"ff",	--6821
		x"ff",	--6822
		x"ff",	--6823
		x"ff",	--6824
		x"ff",	--6825
		x"ff",	--6826
		x"ff",	--6827
		x"ff",	--6828
		x"ff",	--6829
		x"ff",	--6830
		x"ff",	--6831
		x"ff",	--6832
		x"ff",	--6833
		x"ff",	--6834
		x"ff",	--6835
		x"ff",	--6836
		x"ff",	--6837
		x"ff",	--6838
		x"ff",	--6839
		x"ff",	--6840
		x"ff",	--6841
		x"ff",	--6842
		x"ff",	--6843
		x"ff",	--6844
		x"ff",	--6845
		x"ff",	--6846
		x"ff",	--6847
		x"ff",	--6848
		x"ff",	--6849
		x"ff",	--6850
		x"ff",	--6851
		x"ff",	--6852
		x"ff",	--6853
		x"ff",	--6854
		x"ff",	--6855
		x"ff",	--6856
		x"ff",	--6857
		x"ff",	--6858
		x"ff",	--6859
		x"ff",	--6860
		x"ff",	--6861
		x"ff",	--6862
		x"ff",	--6863
		x"ff",	--6864
		x"ff",	--6865
		x"ff",	--6866
		x"ff",	--6867
		x"ff",	--6868
		x"ff",	--6869
		x"ff",	--6870
		x"ff",	--6871
		x"ff",	--6872
		x"ff",	--6873
		x"ff",	--6874
		x"ff",	--6875
		x"ff",	--6876
		x"ff",	--6877
		x"ff",	--6878
		x"ff",	--6879
		x"ff",	--6880
		x"ff",	--6881
		x"ff",	--6882
		x"ff",	--6883
		x"ff",	--6884
		x"ff",	--6885
		x"ff",	--6886
		x"ff",	--6887
		x"ff",	--6888
		x"ff",	--6889
		x"ff",	--6890
		x"ff",	--6891
		x"ff",	--6892
		x"ff",	--6893
		x"ff",	--6894
		x"ff",	--6895
		x"ff",	--6896
		x"ff",	--6897
		x"ff",	--6898
		x"ff",	--6899
		x"ff",	--6900
		x"ff",	--6901
		x"ff",	--6902
		x"ff",	--6903
		x"ff",	--6904
		x"ff",	--6905
		x"ff",	--6906
		x"ff",	--6907
		x"ff",	--6908
		x"ff",	--6909
		x"ff",	--6910
		x"ff",	--6911
		x"ff",	--6912
		x"ff",	--6913
		x"ff",	--6914
		x"ff",	--6915
		x"ff",	--6916
		x"ff",	--6917
		x"ff",	--6918
		x"ff",	--6919
		x"ff",	--6920
		x"ff",	--6921
		x"ff",	--6922
		x"ff",	--6923
		x"ff",	--6924
		x"ff",	--6925
		x"ff",	--6926
		x"ff",	--6927
		x"ff",	--6928
		x"ff",	--6929
		x"ff",	--6930
		x"ff",	--6931
		x"ff",	--6932
		x"ff",	--6933
		x"ff",	--6934
		x"ff",	--6935
		x"ff",	--6936
		x"ff",	--6937
		x"ff",	--6938
		x"ff",	--6939
		x"ff",	--6940
		x"ff",	--6941
		x"ff",	--6942
		x"ff",	--6943
		x"ff",	--6944
		x"ff",	--6945
		x"ff",	--6946
		x"ff",	--6947
		x"ff",	--6948
		x"ff",	--6949
		x"ff",	--6950
		x"ff",	--6951
		x"ff",	--6952
		x"ff",	--6953
		x"ff",	--6954
		x"ff",	--6955
		x"ff",	--6956
		x"ff",	--6957
		x"ff",	--6958
		x"ff",	--6959
		x"ff",	--6960
		x"ff",	--6961
		x"ff",	--6962
		x"ff",	--6963
		x"ff",	--6964
		x"ff",	--6965
		x"ff",	--6966
		x"ff",	--6967
		x"ff",	--6968
		x"ff",	--6969
		x"ff",	--6970
		x"ff",	--6971
		x"ff",	--6972
		x"ff",	--6973
		x"ff",	--6974
		x"ff",	--6975
		x"ff",	--6976
		x"ff",	--6977
		x"ff",	--6978
		x"ff",	--6979
		x"ff",	--6980
		x"ff",	--6981
		x"ff",	--6982
		x"ff",	--6983
		x"ff",	--6984
		x"ff",	--6985
		x"ff",	--6986
		x"ff",	--6987
		x"ff",	--6988
		x"ff",	--6989
		x"ff",	--6990
		x"ff",	--6991
		x"ff",	--6992
		x"ff",	--6993
		x"ff",	--6994
		x"ff",	--6995
		x"ff",	--6996
		x"ff",	--6997
		x"ff",	--6998
		x"ff",	--6999
		x"ff",	--7000
		x"ff",	--7001
		x"ff",	--7002
		x"ff",	--7003
		x"ff",	--7004
		x"ff",	--7005
		x"ff",	--7006
		x"ff",	--7007
		x"ff",	--7008
		x"ff",	--7009
		x"ff",	--7010
		x"ff",	--7011
		x"ff",	--7012
		x"ff",	--7013
		x"ff",	--7014
		x"ff",	--7015
		x"ff",	--7016
		x"ff",	--7017
		x"ff",	--7018
		x"ff",	--7019
		x"ff",	--7020
		x"ff",	--7021
		x"ff",	--7022
		x"ff",	--7023
		x"ff",	--7024
		x"ff",	--7025
		x"ff",	--7026
		x"ff",	--7027
		x"ff",	--7028
		x"ff",	--7029
		x"ff",	--7030
		x"ff",	--7031
		x"ff",	--7032
		x"ff",	--7033
		x"ff",	--7034
		x"ff",	--7035
		x"ff",	--7036
		x"ff",	--7037
		x"ff",	--7038
		x"ff",	--7039
		x"ff",	--7040
		x"ff",	--7041
		x"ff",	--7042
		x"ff",	--7043
		x"ff",	--7044
		x"ff",	--7045
		x"ff",	--7046
		x"ff",	--7047
		x"ff",	--7048
		x"ff",	--7049
		x"ff",	--7050
		x"ff",	--7051
		x"ff",	--7052
		x"ff",	--7053
		x"ff",	--7054
		x"ff",	--7055
		x"ff",	--7056
		x"ff",	--7057
		x"ff",	--7058
		x"ff",	--7059
		x"ff",	--7060
		x"ff",	--7061
		x"ff",	--7062
		x"ff",	--7063
		x"ff",	--7064
		x"ff",	--7065
		x"ff",	--7066
		x"ff",	--7067
		x"ff",	--7068
		x"ff",	--7069
		x"ff",	--7070
		x"ff",	--7071
		x"ff",	--7072
		x"ff",	--7073
		x"ff",	--7074
		x"ff",	--7075
		x"ff",	--7076
		x"ff",	--7077
		x"ff",	--7078
		x"ff",	--7079
		x"ff",	--7080
		x"ff",	--7081
		x"ff",	--7082
		x"ff",	--7083
		x"ff",	--7084
		x"ff",	--7085
		x"ff",	--7086
		x"ff",	--7087
		x"ff",	--7088
		x"ff",	--7089
		x"ff",	--7090
		x"ff",	--7091
		x"ff",	--7092
		x"ff",	--7093
		x"ff",	--7094
		x"ff",	--7095
		x"ff",	--7096
		x"ff",	--7097
		x"ff",	--7098
		x"ff",	--7099
		x"ff",	--7100
		x"ff",	--7101
		x"ff",	--7102
		x"ff",	--7103
		x"ff",	--7104
		x"ff",	--7105
		x"ff",	--7106
		x"ff",	--7107
		x"ff",	--7108
		x"ff",	--7109
		x"ff",	--7110
		x"ff",	--7111
		x"ff",	--7112
		x"ff",	--7113
		x"ff",	--7114
		x"ff",	--7115
		x"ff",	--7116
		x"ff",	--7117
		x"ff",	--7118
		x"ff",	--7119
		x"ff",	--7120
		x"ff",	--7121
		x"ff",	--7122
		x"ff",	--7123
		x"ff",	--7124
		x"ff",	--7125
		x"ff",	--7126
		x"ff",	--7127
		x"ff",	--7128
		x"ff",	--7129
		x"ff",	--7130
		x"ff",	--7131
		x"ff",	--7132
		x"ff",	--7133
		x"ff",	--7134
		x"ff",	--7135
		x"ff",	--7136
		x"ff",	--7137
		x"ff",	--7138
		x"ff",	--7139
		x"ff",	--7140
		x"ff",	--7141
		x"ff",	--7142
		x"ff",	--7143
		x"ff",	--7144
		x"ff",	--7145
		x"ff",	--7146
		x"ff",	--7147
		x"ff",	--7148
		x"ff",	--7149
		x"ff",	--7150
		x"ff",	--7151
		x"ff",	--7152
		x"ff",	--7153
		x"ff",	--7154
		x"ff",	--7155
		x"ff",	--7156
		x"ff",	--7157
		x"ff",	--7158
		x"ff",	--7159
		x"ff",	--7160
		x"ff",	--7161
		x"ff",	--7162
		x"ff",	--7163
		x"ff",	--7164
		x"ff",	--7165
		x"ff",	--7166
		x"ff",	--7167
		x"ff",	--7168
		x"ff",	--7169
		x"ff",	--7170
		x"ff",	--7171
		x"ff",	--7172
		x"ff",	--7173
		x"ff",	--7174
		x"ff",	--7175
		x"ff",	--7176
		x"ff",	--7177
		x"ff",	--7178
		x"ff",	--7179
		x"ff",	--7180
		x"ff",	--7181
		x"ff",	--7182
		x"ff",	--7183
		x"ff",	--7184
		x"ff",	--7185
		x"ff",	--7186
		x"ff",	--7187
		x"ff",	--7188
		x"ff",	--7189
		x"ff",	--7190
		x"ff",	--7191
		x"ff",	--7192
		x"ff",	--7193
		x"ff",	--7194
		x"ff",	--7195
		x"ff",	--7196
		x"ff",	--7197
		x"ff",	--7198
		x"ff",	--7199
		x"ff",	--7200
		x"ff",	--7201
		x"ff",	--7202
		x"ff",	--7203
		x"ff",	--7204
		x"ff",	--7205
		x"ff",	--7206
		x"ff",	--7207
		x"ff",	--7208
		x"ff",	--7209
		x"ff",	--7210
		x"ff",	--7211
		x"ff",	--7212
		x"ff",	--7213
		x"ff",	--7214
		x"ff",	--7215
		x"ff",	--7216
		x"ff",	--7217
		x"ff",	--7218
		x"ff",	--7219
		x"ff",	--7220
		x"ff",	--7221
		x"ff",	--7222
		x"ff",	--7223
		x"ff",	--7224
		x"ff",	--7225
		x"ff",	--7226
		x"ff",	--7227
		x"ff",	--7228
		x"ff",	--7229
		x"ff",	--7230
		x"ff",	--7231
		x"ff",	--7232
		x"ff",	--7233
		x"ff",	--7234
		x"ff",	--7235
		x"ff",	--7236
		x"ff",	--7237
		x"ff",	--7238
		x"ff",	--7239
		x"ff",	--7240
		x"ff",	--7241
		x"ff",	--7242
		x"ff",	--7243
		x"ff",	--7244
		x"ff",	--7245
		x"ff",	--7246
		x"ff",	--7247
		x"ff",	--7248
		x"ff",	--7249
		x"ff",	--7250
		x"ff",	--7251
		x"ff",	--7252
		x"ff",	--7253
		x"ff",	--7254
		x"ff",	--7255
		x"ff",	--7256
		x"ff",	--7257
		x"ff",	--7258
		x"ff",	--7259
		x"ff",	--7260
		x"ff",	--7261
		x"ff",	--7262
		x"ff",	--7263
		x"ff",	--7264
		x"ff",	--7265
		x"ff",	--7266
		x"ff",	--7267
		x"ff",	--7268
		x"ff",	--7269
		x"ff",	--7270
		x"ff",	--7271
		x"ff",	--7272
		x"ff",	--7273
		x"ff",	--7274
		x"ff",	--7275
		x"ff",	--7276
		x"ff",	--7277
		x"ff",	--7278
		x"ff",	--7279
		x"ff",	--7280
		x"ff",	--7281
		x"ff",	--7282
		x"ff",	--7283
		x"ff",	--7284
		x"ff",	--7285
		x"ff",	--7286
		x"ff",	--7287
		x"ff",	--7288
		x"ff",	--7289
		x"ff",	--7290
		x"ff",	--7291
		x"ff",	--7292
		x"ff",	--7293
		x"ff",	--7294
		x"ff",	--7295
		x"ff",	--7296
		x"ff",	--7297
		x"ff",	--7298
		x"ff",	--7299
		x"ff",	--7300
		x"ff",	--7301
		x"ff",	--7302
		x"ff",	--7303
		x"ff",	--7304
		x"ff",	--7305
		x"ff",	--7306
		x"ff",	--7307
		x"ff",	--7308
		x"ff",	--7309
		x"ff",	--7310
		x"ff",	--7311
		x"ff",	--7312
		x"ff",	--7313
		x"ff",	--7314
		x"ff",	--7315
		x"ff",	--7316
		x"ff",	--7317
		x"ff",	--7318
		x"ff",	--7319
		x"ff",	--7320
		x"ff",	--7321
		x"ff",	--7322
		x"ff",	--7323
		x"ff",	--7324
		x"ff",	--7325
		x"ff",	--7326
		x"ff",	--7327
		x"ff",	--7328
		x"ff",	--7329
		x"ff",	--7330
		x"ff",	--7331
		x"ff",	--7332
		x"ff",	--7333
		x"ff",	--7334
		x"ff",	--7335
		x"ff",	--7336
		x"ff",	--7337
		x"ff",	--7338
		x"ff",	--7339
		x"ff",	--7340
		x"ff",	--7341
		x"ff",	--7342
		x"ff",	--7343
		x"ff",	--7344
		x"ff",	--7345
		x"ff",	--7346
		x"ff",	--7347
		x"ff",	--7348
		x"ff",	--7349
		x"ff",	--7350
		x"ff",	--7351
		x"ff",	--7352
		x"ff",	--7353
		x"ff",	--7354
		x"ff",	--7355
		x"ff",	--7356
		x"ff",	--7357
		x"ff",	--7358
		x"ff",	--7359
		x"ff",	--7360
		x"ff",	--7361
		x"ff",	--7362
		x"ff",	--7363
		x"ff",	--7364
		x"ff",	--7365
		x"ff",	--7366
		x"ff",	--7367
		x"ff",	--7368
		x"ff",	--7369
		x"ff",	--7370
		x"ff",	--7371
		x"ff",	--7372
		x"ff",	--7373
		x"ff",	--7374
		x"ff",	--7375
		x"ff",	--7376
		x"ff",	--7377
		x"ff",	--7378
		x"ff",	--7379
		x"ff",	--7380
		x"ff",	--7381
		x"ff",	--7382
		x"ff",	--7383
		x"ff",	--7384
		x"ff",	--7385
		x"ff",	--7386
		x"ff",	--7387
		x"ff",	--7388
		x"ff",	--7389
		x"ff",	--7390
		x"ff",	--7391
		x"ff",	--7392
		x"ff",	--7393
		x"ff",	--7394
		x"ff",	--7395
		x"ff",	--7396
		x"ff",	--7397
		x"ff",	--7398
		x"ff",	--7399
		x"ff",	--7400
		x"ff",	--7401
		x"ff",	--7402
		x"ff",	--7403
		x"ff",	--7404
		x"ff",	--7405
		x"ff",	--7406
		x"ff",	--7407
		x"ff",	--7408
		x"ff",	--7409
		x"ff",	--7410
		x"ff",	--7411
		x"ff",	--7412
		x"ff",	--7413
		x"ff",	--7414
		x"ff",	--7415
		x"ff",	--7416
		x"ff",	--7417
		x"ff",	--7418
		x"ff",	--7419
		x"ff",	--7420
		x"ff",	--7421
		x"ff",	--7422
		x"ff",	--7423
		x"ff",	--7424
		x"ff",	--7425
		x"ff",	--7426
		x"ff",	--7427
		x"ff",	--7428
		x"ff",	--7429
		x"ff",	--7430
		x"ff",	--7431
		x"ff",	--7432
		x"ff",	--7433
		x"ff",	--7434
		x"ff",	--7435
		x"ff",	--7436
		x"ff",	--7437
		x"ff",	--7438
		x"ff",	--7439
		x"ff",	--7440
		x"ff",	--7441
		x"ff",	--7442
		x"ff",	--7443
		x"ff",	--7444
		x"ff",	--7445
		x"ff",	--7446
		x"ff",	--7447
		x"ff",	--7448
		x"ff",	--7449
		x"ff",	--7450
		x"ff",	--7451
		x"ff",	--7452
		x"ff",	--7453
		x"ff",	--7454
		x"ff",	--7455
		x"ff",	--7456
		x"ff",	--7457
		x"ff",	--7458
		x"ff",	--7459
		x"ff",	--7460
		x"ff",	--7461
		x"ff",	--7462
		x"ff",	--7463
		x"ff",	--7464
		x"ff",	--7465
		x"ff",	--7466
		x"ff",	--7467
		x"ff",	--7468
		x"ff",	--7469
		x"ff",	--7470
		x"ff",	--7471
		x"ff",	--7472
		x"ff",	--7473
		x"ff",	--7474
		x"ff",	--7475
		x"ff",	--7476
		x"ff",	--7477
		x"ff",	--7478
		x"ff",	--7479
		x"ff",	--7480
		x"ff",	--7481
		x"ff",	--7482
		x"ff",	--7483
		x"ff",	--7484
		x"ff",	--7485
		x"ff",	--7486
		x"ff",	--7487
		x"ff",	--7488
		x"ff",	--7489
		x"ff",	--7490
		x"ff",	--7491
		x"ff",	--7492
		x"ff",	--7493
		x"ff",	--7494
		x"ff",	--7495
		x"ff",	--7496
		x"ff",	--7497
		x"ff",	--7498
		x"ff",	--7499
		x"ff",	--7500
		x"ff",	--7501
		x"ff",	--7502
		x"ff",	--7503
		x"ff",	--7504
		x"ff",	--7505
		x"ff",	--7506
		x"ff",	--7507
		x"ff",	--7508
		x"ff",	--7509
		x"ff",	--7510
		x"ff",	--7511
		x"ff",	--7512
		x"ff",	--7513
		x"ff",	--7514
		x"ff",	--7515
		x"ff",	--7516
		x"ff",	--7517
		x"ff",	--7518
		x"ff",	--7519
		x"ff",	--7520
		x"ff",	--7521
		x"ff",	--7522
		x"ff",	--7523
		x"ff",	--7524
		x"ff",	--7525
		x"ff",	--7526
		x"ff",	--7527
		x"ff",	--7528
		x"ff",	--7529
		x"ff",	--7530
		x"ff",	--7531
		x"ff",	--7532
		x"ff",	--7533
		x"ff",	--7534
		x"ff",	--7535
		x"ff",	--7536
		x"ff",	--7537
		x"ff",	--7538
		x"ff",	--7539
		x"ff",	--7540
		x"ff",	--7541
		x"ff",	--7542
		x"ff",	--7543
		x"ff",	--7544
		x"ff",	--7545
		x"ff",	--7546
		x"ff",	--7547
		x"ff",	--7548
		x"ff",	--7549
		x"ff",	--7550
		x"ff",	--7551
		x"ff",	--7552
		x"ff",	--7553
		x"ff",	--7554
		x"ff",	--7555
		x"ff",	--7556
		x"ff",	--7557
		x"ff",	--7558
		x"ff",	--7559
		x"ff",	--7560
		x"ff",	--7561
		x"ff",	--7562
		x"ff",	--7563
		x"ff",	--7564
		x"ff",	--7565
		x"ff",	--7566
		x"ff",	--7567
		x"ff",	--7568
		x"ff",	--7569
		x"ff",	--7570
		x"ff",	--7571
		x"ff",	--7572
		x"ff",	--7573
		x"ff",	--7574
		x"ff",	--7575
		x"ff",	--7576
		x"ff",	--7577
		x"ff",	--7578
		x"ff",	--7579
		x"ff",	--7580
		x"ff",	--7581
		x"ff",	--7582
		x"ff",	--7583
		x"ff",	--7584
		x"ff",	--7585
		x"ff",	--7586
		x"ff",	--7587
		x"ff",	--7588
		x"ff",	--7589
		x"ff",	--7590
		x"ff",	--7591
		x"ff",	--7592
		x"ff",	--7593
		x"ff",	--7594
		x"ff",	--7595
		x"ff",	--7596
		x"ff",	--7597
		x"ff",	--7598
		x"ff",	--7599
		x"ff",	--7600
		x"ff",	--7601
		x"ff",	--7602
		x"ff",	--7603
		x"ff",	--7604
		x"ff",	--7605
		x"ff",	--7606
		x"ff",	--7607
		x"ff",	--7608
		x"ff",	--7609
		x"ff",	--7610
		x"ff",	--7611
		x"ff",	--7612
		x"ff",	--7613
		x"ff",	--7614
		x"ff",	--7615
		x"ff",	--7616
		x"ff",	--7617
		x"ff",	--7618
		x"ff",	--7619
		x"ff",	--7620
		x"ff",	--7621
		x"ff",	--7622
		x"ff",	--7623
		x"ff",	--7624
		x"ff",	--7625
		x"ff",	--7626
		x"ff",	--7627
		x"ff",	--7628
		x"ff",	--7629
		x"ff",	--7630
		x"ff",	--7631
		x"ff",	--7632
		x"ff",	--7633
		x"ff",	--7634
		x"ff",	--7635
		x"ff",	--7636
		x"ff",	--7637
		x"ff",	--7638
		x"ff",	--7639
		x"ff",	--7640
		x"ff",	--7641
		x"ff",	--7642
		x"ff",	--7643
		x"ff",	--7644
		x"ff",	--7645
		x"ff",	--7646
		x"ff",	--7647
		x"ff",	--7648
		x"ff",	--7649
		x"ff",	--7650
		x"ff",	--7651
		x"ff",	--7652
		x"ff",	--7653
		x"ff",	--7654
		x"ff",	--7655
		x"ff",	--7656
		x"ff",	--7657
		x"ff",	--7658
		x"ff",	--7659
		x"ff",	--7660
		x"ff",	--7661
		x"ff",	--7662
		x"ff",	--7663
		x"ff",	--7664
		x"ff",	--7665
		x"ff",	--7666
		x"ff",	--7667
		x"ff",	--7668
		x"ff",	--7669
		x"ff",	--7670
		x"ff",	--7671
		x"ff",	--7672
		x"ff",	--7673
		x"ff",	--7674
		x"ff",	--7675
		x"ff",	--7676
		x"ff",	--7677
		x"ff",	--7678
		x"ff",	--7679
		x"ff",	--7680
		x"ff",	--7681
		x"ff",	--7682
		x"ff",	--7683
		x"ff",	--7684
		x"ff",	--7685
		x"ff",	--7686
		x"ff",	--7687
		x"ff",	--7688
		x"ff",	--7689
		x"ff",	--7690
		x"ff",	--7691
		x"ff",	--7692
		x"ff",	--7693
		x"ff",	--7694
		x"ff",	--7695
		x"ff",	--7696
		x"ff",	--7697
		x"ff",	--7698
		x"ff",	--7699
		x"ff",	--7700
		x"ff",	--7701
		x"ff",	--7702
		x"ff",	--7703
		x"ff",	--7704
		x"ff",	--7705
		x"ff",	--7706
		x"ff",	--7707
		x"ff",	--7708
		x"ff",	--7709
		x"ff",	--7710
		x"ff",	--7711
		x"ff",	--7712
		x"ff",	--7713
		x"ff",	--7714
		x"ff",	--7715
		x"ff",	--7716
		x"ff",	--7717
		x"ff",	--7718
		x"ff",	--7719
		x"ff",	--7720
		x"ff",	--7721
		x"ff",	--7722
		x"ff",	--7723
		x"ff",	--7724
		x"ff",	--7725
		x"ff",	--7726
		x"ff",	--7727
		x"ff",	--7728
		x"ff",	--7729
		x"ff",	--7730
		x"ff",	--7731
		x"ff",	--7732
		x"ff",	--7733
		x"ff",	--7734
		x"ff",	--7735
		x"ff",	--7736
		x"ff",	--7737
		x"ff",	--7738
		x"ff",	--7739
		x"ff",	--7740
		x"ff",	--7741
		x"ff",	--7742
		x"ff",	--7743
		x"ff",	--7744
		x"ff",	--7745
		x"ff",	--7746
		x"ff",	--7747
		x"ff",	--7748
		x"ff",	--7749
		x"ff",	--7750
		x"ff",	--7751
		x"ff",	--7752
		x"ff",	--7753
		x"ff",	--7754
		x"ff",	--7755
		x"ff",	--7756
		x"ff",	--7757
		x"ff",	--7758
		x"ff",	--7759
		x"ff",	--7760
		x"ff",	--7761
		x"ff",	--7762
		x"ff",	--7763
		x"ff",	--7764
		x"ff",	--7765
		x"ff",	--7766
		x"ff",	--7767
		x"ff",	--7768
		x"ff",	--7769
		x"ff",	--7770
		x"ff",	--7771
		x"ff",	--7772
		x"ff",	--7773
		x"ff",	--7774
		x"ff",	--7775
		x"ff",	--7776
		x"ff",	--7777
		x"ff",	--7778
		x"ff",	--7779
		x"ff",	--7780
		x"ff",	--7781
		x"ff",	--7782
		x"ff",	--7783
		x"ff",	--7784
		x"ff",	--7785
		x"ff",	--7786
		x"ff",	--7787
		x"ff",	--7788
		x"ff",	--7789
		x"ff",	--7790
		x"ff",	--7791
		x"ff",	--7792
		x"ff",	--7793
		x"ff",	--7794
		x"ff",	--7795
		x"ff",	--7796
		x"ff",	--7797
		x"ff",	--7798
		x"ff",	--7799
		x"ff",	--7800
		x"ff",	--7801
		x"ff",	--7802
		x"ff",	--7803
		x"ff",	--7804
		x"ff",	--7805
		x"ff",	--7806
		x"ff",	--7807
		x"ff",	--7808
		x"ff",	--7809
		x"ff",	--7810
		x"ff",	--7811
		x"ff",	--7812
		x"ff",	--7813
		x"ff",	--7814
		x"ff",	--7815
		x"ff",	--7816
		x"ff",	--7817
		x"ff",	--7818
		x"ff",	--7819
		x"ff",	--7820
		x"ff",	--7821
		x"ff",	--7822
		x"ff",	--7823
		x"ff",	--7824
		x"ff",	--7825
		x"ff",	--7826
		x"ff",	--7827
		x"ff",	--7828
		x"ff",	--7829
		x"ff",	--7830
		x"ff",	--7831
		x"ff",	--7832
		x"ff",	--7833
		x"ff",	--7834
		x"ff",	--7835
		x"ff",	--7836
		x"ff",	--7837
		x"ff",	--7838
		x"ff",	--7839
		x"ff",	--7840
		x"ff",	--7841
		x"ff",	--7842
		x"ff",	--7843
		x"ff",	--7844
		x"ff",	--7845
		x"ff",	--7846
		x"ff",	--7847
		x"ff",	--7848
		x"ff",	--7849
		x"ff",	--7850
		x"ff",	--7851
		x"ff",	--7852
		x"ff",	--7853
		x"ff",	--7854
		x"ff",	--7855
		x"ff",	--7856
		x"ff",	--7857
		x"ff",	--7858
		x"ff",	--7859
		x"ff",	--7860
		x"ff",	--7861
		x"ff",	--7862
		x"ff",	--7863
		x"ff",	--7864
		x"ff",	--7865
		x"ff",	--7866
		x"ff",	--7867
		x"ff",	--7868
		x"ff",	--7869
		x"ff",	--7870
		x"ff",	--7871
		x"ff",	--7872
		x"ff",	--7873
		x"ff",	--7874
		x"ff",	--7875
		x"ff",	--7876
		x"ff",	--7877
		x"ff",	--7878
		x"ff",	--7879
		x"ff",	--7880
		x"ff",	--7881
		x"ff",	--7882
		x"ff",	--7883
		x"ff",	--7884
		x"ff",	--7885
		x"ff",	--7886
		x"ff",	--7887
		x"ff",	--7888
		x"ff",	--7889
		x"ff",	--7890
		x"ff",	--7891
		x"ff",	--7892
		x"ff",	--7893
		x"ff",	--7894
		x"ff",	--7895
		x"ff",	--7896
		x"ff",	--7897
		x"ff",	--7898
		x"ff",	--7899
		x"ff",	--7900
		x"ff",	--7901
		x"ff",	--7902
		x"ff",	--7903
		x"ff",	--7904
		x"ff",	--7905
		x"ff",	--7906
		x"ff",	--7907
		x"ff",	--7908
		x"ff",	--7909
		x"ff",	--7910
		x"ff",	--7911
		x"ff",	--7912
		x"ff",	--7913
		x"ff",	--7914
		x"ff",	--7915
		x"ff",	--7916
		x"ff",	--7917
		x"ff",	--7918
		x"ff",	--7919
		x"ff",	--7920
		x"ff",	--7921
		x"ff",	--7922
		x"ff",	--7923
		x"ff",	--7924
		x"ff",	--7925
		x"ff",	--7926
		x"ff",	--7927
		x"ff",	--7928
		x"ff",	--7929
		x"ff",	--7930
		x"ff",	--7931
		x"ff",	--7932
		x"ff",	--7933
		x"ff",	--7934
		x"ff",	--7935
		x"ff",	--7936
		x"ff",	--7937
		x"ff",	--7938
		x"ff",	--7939
		x"ff",	--7940
		x"ff",	--7941
		x"ff",	--7942
		x"ff",	--7943
		x"ff",	--7944
		x"ff",	--7945
		x"ff",	--7946
		x"ff",	--7947
		x"ff",	--7948
		x"ff",	--7949
		x"ff",	--7950
		x"ff",	--7951
		x"ff",	--7952
		x"ff",	--7953
		x"ff",	--7954
		x"ff",	--7955
		x"ff",	--7956
		x"ff",	--7957
		x"ff",	--7958
		x"ff",	--7959
		x"ff",	--7960
		x"ff",	--7961
		x"ff",	--7962
		x"ff",	--7963
		x"ff",	--7964
		x"ff",	--7965
		x"ff",	--7966
		x"ff",	--7967
		x"ff",	--7968
		x"ff",	--7969
		x"ff",	--7970
		x"ff",	--7971
		x"ff",	--7972
		x"ff",	--7973
		x"ff",	--7974
		x"ff",	--7975
		x"ff",	--7976
		x"ff",	--7977
		x"ff",	--7978
		x"ff",	--7979
		x"ff",	--7980
		x"ff",	--7981
		x"ff",	--7982
		x"ff",	--7983
		x"ff",	--7984
		x"ff",	--7985
		x"ff",	--7986
		x"ff",	--7987
		x"ff",	--7988
		x"ff",	--7989
		x"ff",	--7990
		x"ff",	--7991
		x"ff",	--7992
		x"ff",	--7993
		x"ff",	--7994
		x"ff",	--7995
		x"ff",	--7996
		x"ff",	--7997
		x"ff",	--7998
		x"ff",	--7999
		x"ff",	--8000
		x"ff",	--8001
		x"ff",	--8002
		x"ff",	--8003
		x"ff",	--8004
		x"ff",	--8005
		x"ff",	--8006
		x"ff",	--8007
		x"ff",	--8008
		x"ff",	--8009
		x"ff",	--8010
		x"ff",	--8011
		x"ff",	--8012
		x"ff",	--8013
		x"ff",	--8014
		x"ff",	--8015
		x"ff",	--8016
		x"ff",	--8017
		x"ff",	--8018
		x"ff",	--8019
		x"ff",	--8020
		x"ff",	--8021
		x"ff",	--8022
		x"ff",	--8023
		x"ff",	--8024
		x"ff",	--8025
		x"ff",	--8026
		x"ff",	--8027
		x"ff",	--8028
		x"ff",	--8029
		x"ff",	--8030
		x"ff",	--8031
		x"ff",	--8032
		x"ff",	--8033
		x"ff",	--8034
		x"ff",	--8035
		x"ff",	--8036
		x"ff",	--8037
		x"ff",	--8038
		x"ff",	--8039
		x"ff",	--8040
		x"ff",	--8041
		x"ff",	--8042
		x"ff",	--8043
		x"ff",	--8044
		x"ff",	--8045
		x"ff",	--8046
		x"ff",	--8047
		x"ff",	--8048
		x"ff",	--8049
		x"ff",	--8050
		x"ff",	--8051
		x"ff",	--8052
		x"ff",	--8053
		x"ff",	--8054
		x"ff",	--8055
		x"ff",	--8056
		x"ff",	--8057
		x"ff",	--8058
		x"ff",	--8059
		x"ff",	--8060
		x"ff",	--8061
		x"ff",	--8062
		x"ff",	--8063
		x"ff",	--8064
		x"ff",	--8065
		x"ff",	--8066
		x"ff",	--8067
		x"ff",	--8068
		x"ff",	--8069
		x"ff",	--8070
		x"ff",	--8071
		x"ff",	--8072
		x"ff",	--8073
		x"ff",	--8074
		x"ff",	--8075
		x"ff",	--8076
		x"ff",	--8077
		x"ff",	--8078
		x"ff",	--8079
		x"ff",	--8080
		x"ff",	--8081
		x"ff",	--8082
		x"ff",	--8083
		x"ff",	--8084
		x"ff",	--8085
		x"ff",	--8086
		x"ff",	--8087
		x"ff",	--8088
		x"ff",	--8089
		x"ff",	--8090
		x"ff",	--8091
		x"ff",	--8092
		x"ff",	--8093
		x"ff",	--8094
		x"ff",	--8095
		x"ff",	--8096
		x"ff",	--8097
		x"ff",	--8098
		x"ff",	--8099
		x"ff",	--8100
		x"ff",	--8101
		x"ff",	--8102
		x"ff",	--8103
		x"ff",	--8104
		x"ff",	--8105
		x"ff",	--8106
		x"ff",	--8107
		x"ff",	--8108
		x"ff",	--8109
		x"ff",	--8110
		x"ff",	--8111
		x"ff",	--8112
		x"ff",	--8113
		x"ff",	--8114
		x"ff",	--8115
		x"ff",	--8116
		x"ff",	--8117
		x"ff",	--8118
		x"ff",	--8119
		x"ff",	--8120
		x"ff",	--8121
		x"ff",	--8122
		x"ff",	--8123
		x"ff",	--8124
		x"ff",	--8125
		x"ff",	--8126
		x"ff",	--8127
		x"ff",	--8128
		x"ff",	--8129
		x"ff",	--8130
		x"ff",	--8131
		x"ff",	--8132
		x"ff",	--8133
		x"ff",	--8134
		x"ff",	--8135
		x"ff",	--8136
		x"ff",	--8137
		x"ff",	--8138
		x"ff",	--8139
		x"ff",	--8140
		x"ff",	--8141
		x"ff",	--8142
		x"ff",	--8143
		x"ff",	--8144
		x"ff",	--8145
		x"ff",	--8146
		x"ff",	--8147
		x"ff",	--8148
		x"ff",	--8149
		x"ff",	--8150
		x"ff",	--8151
		x"ff",	--8152
		x"ff",	--8153
		x"ff",	--8154
		x"ff",	--8155
		x"ff",	--8156
		x"ff",	--8157
		x"ff",	--8158
		x"ff",	--8159
		x"ff",	--8160
		x"ff",	--8161
		x"ff",	--8162
		x"ff",	--8163
		x"ff",	--8164
		x"ff",	--8165
		x"ff",	--8166
		x"ff",	--8167
		x"ff",	--8168
		x"ff",	--8169
		x"ff",	--8170
		x"ff",	--8171
		x"ff",	--8172
		x"ff",	--8173
		x"ff",	--8174
		x"ff",	--8175
		x"c3",	--8176
		x"c3",	--8177
		x"c3",	--8178
		x"c3",	--8179
		x"c3",	--8180
		x"c3",	--8181
		x"c3",	--8182
		x"d4",	--8183
		x"d1",	--8184
		x"c3",	--8185
		x"c3",	--8186
		x"c3",	--8187
		x"c3",	--8188
		x"c3",	--8189
		x"c3",	--8190
		x"c0");	--8191

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
