library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"d0",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"06",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"d0",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"12",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"ca",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"d0",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"06",	--29
		x"f9",	--30
		x"31",	--31
		x"c2",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"80",	--41
		x"0f",	--42
		x"b0",	--43
		x"d8",	--44
		x"b0",	--45
		x"06",	--46
		x"c2",	--47
		x"19",	--48
		x"30",	--49
		x"63",	--50
		x"b0",	--51
		x"96",	--52
		x"21",	--53
		x"3d",	--54
		x"80",	--55
		x"3e",	--56
		x"a4",	--57
		x"7f",	--58
		x"77",	--59
		x"b0",	--60
		x"36",	--61
		x"3d",	--62
		x"86",	--63
		x"3e",	--64
		x"44",	--65
		x"7f",	--66
		x"72",	--67
		x"b0",	--68
		x"36",	--69
		x"3d",	--70
		x"8b",	--71
		x"3e",	--72
		x"f2",	--73
		x"7f",	--74
		x"70",	--75
		x"b0",	--76
		x"36",	--77
		x"3d",	--78
		x"8f",	--79
		x"3e",	--80
		x"bc",	--81
		x"7f",	--82
		x"62",	--83
		x"b0",	--84
		x"36",	--85
		x"0f",	--86
		x"b0",	--87
		x"cc",	--88
		x"2c",	--89
		x"3d",	--90
		x"20",	--91
		x"3e",	--92
		x"80",	--93
		x"0f",	--94
		x"3f",	--95
		x"0a",	--96
		x"b0",	--97
		x"dc",	--98
		x"0f",	--99
		x"3f",	--100
		x"0a",	--101
		x"b0",	--102
		x"24",	--103
		x"2c",	--104
		x"3d",	--105
		x"20",	--106
		x"3e",	--107
		x"88",	--108
		x"0f",	--109
		x"b0",	--110
		x"dc",	--111
		x"0f",	--112
		x"b0",	--113
		x"24",	--114
		x"0e",	--115
		x"0f",	--116
		x"3f",	--117
		x"0a",	--118
		x"b0",	--119
		x"e8",	--120
		x"f2",	--121
		x"80",	--122
		x"19",	--123
		x"32",	--124
		x"0b",	--125
		x"30",	--126
		x"9a",	--127
		x"b0",	--128
		x"96",	--129
		x"21",	--130
		x"0a",	--131
		x"32",	--132
		x"10",	--133
		x"1b",	--134
		x"3b",	--135
		x"09",	--136
		x"0a",	--137
		x"1f",	--138
		x"4e",	--139
		x"7e",	--140
		x"0f",	--141
		x"03",	--142
		x"0f",	--143
		x"7e",	--144
		x"fd",	--145
		x"4f",	--146
		x"02",	--147
		x"5f",	--148
		x"0b",	--149
		x"c2",	--150
		x"19",	--151
		x"b0",	--152
		x"e6",	--153
		x"0f",	--154
		x"e8",	--155
		x"b0",	--156
		x"0e",	--157
		x"7f",	--158
		x"1c",	--159
		x"7f",	--160
		x"0d",	--161
		x"22",	--162
		x"30",	--163
		x"9d",	--164
		x"b0",	--165
		x"96",	--166
		x"21",	--167
		x"3f",	--168
		x"14",	--169
		x"0f",	--170
		x"0a",	--171
		x"ca",	--172
		x"00",	--173
		x"0f",	--174
		x"30",	--175
		x"a0",	--176
		x"b0",	--177
		x"96",	--178
		x"21",	--179
		x"0e",	--180
		x"3e",	--181
		x"14",	--182
		x"5f",	--183
		x"14",	--184
		x"b0",	--185
		x"6a",	--186
		x"c2",	--187
		x"0a",	--188
		x"c6",	--189
		x"3a",	--190
		x"30",	--191
		x"a6",	--192
		x"b0",	--193
		x"96",	--194
		x"21",	--195
		x"bf",	--196
		x"3a",	--197
		x"28",	--198
		x"bc",	--199
		x"4e",	--200
		x"8e",	--201
		x"0e",	--202
		x"30",	--203
		x"aa",	--204
		x"81",	--205
		x"40",	--206
		x"b0",	--207
		x"96",	--208
		x"21",	--209
		x"3e",	--210
		x"14",	--211
		x"0e",	--212
		x"0e",	--213
		x"1f",	--214
		x"3c",	--215
		x"ce",	--216
		x"00",	--217
		x"1a",	--218
		x"a8",	--219
		x"30",	--220
		x"e2",	--221
		x"b2",	--222
		x"00",	--223
		x"92",	--224
		x"a2",	--225
		x"94",	--226
		x"b2",	--227
		x"6d",	--228
		x"96",	--229
		x"30",	--230
		x"ea",	--231
		x"b0",	--232
		x"96",	--233
		x"92",	--234
		x"90",	--235
		x"b1",	--236
		x"08",	--237
		x"00",	--238
		x"b0",	--239
		x"96",	--240
		x"21",	--241
		x"0f",	--242
		x"30",	--243
		x"82",	--244
		x"0e",	--245
		x"82",	--246
		x"0c",	--247
		x"30",	--248
		x"31",	--249
		x"ff",	--250
		x"20",	--251
		x"01",	--252
		x"39",	--253
		x"cf",	--254
		x"02",	--255
		x"36",	--256
		x"0d",	--257
		x"0e",	--258
		x"2e",	--259
		x"0f",	--260
		x"2f",	--261
		x"b0",	--262
		x"c2",	--263
		x"81",	--264
		x"00",	--265
		x"40",	--266
		x"0d",	--267
		x"0e",	--268
		x"0f",	--269
		x"2f",	--270
		x"b0",	--271
		x"c2",	--272
		x"81",	--273
		x"00",	--274
		x"37",	--275
		x"1e",	--276
		x"04",	--277
		x"0f",	--278
		x"b0",	--279
		x"00",	--280
		x"0c",	--281
		x"3d",	--282
		x"c8",	--283
		x"b0",	--284
		x"d0",	--285
		x"0d",	--286
		x"0e",	--287
		x"1f",	--288
		x"0e",	--289
		x"b0",	--290
		x"78",	--291
		x"1e",	--292
		x"02",	--293
		x"0f",	--294
		x"b0",	--295
		x"00",	--296
		x"0c",	--297
		x"3d",	--298
		x"c8",	--299
		x"b0",	--300
		x"d0",	--301
		x"0d",	--302
		x"0e",	--303
		x"1f",	--304
		x"0c",	--305
		x"b0",	--306
		x"78",	--307
		x"0f",	--308
		x"31",	--309
		x"30",	--310
		x"30",	--311
		x"21",	--312
		x"81",	--313
		x"08",	--314
		x"b0",	--315
		x"96",	--316
		x"1f",	--317
		x"08",	--318
		x"6f",	--319
		x"8f",	--320
		x"81",	--321
		x"00",	--322
		x"30",	--323
		x"32",	--324
		x"b0",	--325
		x"96",	--326
		x"21",	--327
		x"3f",	--328
		x"31",	--329
		x"30",	--330
		x"30",	--331
		x"43",	--332
		x"b0",	--333
		x"96",	--334
		x"21",	--335
		x"3f",	--336
		x"e3",	--337
		x"0b",	--338
		x"31",	--339
		x"fa",	--340
		x"0b",	--341
		x"30",	--342
		x"ad",	--343
		x"b0",	--344
		x"96",	--345
		x"21",	--346
		x"fb",	--347
		x"20",	--348
		x"01",	--349
		x"2a",	--350
		x"cb",	--351
		x"02",	--352
		x"27",	--353
		x"0d",	--354
		x"0e",	--355
		x"2e",	--356
		x"0f",	--357
		x"2f",	--358
		x"b0",	--359
		x"c2",	--360
		x"81",	--361
		x"00",	--362
		x"2f",	--363
		x"0d",	--364
		x"0e",	--365
		x"0f",	--366
		x"2f",	--367
		x"b0",	--368
		x"c2",	--369
		x"81",	--370
		x"00",	--371
		x"26",	--372
		x"11",	--373
		x"04",	--374
		x"11",	--375
		x"08",	--376
		x"30",	--377
		x"fb",	--378
		x"b0",	--379
		x"96",	--380
		x"31",	--381
		x"06",	--382
		x"1f",	--383
		x"04",	--384
		x"9f",	--385
		x"02",	--386
		x"00",	--387
		x"0f",	--388
		x"31",	--389
		x"06",	--390
		x"3b",	--391
		x"30",	--392
		x"30",	--393
		x"b5",	--394
		x"b0",	--395
		x"96",	--396
		x"6f",	--397
		x"8f",	--398
		x"81",	--399
		x"00",	--400
		x"30",	--401
		x"c6",	--402
		x"b0",	--403
		x"96",	--404
		x"21",	--405
		x"3f",	--406
		x"31",	--407
		x"06",	--408
		x"3b",	--409
		x"30",	--410
		x"30",	--411
		x"db",	--412
		x"b0",	--413
		x"96",	--414
		x"21",	--415
		x"3f",	--416
		x"e3",	--417
		x"0b",	--418
		x"21",	--419
		x"0b",	--420
		x"30",	--421
		x"07",	--422
		x"b0",	--423
		x"96",	--424
		x"21",	--425
		x"fb",	--426
		x"20",	--427
		x"01",	--428
		x"1b",	--429
		x"cb",	--430
		x"02",	--431
		x"18",	--432
		x"0d",	--433
		x"0e",	--434
		x"2e",	--435
		x"0f",	--436
		x"2f",	--437
		x"b0",	--438
		x"c2",	--439
		x"81",	--440
		x"00",	--441
		x"1f",	--442
		x"1f",	--443
		x"02",	--444
		x"2f",	--445
		x"0f",	--446
		x"30",	--447
		x"fb",	--448
		x"b0",	--449
		x"96",	--450
		x"31",	--451
		x"06",	--452
		x"0f",	--453
		x"21",	--454
		x"3b",	--455
		x"30",	--456
		x"30",	--457
		x"b5",	--458
		x"b0",	--459
		x"96",	--460
		x"6f",	--461
		x"8f",	--462
		x"81",	--463
		x"00",	--464
		x"30",	--465
		x"0e",	--466
		x"b0",	--467
		x"96",	--468
		x"21",	--469
		x"3f",	--470
		x"21",	--471
		x"3b",	--472
		x"30",	--473
		x"30",	--474
		x"db",	--475
		x"b0",	--476
		x"96",	--477
		x"21",	--478
		x"3f",	--479
		x"e5",	--480
		x"0b",	--481
		x"0a",	--482
		x"09",	--483
		x"08",	--484
		x"07",	--485
		x"8f",	--486
		x"00",	--487
		x"8d",	--488
		x"00",	--489
		x"6c",	--490
		x"4c",	--491
		x"5f",	--492
		x"0b",	--493
		x"1b",	--494
		x"08",	--495
		x"0a",	--496
		x"07",	--497
		x"09",	--498
		x"18",	--499
		x"7a",	--500
		x"0a",	--501
		x"35",	--502
		x"2c",	--503
		x"0c",	--504
		x"0c",	--505
		x"0c",	--506
		x"0c",	--507
		x"8f",	--508
		x"00",	--509
		x"3c",	--510
		x"d0",	--511
		x"6a",	--512
		x"8a",	--513
		x"0c",	--514
		x"8f",	--515
		x"00",	--516
		x"17",	--517
		x"19",	--518
		x"0a",	--519
		x"08",	--520
		x"7c",	--521
		x"4c",	--522
		x"40",	--523
		x"7c",	--524
		x"78",	--525
		x"1b",	--526
		x"7c",	--527
		x"20",	--528
		x"43",	--529
		x"4a",	--530
		x"7a",	--531
		x"d0",	--532
		x"07",	--533
		x"dd",	--534
		x"7a",	--535
		x"0a",	--536
		x"46",	--537
		x"2a",	--538
		x"0a",	--539
		x"0c",	--540
		x"0c",	--541
		x"0c",	--542
		x"0c",	--543
		x"8f",	--544
		x"00",	--545
		x"3c",	--546
		x"d0",	--547
		x"68",	--548
		x"88",	--549
		x"0c",	--550
		x"8f",	--551
		x"00",	--552
		x"dc",	--553
		x"17",	--554
		x"da",	--555
		x"4a",	--556
		x"7a",	--557
		x"9f",	--558
		x"7a",	--559
		x"06",	--560
		x"0a",	--561
		x"2c",	--562
		x"0c",	--563
		x"0c",	--564
		x"0c",	--565
		x"0c",	--566
		x"8f",	--567
		x"00",	--568
		x"3c",	--569
		x"a9",	--570
		x"c4",	--571
		x"4a",	--572
		x"7a",	--573
		x"bf",	--574
		x"7a",	--575
		x"06",	--576
		x"1e",	--577
		x"2c",	--578
		x"0c",	--579
		x"0c",	--580
		x"0c",	--581
		x"0c",	--582
		x"8f",	--583
		x"00",	--584
		x"3c",	--585
		x"c9",	--586
		x"b4",	--587
		x"9d",	--588
		x"00",	--589
		x"0f",	--590
		x"37",	--591
		x"38",	--592
		x"39",	--593
		x"3a",	--594
		x"3b",	--595
		x"30",	--596
		x"9d",	--597
		x"00",	--598
		x"0f",	--599
		x"1f",	--600
		x"0f",	--601
		x"37",	--602
		x"38",	--603
		x"39",	--604
		x"3a",	--605
		x"3b",	--606
		x"30",	--607
		x"8c",	--608
		x"0c",	--609
		x"30",	--610
		x"1d",	--611
		x"b0",	--612
		x"96",	--613
		x"21",	--614
		x"0f",	--615
		x"37",	--616
		x"38",	--617
		x"39",	--618
		x"3a",	--619
		x"3b",	--620
		x"30",	--621
		x"0b",	--622
		x"0a",	--623
		x"0b",	--624
		x"0a",	--625
		x"8f",	--626
		x"00",	--627
		x"8f",	--628
		x"02",	--629
		x"8f",	--630
		x"04",	--631
		x"0c",	--632
		x"0d",	--633
		x"3e",	--634
		x"00",	--635
		x"3f",	--636
		x"6e",	--637
		x"b0",	--638
		x"34",	--639
		x"8b",	--640
		x"02",	--641
		x"02",	--642
		x"32",	--643
		x"03",	--644
		x"82",	--645
		x"32",	--646
		x"b2",	--647
		x"18",	--648
		x"38",	--649
		x"9b",	--650
		x"3a",	--651
		x"06",	--652
		x"32",	--653
		x"0f",	--654
		x"3a",	--655
		x"3b",	--656
		x"30",	--657
		x"0b",	--658
		x"09",	--659
		x"08",	--660
		x"8f",	--661
		x"06",	--662
		x"bf",	--663
		x"00",	--664
		x"08",	--665
		x"2b",	--666
		x"1e",	--667
		x"02",	--668
		x"0f",	--669
		x"b0",	--670
		x"00",	--671
		x"0c",	--672
		x"3d",	--673
		x"00",	--674
		x"b0",	--675
		x"ac",	--676
		x"08",	--677
		x"09",	--678
		x"1e",	--679
		x"06",	--680
		x"0f",	--681
		x"b0",	--682
		x"00",	--683
		x"0c",	--684
		x"0d",	--685
		x"0e",	--686
		x"0f",	--687
		x"b0",	--688
		x"5c",	--689
		x"b0",	--690
		x"3c",	--691
		x"8b",	--692
		x"04",	--693
		x"9b",	--694
		x"00",	--695
		x"38",	--696
		x"39",	--697
		x"3b",	--698
		x"30",	--699
		x"0b",	--700
		x"0a",	--701
		x"09",	--702
		x"0a",	--703
		x"0b",	--704
		x"8f",	--705
		x"06",	--706
		x"8f",	--707
		x"08",	--708
		x"29",	--709
		x"1e",	--710
		x"02",	--711
		x"0f",	--712
		x"b0",	--713
		x"00",	--714
		x"0c",	--715
		x"0d",	--716
		x"0e",	--717
		x"0f",	--718
		x"b0",	--719
		x"ac",	--720
		x"0a",	--721
		x"0b",	--722
		x"1e",	--723
		x"06",	--724
		x"0f",	--725
		x"b0",	--726
		x"00",	--727
		x"0c",	--728
		x"0d",	--729
		x"0e",	--730
		x"0f",	--731
		x"b0",	--732
		x"5c",	--733
		x"b0",	--734
		x"3c",	--735
		x"89",	--736
		x"04",	--737
		x"39",	--738
		x"3a",	--739
		x"3b",	--740
		x"30",	--741
		x"0b",	--742
		x"0a",	--743
		x"92",	--744
		x"06",	--745
		x"14",	--746
		x"3b",	--747
		x"14",	--748
		x"0a",	--749
		x"2b",	--750
		x"5f",	--751
		x"fc",	--752
		x"8f",	--753
		x"0f",	--754
		x"30",	--755
		x"32",	--756
		x"b0",	--757
		x"96",	--758
		x"31",	--759
		x"06",	--760
		x"1a",	--761
		x"3b",	--762
		x"06",	--763
		x"1a",	--764
		x"06",	--765
		x"ef",	--766
		x"0f",	--767
		x"3a",	--768
		x"3b",	--769
		x"30",	--770
		x"1e",	--771
		x"06",	--772
		x"3e",	--773
		x"40",	--774
		x"12",	--775
		x"0f",	--776
		x"0f",	--777
		x"0f",	--778
		x"0f",	--779
		x"3f",	--780
		x"10",	--781
		x"ff",	--782
		x"68",	--783
		x"00",	--784
		x"bf",	--785
		x"cc",	--786
		x"02",	--787
		x"bf",	--788
		x"00",	--789
		x"04",	--790
		x"1e",	--791
		x"82",	--792
		x"06",	--793
		x"30",	--794
		x"0b",	--795
		x"1b",	--796
		x"06",	--797
		x"3b",	--798
		x"40",	--799
		x"12",	--800
		x"0c",	--801
		x"0c",	--802
		x"0c",	--803
		x"0c",	--804
		x"3c",	--805
		x"10",	--806
		x"cc",	--807
		x"00",	--808
		x"8c",	--809
		x"02",	--810
		x"8c",	--811
		x"04",	--812
		x"1b",	--813
		x"82",	--814
		x"06",	--815
		x"0f",	--816
		x"3b",	--817
		x"30",	--818
		x"3f",	--819
		x"fc",	--820
		x"0b",	--821
		x"1b",	--822
		x"06",	--823
		x"1b",	--824
		x"0f",	--825
		x"5f",	--826
		x"10",	--827
		x"14",	--828
		x"3d",	--829
		x"16",	--830
		x"0c",	--831
		x"05",	--832
		x"3d",	--833
		x"06",	--834
		x"cd",	--835
		x"fa",	--836
		x"0c",	--837
		x"1c",	--838
		x"0c",	--839
		x"f8",	--840
		x"30",	--841
		x"3a",	--842
		x"b0",	--843
		x"96",	--844
		x"21",	--845
		x"3f",	--846
		x"3b",	--847
		x"30",	--848
		x"0c",	--849
		x"0d",	--850
		x"0d",	--851
		x"0c",	--852
		x"0c",	--853
		x"3c",	--854
		x"10",	--855
		x"0f",	--856
		x"9c",	--857
		x"02",	--858
		x"3b",	--859
		x"30",	--860
		x"5e",	--861
		x"81",	--862
		x"3e",	--863
		x"fc",	--864
		x"c2",	--865
		x"84",	--866
		x"0f",	--867
		x"30",	--868
		x"3f",	--869
		x"0f",	--870
		x"5f",	--871
		x"f8",	--872
		x"8f",	--873
		x"b0",	--874
		x"ba",	--875
		x"30",	--876
		x"0b",	--877
		x"0b",	--878
		x"0e",	--879
		x"0e",	--880
		x"0e",	--881
		x"0e",	--882
		x"0e",	--883
		x"0f",	--884
		x"b0",	--885
		x"ca",	--886
		x"0f",	--887
		x"b0",	--888
		x"ca",	--889
		x"3b",	--890
		x"30",	--891
		x"0b",	--892
		x"0a",	--893
		x"0a",	--894
		x"3b",	--895
		x"07",	--896
		x"0e",	--897
		x"4d",	--898
		x"7d",	--899
		x"0f",	--900
		x"03",	--901
		x"0e",	--902
		x"7d",	--903
		x"fd",	--904
		x"1e",	--905
		x"0a",	--906
		x"3f",	--907
		x"31",	--908
		x"b0",	--909
		x"ba",	--910
		x"3b",	--911
		x"3b",	--912
		x"ef",	--913
		x"3a",	--914
		x"3b",	--915
		x"30",	--916
		x"3f",	--917
		x"30",	--918
		x"f5",	--919
		x"0b",	--920
		x"0b",	--921
		x"0e",	--922
		x"8e",	--923
		x"8e",	--924
		x"0f",	--925
		x"b0",	--926
		x"da",	--927
		x"0f",	--928
		x"b0",	--929
		x"da",	--930
		x"3b",	--931
		x"30",	--932
		x"0b",	--933
		x"0a",	--934
		x"0a",	--935
		x"0b",	--936
		x"0d",	--937
		x"8d",	--938
		x"8d",	--939
		x"0f",	--940
		x"b0",	--941
		x"da",	--942
		x"0f",	--943
		x"b0",	--944
		x"da",	--945
		x"0c",	--946
		x"0d",	--947
		x"8d",	--948
		x"8c",	--949
		x"4d",	--950
		x"0d",	--951
		x"0f",	--952
		x"b0",	--953
		x"da",	--954
		x"0f",	--955
		x"b0",	--956
		x"da",	--957
		x"3a",	--958
		x"3b",	--959
		x"30",	--960
		x"0b",	--961
		x"0a",	--962
		x"09",	--963
		x"0a",	--964
		x"0e",	--965
		x"19",	--966
		x"09",	--967
		x"39",	--968
		x"0b",	--969
		x"0d",	--970
		x"0d",	--971
		x"6f",	--972
		x"8f",	--973
		x"b0",	--974
		x"da",	--975
		x"0b",	--976
		x"0e",	--977
		x"1b",	--978
		x"3b",	--979
		x"07",	--980
		x"05",	--981
		x"3f",	--982
		x"20",	--983
		x"b0",	--984
		x"ba",	--985
		x"ef",	--986
		x"3f",	--987
		x"3a",	--988
		x"b0",	--989
		x"ba",	--990
		x"ea",	--991
		x"39",	--992
		x"3a",	--993
		x"3b",	--994
		x"30",	--995
		x"0b",	--996
		x"0a",	--997
		x"09",	--998
		x"0a",	--999
		x"0e",	--1000
		x"17",	--1001
		x"09",	--1002
		x"39",	--1003
		x"0b",	--1004
		x"6f",	--1005
		x"8f",	--1006
		x"b0",	--1007
		x"ca",	--1008
		x"0b",	--1009
		x"0e",	--1010
		x"1b",	--1011
		x"3b",	--1012
		x"07",	--1013
		x"f6",	--1014
		x"3f",	--1015
		x"20",	--1016
		x"b0",	--1017
		x"ba",	--1018
		x"6f",	--1019
		x"8f",	--1020
		x"b0",	--1021
		x"ca",	--1022
		x"0b",	--1023
		x"f2",	--1024
		x"39",	--1025
		x"3a",	--1026
		x"3b",	--1027
		x"30",	--1028
		x"0b",	--1029
		x"0a",	--1030
		x"09",	--1031
		x"31",	--1032
		x"ec",	--1033
		x"0b",	--1034
		x"0f",	--1035
		x"34",	--1036
		x"3b",	--1037
		x"0a",	--1038
		x"38",	--1039
		x"09",	--1040
		x"0a",	--1041
		x"0a",	--1042
		x"3e",	--1043
		x"0a",	--1044
		x"0f",	--1045
		x"b0",	--1046
		x"2c",	--1047
		x"7f",	--1048
		x"30",	--1049
		x"ca",	--1050
		x"00",	--1051
		x"19",	--1052
		x"3e",	--1053
		x"0a",	--1054
		x"0f",	--1055
		x"b0",	--1056
		x"fa",	--1057
		x"0b",	--1058
		x"3f",	--1059
		x"0a",	--1060
		x"eb",	--1061
		x"0a",	--1062
		x"1a",	--1063
		x"09",	--1064
		x"3e",	--1065
		x"0a",	--1066
		x"0f",	--1067
		x"b0",	--1068
		x"2c",	--1069
		x"7f",	--1070
		x"30",	--1071
		x"c9",	--1072
		x"00",	--1073
		x"3a",	--1074
		x"0f",	--1075
		x"0f",	--1076
		x"6f",	--1077
		x"8f",	--1078
		x"b0",	--1079
		x"ba",	--1080
		x"0a",	--1081
		x"f7",	--1082
		x"31",	--1083
		x"14",	--1084
		x"39",	--1085
		x"3a",	--1086
		x"3b",	--1087
		x"30",	--1088
		x"3f",	--1089
		x"2d",	--1090
		x"b0",	--1091
		x"ba",	--1092
		x"3b",	--1093
		x"1b",	--1094
		x"c5",	--1095
		x"1a",	--1096
		x"09",	--1097
		x"dd",	--1098
		x"0b",	--1099
		x"0a",	--1100
		x"09",	--1101
		x"0b",	--1102
		x"3b",	--1103
		x"39",	--1104
		x"6f",	--1105
		x"4f",	--1106
		x"0b",	--1107
		x"1a",	--1108
		x"8f",	--1109
		x"b0",	--1110
		x"ba",	--1111
		x"0a",	--1112
		x"09",	--1113
		x"19",	--1114
		x"5f",	--1115
		x"01",	--1116
		x"4f",	--1117
		x"10",	--1118
		x"7f",	--1119
		x"25",	--1120
		x"f3",	--1121
		x"0a",	--1122
		x"1a",	--1123
		x"5f",	--1124
		x"01",	--1125
		x"7f",	--1126
		x"db",	--1127
		x"7f",	--1128
		x"54",	--1129
		x"ee",	--1130
		x"4f",	--1131
		x"0f",	--1132
		x"10",	--1133
		x"50",	--1134
		x"39",	--1135
		x"3a",	--1136
		x"3b",	--1137
		x"30",	--1138
		x"09",	--1139
		x"29",	--1140
		x"1e",	--1141
		x"02",	--1142
		x"2f",	--1143
		x"b0",	--1144
		x"82",	--1145
		x"0b",	--1146
		x"dd",	--1147
		x"09",	--1148
		x"29",	--1149
		x"2f",	--1150
		x"b0",	--1151
		x"30",	--1152
		x"0b",	--1153
		x"d6",	--1154
		x"0f",	--1155
		x"2b",	--1156
		x"29",	--1157
		x"6f",	--1158
		x"4f",	--1159
		x"d0",	--1160
		x"19",	--1161
		x"8f",	--1162
		x"b0",	--1163
		x"ba",	--1164
		x"7f",	--1165
		x"4f",	--1166
		x"fa",	--1167
		x"c8",	--1168
		x"09",	--1169
		x"29",	--1170
		x"1e",	--1171
		x"02",	--1172
		x"2f",	--1173
		x"b0",	--1174
		x"c8",	--1175
		x"0b",	--1176
		x"bf",	--1177
		x"09",	--1178
		x"29",	--1179
		x"2e",	--1180
		x"0f",	--1181
		x"8f",	--1182
		x"8f",	--1183
		x"8f",	--1184
		x"8f",	--1185
		x"b0",	--1186
		x"4a",	--1187
		x"0b",	--1188
		x"b3",	--1189
		x"09",	--1190
		x"29",	--1191
		x"2f",	--1192
		x"b0",	--1193
		x"0a",	--1194
		x"0b",	--1195
		x"ac",	--1196
		x"09",	--1197
		x"29",	--1198
		x"2f",	--1199
		x"b0",	--1200
		x"ba",	--1201
		x"0b",	--1202
		x"a5",	--1203
		x"09",	--1204
		x"29",	--1205
		x"2f",	--1206
		x"b0",	--1207
		x"da",	--1208
		x"0b",	--1209
		x"9e",	--1210
		x"09",	--1211
		x"29",	--1212
		x"2f",	--1213
		x"b0",	--1214
		x"f8",	--1215
		x"0b",	--1216
		x"97",	--1217
		x"3f",	--1218
		x"25",	--1219
		x"b0",	--1220
		x"ba",	--1221
		x"92",	--1222
		x"0f",	--1223
		x"0e",	--1224
		x"1f",	--1225
		x"08",	--1226
		x"df",	--1227
		x"85",	--1228
		x"90",	--1229
		x"1f",	--1230
		x"08",	--1231
		x"3f",	--1232
		x"3f",	--1233
		x"16",	--1234
		x"92",	--1235
		x"08",	--1236
		x"1e",	--1237
		x"08",	--1238
		x"1f",	--1239
		x"0a",	--1240
		x"0e",	--1241
		x"02",	--1242
		x"92",	--1243
		x"0a",	--1244
		x"f2",	--1245
		x"10",	--1246
		x"81",	--1247
		x"b1",	--1248
		x"10",	--1249
		x"04",	--1250
		x"3e",	--1251
		x"3f",	--1252
		x"b1",	--1253
		x"f0",	--1254
		x"00",	--1255
		x"00",	--1256
		x"82",	--1257
		x"08",	--1258
		x"e9",	--1259
		x"b2",	--1260
		x"c3",	--1261
		x"82",	--1262
		x"f2",	--1263
		x"11",	--1264
		x"80",	--1265
		x"30",	--1266
		x"1e",	--1267
		x"08",	--1268
		x"1f",	--1269
		x"0a",	--1270
		x"0e",	--1271
		x"05",	--1272
		x"1f",	--1273
		x"08",	--1274
		x"1f",	--1275
		x"0a",	--1276
		x"30",	--1277
		x"1d",	--1278
		x"08",	--1279
		x"1e",	--1280
		x"0a",	--1281
		x"3f",	--1282
		x"40",	--1283
		x"0f",	--1284
		x"0f",	--1285
		x"30",	--1286
		x"1f",	--1287
		x"0a",	--1288
		x"5f",	--1289
		x"90",	--1290
		x"1d",	--1291
		x"0a",	--1292
		x"1e",	--1293
		x"08",	--1294
		x"0d",	--1295
		x"0b",	--1296
		x"1e",	--1297
		x"0a",	--1298
		x"3e",	--1299
		x"3f",	--1300
		x"03",	--1301
		x"82",	--1302
		x"0a",	--1303
		x"30",	--1304
		x"92",	--1305
		x"0a",	--1306
		x"30",	--1307
		x"4f",	--1308
		x"30",	--1309
		x"0b",	--1310
		x"0a",	--1311
		x"0a",	--1312
		x"0b",	--1313
		x"0c",	--1314
		x"3d",	--1315
		x"00",	--1316
		x"b0",	--1317
		x"20",	--1318
		x"0f",	--1319
		x"07",	--1320
		x"0e",	--1321
		x"0f",	--1322
		x"b0",	--1323
		x"70",	--1324
		x"3a",	--1325
		x"3b",	--1326
		x"30",	--1327
		x"0c",	--1328
		x"3d",	--1329
		x"00",	--1330
		x"0e",	--1331
		x"0f",	--1332
		x"b0",	--1333
		x"5c",	--1334
		x"b0",	--1335
		x"70",	--1336
		x"0e",	--1337
		x"3f",	--1338
		x"00",	--1339
		x"3a",	--1340
		x"3b",	--1341
		x"30",	--1342
		x"0b",	--1343
		x"0a",	--1344
		x"09",	--1345
		x"08",	--1346
		x"07",	--1347
		x"06",	--1348
		x"05",	--1349
		x"04",	--1350
		x"31",	--1351
		x"fa",	--1352
		x"08",	--1353
		x"6b",	--1354
		x"6b",	--1355
		x"67",	--1356
		x"6c",	--1357
		x"6c",	--1358
		x"e9",	--1359
		x"6b",	--1360
		x"02",	--1361
		x"30",	--1362
		x"fe",	--1363
		x"6c",	--1364
		x"e3",	--1365
		x"6c",	--1366
		x"bb",	--1367
		x"6b",	--1368
		x"df",	--1369
		x"91",	--1370
		x"02",	--1371
		x"00",	--1372
		x"1b",	--1373
		x"02",	--1374
		x"14",	--1375
		x"04",	--1376
		x"15",	--1377
		x"06",	--1378
		x"16",	--1379
		x"04",	--1380
		x"17",	--1381
		x"06",	--1382
		x"2c",	--1383
		x"0c",	--1384
		x"09",	--1385
		x"0c",	--1386
		x"bf",	--1387
		x"39",	--1388
		x"20",	--1389
		x"50",	--1390
		x"1c",	--1391
		x"d7",	--1392
		x"81",	--1393
		x"02",	--1394
		x"81",	--1395
		x"04",	--1396
		x"4c",	--1397
		x"7c",	--1398
		x"1f",	--1399
		x"0b",	--1400
		x"0a",	--1401
		x"0b",	--1402
		x"12",	--1403
		x"0b",	--1404
		x"0a",	--1405
		x"7c",	--1406
		x"fb",	--1407
		x"81",	--1408
		x"02",	--1409
		x"81",	--1410
		x"04",	--1411
		x"1c",	--1412
		x"0d",	--1413
		x"79",	--1414
		x"1f",	--1415
		x"04",	--1416
		x"0c",	--1417
		x"0d",	--1418
		x"79",	--1419
		x"fc",	--1420
		x"3c",	--1421
		x"3d",	--1422
		x"0c",	--1423
		x"0d",	--1424
		x"1a",	--1425
		x"0b",	--1426
		x"0c",	--1427
		x"02",	--1428
		x"0d",	--1429
		x"e5",	--1430
		x"16",	--1431
		x"02",	--1432
		x"17",	--1433
		x"04",	--1434
		x"06",	--1435
		x"07",	--1436
		x"5f",	--1437
		x"01",	--1438
		x"5f",	--1439
		x"01",	--1440
		x"28",	--1441
		x"c8",	--1442
		x"01",	--1443
		x"a8",	--1444
		x"02",	--1445
		x"0e",	--1446
		x"0f",	--1447
		x"0e",	--1448
		x"0f",	--1449
		x"88",	--1450
		x"04",	--1451
		x"88",	--1452
		x"06",	--1453
		x"f8",	--1454
		x"03",	--1455
		x"00",	--1456
		x"0f",	--1457
		x"4d",	--1458
		x"0f",	--1459
		x"31",	--1460
		x"06",	--1461
		x"34",	--1462
		x"35",	--1463
		x"36",	--1464
		x"37",	--1465
		x"38",	--1466
		x"39",	--1467
		x"3a",	--1468
		x"3b",	--1469
		x"30",	--1470
		x"2b",	--1471
		x"67",	--1472
		x"81",	--1473
		x"00",	--1474
		x"04",	--1475
		x"05",	--1476
		x"5f",	--1477
		x"01",	--1478
		x"5f",	--1479
		x"01",	--1480
		x"d8",	--1481
		x"4f",	--1482
		x"68",	--1483
		x"0e",	--1484
		x"0f",	--1485
		x"0e",	--1486
		x"0f",	--1487
		x"0f",	--1488
		x"69",	--1489
		x"c8",	--1490
		x"01",	--1491
		x"a8",	--1492
		x"02",	--1493
		x"88",	--1494
		x"04",	--1495
		x"88",	--1496
		x"06",	--1497
		x"0c",	--1498
		x"0d",	--1499
		x"3c",	--1500
		x"3d",	--1501
		x"3d",	--1502
		x"ff",	--1503
		x"05",	--1504
		x"3d",	--1505
		x"00",	--1506
		x"17",	--1507
		x"3c",	--1508
		x"15",	--1509
		x"1b",	--1510
		x"02",	--1511
		x"3b",	--1512
		x"0e",	--1513
		x"0f",	--1514
		x"0a",	--1515
		x"3b",	--1516
		x"0c",	--1517
		x"0d",	--1518
		x"3c",	--1519
		x"3d",	--1520
		x"3d",	--1521
		x"ff",	--1522
		x"f5",	--1523
		x"3c",	--1524
		x"88",	--1525
		x"04",	--1526
		x"88",	--1527
		x"06",	--1528
		x"88",	--1529
		x"02",	--1530
		x"f8",	--1531
		x"03",	--1532
		x"00",	--1533
		x"0f",	--1534
		x"b3",	--1535
		x"0c",	--1536
		x"0d",	--1537
		x"1c",	--1538
		x"0d",	--1539
		x"12",	--1540
		x"0f",	--1541
		x"0e",	--1542
		x"0a",	--1543
		x"0b",	--1544
		x"0a",	--1545
		x"0b",	--1546
		x"88",	--1547
		x"04",	--1548
		x"88",	--1549
		x"06",	--1550
		x"98",	--1551
		x"02",	--1552
		x"0f",	--1553
		x"a1",	--1554
		x"6b",	--1555
		x"9f",	--1556
		x"ad",	--1557
		x"00",	--1558
		x"9d",	--1559
		x"02",	--1560
		x"02",	--1561
		x"9d",	--1562
		x"04",	--1563
		x"04",	--1564
		x"9d",	--1565
		x"06",	--1566
		x"06",	--1567
		x"5e",	--1568
		x"01",	--1569
		x"5e",	--1570
		x"01",	--1571
		x"cd",	--1572
		x"01",	--1573
		x"0f",	--1574
		x"8c",	--1575
		x"06",	--1576
		x"07",	--1577
		x"9a",	--1578
		x"39",	--1579
		x"19",	--1580
		x"39",	--1581
		x"20",	--1582
		x"8f",	--1583
		x"3e",	--1584
		x"3c",	--1585
		x"b6",	--1586
		x"c1",	--1587
		x"0e",	--1588
		x"0f",	--1589
		x"0e",	--1590
		x"0f",	--1591
		x"97",	--1592
		x"0f",	--1593
		x"79",	--1594
		x"d8",	--1595
		x"01",	--1596
		x"a8",	--1597
		x"02",	--1598
		x"3e",	--1599
		x"3f",	--1600
		x"1e",	--1601
		x"0f",	--1602
		x"88",	--1603
		x"04",	--1604
		x"88",	--1605
		x"06",	--1606
		x"92",	--1607
		x"0c",	--1608
		x"7b",	--1609
		x"81",	--1610
		x"00",	--1611
		x"81",	--1612
		x"02",	--1613
		x"81",	--1614
		x"04",	--1615
		x"4d",	--1616
		x"7d",	--1617
		x"1f",	--1618
		x"0c",	--1619
		x"4b",	--1620
		x"0c",	--1621
		x"0d",	--1622
		x"12",	--1623
		x"0d",	--1624
		x"0c",	--1625
		x"7b",	--1626
		x"fb",	--1627
		x"81",	--1628
		x"02",	--1629
		x"81",	--1630
		x"04",	--1631
		x"1c",	--1632
		x"0d",	--1633
		x"79",	--1634
		x"1f",	--1635
		x"04",	--1636
		x"0c",	--1637
		x"0d",	--1638
		x"79",	--1639
		x"fc",	--1640
		x"3c",	--1641
		x"3d",	--1642
		x"0c",	--1643
		x"0d",	--1644
		x"1a",	--1645
		x"0b",	--1646
		x"0c",	--1647
		x"04",	--1648
		x"0d",	--1649
		x"02",	--1650
		x"0a",	--1651
		x"0b",	--1652
		x"14",	--1653
		x"02",	--1654
		x"15",	--1655
		x"04",	--1656
		x"04",	--1657
		x"05",	--1658
		x"49",	--1659
		x"0a",	--1660
		x"0b",	--1661
		x"18",	--1662
		x"6c",	--1663
		x"33",	--1664
		x"df",	--1665
		x"01",	--1666
		x"01",	--1667
		x"2f",	--1668
		x"3f",	--1669
		x"0a",	--1670
		x"2c",	--1671
		x"31",	--1672
		x"e0",	--1673
		x"81",	--1674
		x"04",	--1675
		x"81",	--1676
		x"06",	--1677
		x"81",	--1678
		x"00",	--1679
		x"81",	--1680
		x"02",	--1681
		x"0e",	--1682
		x"3e",	--1683
		x"18",	--1684
		x"0f",	--1685
		x"2f",	--1686
		x"b0",	--1687
		x"32",	--1688
		x"0e",	--1689
		x"3e",	--1690
		x"10",	--1691
		x"0f",	--1692
		x"b0",	--1693
		x"32",	--1694
		x"0d",	--1695
		x"3d",	--1696
		x"0e",	--1697
		x"3e",	--1698
		x"10",	--1699
		x"0f",	--1700
		x"3f",	--1701
		x"18",	--1702
		x"b0",	--1703
		x"7e",	--1704
		x"b0",	--1705
		x"54",	--1706
		x"31",	--1707
		x"20",	--1708
		x"30",	--1709
		x"31",	--1710
		x"e0",	--1711
		x"81",	--1712
		x"04",	--1713
		x"81",	--1714
		x"06",	--1715
		x"81",	--1716
		x"00",	--1717
		x"81",	--1718
		x"02",	--1719
		x"0e",	--1720
		x"3e",	--1721
		x"18",	--1722
		x"0f",	--1723
		x"2f",	--1724
		x"b0",	--1725
		x"32",	--1726
		x"0e",	--1727
		x"3e",	--1728
		x"10",	--1729
		x"0f",	--1730
		x"b0",	--1731
		x"32",	--1732
		x"d1",	--1733
		x"11",	--1734
		x"0d",	--1735
		x"3d",	--1736
		x"0e",	--1737
		x"3e",	--1738
		x"10",	--1739
		x"0f",	--1740
		x"3f",	--1741
		x"18",	--1742
		x"b0",	--1743
		x"7e",	--1744
		x"b0",	--1745
		x"54",	--1746
		x"31",	--1747
		x"20",	--1748
		x"30",	--1749
		x"0b",	--1750
		x"0a",	--1751
		x"09",	--1752
		x"08",	--1753
		x"07",	--1754
		x"06",	--1755
		x"05",	--1756
		x"04",	--1757
		x"31",	--1758
		x"dc",	--1759
		x"81",	--1760
		x"04",	--1761
		x"81",	--1762
		x"06",	--1763
		x"81",	--1764
		x"00",	--1765
		x"81",	--1766
		x"02",	--1767
		x"0e",	--1768
		x"3e",	--1769
		x"18",	--1770
		x"0f",	--1771
		x"2f",	--1772
		x"b0",	--1773
		x"32",	--1774
		x"0e",	--1775
		x"3e",	--1776
		x"10",	--1777
		x"0f",	--1778
		x"b0",	--1779
		x"32",	--1780
		x"5f",	--1781
		x"18",	--1782
		x"6f",	--1783
		x"b6",	--1784
		x"5e",	--1785
		x"10",	--1786
		x"6e",	--1787
		x"d9",	--1788
		x"6f",	--1789
		x"ae",	--1790
		x"6e",	--1791
		x"e2",	--1792
		x"6f",	--1793
		x"ac",	--1794
		x"6e",	--1795
		x"d1",	--1796
		x"14",	--1797
		x"1c",	--1798
		x"15",	--1799
		x"1e",	--1800
		x"18",	--1801
		x"14",	--1802
		x"19",	--1803
		x"16",	--1804
		x"3c",	--1805
		x"20",	--1806
		x"0e",	--1807
		x"0f",	--1808
		x"06",	--1809
		x"07",	--1810
		x"81",	--1811
		x"20",	--1812
		x"81",	--1813
		x"22",	--1814
		x"0a",	--1815
		x"0b",	--1816
		x"81",	--1817
		x"20",	--1818
		x"08",	--1819
		x"08",	--1820
		x"09",	--1821
		x"12",	--1822
		x"05",	--1823
		x"04",	--1824
		x"b1",	--1825
		x"20",	--1826
		x"19",	--1827
		x"14",	--1828
		x"0d",	--1829
		x"0a",	--1830
		x"0b",	--1831
		x"0e",	--1832
		x"0f",	--1833
		x"1c",	--1834
		x"0d",	--1835
		x"0b",	--1836
		x"03",	--1837
		x"0b",	--1838
		x"0c",	--1839
		x"0d",	--1840
		x"0e",	--1841
		x"0f",	--1842
		x"06",	--1843
		x"07",	--1844
		x"09",	--1845
		x"e5",	--1846
		x"16",	--1847
		x"07",	--1848
		x"e2",	--1849
		x"0a",	--1850
		x"f5",	--1851
		x"f2",	--1852
		x"81",	--1853
		x"20",	--1854
		x"81",	--1855
		x"22",	--1856
		x"0c",	--1857
		x"1a",	--1858
		x"1a",	--1859
		x"1a",	--1860
		x"12",	--1861
		x"06",	--1862
		x"26",	--1863
		x"81",	--1864
		x"0a",	--1865
		x"5d",	--1866
		x"d1",	--1867
		x"11",	--1868
		x"19",	--1869
		x"83",	--1870
		x"c1",	--1871
		x"09",	--1872
		x"0c",	--1873
		x"3c",	--1874
		x"3f",	--1875
		x"00",	--1876
		x"18",	--1877
		x"1d",	--1878
		x"0a",	--1879
		x"3d",	--1880
		x"1a",	--1881
		x"20",	--1882
		x"1b",	--1883
		x"22",	--1884
		x"0c",	--1885
		x"0e",	--1886
		x"0f",	--1887
		x"0b",	--1888
		x"2a",	--1889
		x"0a",	--1890
		x"0b",	--1891
		x"3d",	--1892
		x"3f",	--1893
		x"00",	--1894
		x"f5",	--1895
		x"81",	--1896
		x"20",	--1897
		x"81",	--1898
		x"22",	--1899
		x"81",	--1900
		x"0a",	--1901
		x"0c",	--1902
		x"0d",	--1903
		x"3c",	--1904
		x"7f",	--1905
		x"0d",	--1906
		x"3c",	--1907
		x"40",	--1908
		x"44",	--1909
		x"81",	--1910
		x"0c",	--1911
		x"81",	--1912
		x"0e",	--1913
		x"f1",	--1914
		x"03",	--1915
		x"08",	--1916
		x"0f",	--1917
		x"3f",	--1918
		x"b0",	--1919
		x"54",	--1920
		x"31",	--1921
		x"24",	--1922
		x"34",	--1923
		x"35",	--1924
		x"36",	--1925
		x"37",	--1926
		x"38",	--1927
		x"39",	--1928
		x"3a",	--1929
		x"3b",	--1930
		x"30",	--1931
		x"1e",	--1932
		x"0f",	--1933
		x"d3",	--1934
		x"3a",	--1935
		x"03",	--1936
		x"08",	--1937
		x"1e",	--1938
		x"10",	--1939
		x"1c",	--1940
		x"20",	--1941
		x"1d",	--1942
		x"22",	--1943
		x"12",	--1944
		x"0d",	--1945
		x"0c",	--1946
		x"06",	--1947
		x"07",	--1948
		x"06",	--1949
		x"37",	--1950
		x"00",	--1951
		x"81",	--1952
		x"20",	--1953
		x"81",	--1954
		x"22",	--1955
		x"12",	--1956
		x"0f",	--1957
		x"0e",	--1958
		x"1a",	--1959
		x"0f",	--1960
		x"e7",	--1961
		x"81",	--1962
		x"0a",	--1963
		x"a6",	--1964
		x"6e",	--1965
		x"36",	--1966
		x"5f",	--1967
		x"d1",	--1968
		x"11",	--1969
		x"19",	--1970
		x"20",	--1971
		x"c1",	--1972
		x"19",	--1973
		x"0f",	--1974
		x"3f",	--1975
		x"18",	--1976
		x"c5",	--1977
		x"0d",	--1978
		x"ba",	--1979
		x"0c",	--1980
		x"0d",	--1981
		x"3c",	--1982
		x"80",	--1983
		x"0d",	--1984
		x"0c",	--1985
		x"b3",	--1986
		x"0d",	--1987
		x"b1",	--1988
		x"81",	--1989
		x"20",	--1990
		x"03",	--1991
		x"81",	--1992
		x"22",	--1993
		x"ab",	--1994
		x"3e",	--1995
		x"40",	--1996
		x"0f",	--1997
		x"3e",	--1998
		x"80",	--1999
		x"3f",	--2000
		x"a4",	--2001
		x"4d",	--2002
		x"7b",	--2003
		x"4f",	--2004
		x"de",	--2005
		x"5f",	--2006
		x"d1",	--2007
		x"11",	--2008
		x"19",	--2009
		x"06",	--2010
		x"c1",	--2011
		x"11",	--2012
		x"0f",	--2013
		x"3f",	--2014
		x"10",	--2015
		x"9e",	--2016
		x"4f",	--2017
		x"f8",	--2018
		x"6f",	--2019
		x"f1",	--2020
		x"3f",	--2021
		x"0a",	--2022
		x"97",	--2023
		x"0b",	--2024
		x"0a",	--2025
		x"09",	--2026
		x"08",	--2027
		x"07",	--2028
		x"31",	--2029
		x"e8",	--2030
		x"81",	--2031
		x"04",	--2032
		x"81",	--2033
		x"06",	--2034
		x"81",	--2035
		x"00",	--2036
		x"81",	--2037
		x"02",	--2038
		x"0e",	--2039
		x"3e",	--2040
		x"10",	--2041
		x"0f",	--2042
		x"2f",	--2043
		x"b0",	--2044
		x"32",	--2045
		x"0e",	--2046
		x"3e",	--2047
		x"0f",	--2048
		x"b0",	--2049
		x"32",	--2050
		x"5f",	--2051
		x"10",	--2052
		x"6f",	--2053
		x"5d",	--2054
		x"5e",	--2055
		x"08",	--2056
		x"6e",	--2057
		x"82",	--2058
		x"d1",	--2059
		x"09",	--2060
		x"11",	--2061
		x"6f",	--2062
		x"58",	--2063
		x"6f",	--2064
		x"56",	--2065
		x"6e",	--2066
		x"6f",	--2067
		x"6e",	--2068
		x"4c",	--2069
		x"1d",	--2070
		x"12",	--2071
		x"1d",	--2072
		x"0a",	--2073
		x"81",	--2074
		x"12",	--2075
		x"1e",	--2076
		x"14",	--2077
		x"1f",	--2078
		x"16",	--2079
		x"18",	--2080
		x"0c",	--2081
		x"19",	--2082
		x"0e",	--2083
		x"0f",	--2084
		x"1e",	--2085
		x"0e",	--2086
		x"0f",	--2087
		x"3d",	--2088
		x"81",	--2089
		x"12",	--2090
		x"37",	--2091
		x"1f",	--2092
		x"0c",	--2093
		x"3d",	--2094
		x"00",	--2095
		x"0a",	--2096
		x"0b",	--2097
		x"0b",	--2098
		x"0a",	--2099
		x"0b",	--2100
		x"0e",	--2101
		x"0f",	--2102
		x"12",	--2103
		x"0d",	--2104
		x"0c",	--2105
		x"0e",	--2106
		x"0f",	--2107
		x"37",	--2108
		x"0b",	--2109
		x"0f",	--2110
		x"f7",	--2111
		x"f2",	--2112
		x"0e",	--2113
		x"f4",	--2114
		x"ef",	--2115
		x"09",	--2116
		x"e5",	--2117
		x"0e",	--2118
		x"e3",	--2119
		x"dd",	--2120
		x"0c",	--2121
		x"0d",	--2122
		x"3c",	--2123
		x"7f",	--2124
		x"0d",	--2125
		x"3c",	--2126
		x"40",	--2127
		x"1c",	--2128
		x"81",	--2129
		x"14",	--2130
		x"81",	--2131
		x"16",	--2132
		x"0f",	--2133
		x"3f",	--2134
		x"10",	--2135
		x"b0",	--2136
		x"54",	--2137
		x"31",	--2138
		x"18",	--2139
		x"37",	--2140
		x"38",	--2141
		x"39",	--2142
		x"3a",	--2143
		x"3b",	--2144
		x"30",	--2145
		x"e1",	--2146
		x"10",	--2147
		x"0f",	--2148
		x"3f",	--2149
		x"10",	--2150
		x"f0",	--2151
		x"4f",	--2152
		x"fa",	--2153
		x"3f",	--2154
		x"0a",	--2155
		x"eb",	--2156
		x"0d",	--2157
		x"e2",	--2158
		x"0c",	--2159
		x"0d",	--2160
		x"3c",	--2161
		x"80",	--2162
		x"0d",	--2163
		x"0c",	--2164
		x"db",	--2165
		x"0d",	--2166
		x"d9",	--2167
		x"0e",	--2168
		x"02",	--2169
		x"0f",	--2170
		x"d5",	--2171
		x"3a",	--2172
		x"40",	--2173
		x"0b",	--2174
		x"3a",	--2175
		x"80",	--2176
		x"3b",	--2177
		x"ce",	--2178
		x"81",	--2179
		x"14",	--2180
		x"81",	--2181
		x"16",	--2182
		x"81",	--2183
		x"12",	--2184
		x"0f",	--2185
		x"3f",	--2186
		x"10",	--2187
		x"cb",	--2188
		x"0f",	--2189
		x"3f",	--2190
		x"c8",	--2191
		x"31",	--2192
		x"e8",	--2193
		x"81",	--2194
		x"04",	--2195
		x"81",	--2196
		x"06",	--2197
		x"81",	--2198
		x"00",	--2199
		x"81",	--2200
		x"02",	--2201
		x"0e",	--2202
		x"3e",	--2203
		x"10",	--2204
		x"0f",	--2205
		x"2f",	--2206
		x"b0",	--2207
		x"32",	--2208
		x"0e",	--2209
		x"3e",	--2210
		x"0f",	--2211
		x"b0",	--2212
		x"32",	--2213
		x"e1",	--2214
		x"10",	--2215
		x"0d",	--2216
		x"e1",	--2217
		x"08",	--2218
		x"0a",	--2219
		x"0e",	--2220
		x"3e",	--2221
		x"0f",	--2222
		x"3f",	--2223
		x"10",	--2224
		x"b0",	--2225
		x"56",	--2226
		x"31",	--2227
		x"18",	--2228
		x"30",	--2229
		x"3f",	--2230
		x"fb",	--2231
		x"31",	--2232
		x"f4",	--2233
		x"81",	--2234
		x"00",	--2235
		x"81",	--2236
		x"02",	--2237
		x"0e",	--2238
		x"2e",	--2239
		x"0f",	--2240
		x"b0",	--2241
		x"32",	--2242
		x"5f",	--2243
		x"04",	--2244
		x"6f",	--2245
		x"28",	--2246
		x"27",	--2247
		x"6f",	--2248
		x"07",	--2249
		x"1d",	--2250
		x"06",	--2251
		x"0d",	--2252
		x"21",	--2253
		x"3d",	--2254
		x"1f",	--2255
		x"09",	--2256
		x"c1",	--2257
		x"05",	--2258
		x"26",	--2259
		x"3e",	--2260
		x"3f",	--2261
		x"ff",	--2262
		x"31",	--2263
		x"0c",	--2264
		x"30",	--2265
		x"1e",	--2266
		x"08",	--2267
		x"1f",	--2268
		x"0a",	--2269
		x"3c",	--2270
		x"1e",	--2271
		x"4c",	--2272
		x"4d",	--2273
		x"7d",	--2274
		x"1f",	--2275
		x"0f",	--2276
		x"c1",	--2277
		x"05",	--2278
		x"ef",	--2279
		x"3e",	--2280
		x"3f",	--2281
		x"1e",	--2282
		x"0f",	--2283
		x"31",	--2284
		x"0c",	--2285
		x"30",	--2286
		x"0e",	--2287
		x"0f",	--2288
		x"31",	--2289
		x"0c",	--2290
		x"30",	--2291
		x"12",	--2292
		x"0f",	--2293
		x"0e",	--2294
		x"7d",	--2295
		x"fb",	--2296
		x"eb",	--2297
		x"0e",	--2298
		x"3f",	--2299
		x"00",	--2300
		x"31",	--2301
		x"0c",	--2302
		x"30",	--2303
		x"0b",	--2304
		x"0a",	--2305
		x"09",	--2306
		x"08",	--2307
		x"31",	--2308
		x"0a",	--2309
		x"0b",	--2310
		x"c1",	--2311
		x"01",	--2312
		x"0e",	--2313
		x"0d",	--2314
		x"0b",	--2315
		x"0b",	--2316
		x"e1",	--2317
		x"00",	--2318
		x"0f",	--2319
		x"b0",	--2320
		x"54",	--2321
		x"31",	--2322
		x"38",	--2323
		x"39",	--2324
		x"3a",	--2325
		x"3b",	--2326
		x"30",	--2327
		x"f1",	--2328
		x"03",	--2329
		x"00",	--2330
		x"b1",	--2331
		x"1e",	--2332
		x"02",	--2333
		x"81",	--2334
		x"04",	--2335
		x"81",	--2336
		x"06",	--2337
		x"0e",	--2338
		x"0f",	--2339
		x"b0",	--2340
		x"e2",	--2341
		x"3f",	--2342
		x"0f",	--2343
		x"18",	--2344
		x"e5",	--2345
		x"81",	--2346
		x"04",	--2347
		x"81",	--2348
		x"06",	--2349
		x"4e",	--2350
		x"7e",	--2351
		x"1f",	--2352
		x"06",	--2353
		x"3e",	--2354
		x"1e",	--2355
		x"0e",	--2356
		x"81",	--2357
		x"02",	--2358
		x"d7",	--2359
		x"91",	--2360
		x"04",	--2361
		x"04",	--2362
		x"91",	--2363
		x"06",	--2364
		x"06",	--2365
		x"7e",	--2366
		x"f8",	--2367
		x"f1",	--2368
		x"0e",	--2369
		x"3e",	--2370
		x"1e",	--2371
		x"1c",	--2372
		x"0d",	--2373
		x"48",	--2374
		x"78",	--2375
		x"1f",	--2376
		x"04",	--2377
		x"0c",	--2378
		x"0d",	--2379
		x"78",	--2380
		x"fc",	--2381
		x"3c",	--2382
		x"3d",	--2383
		x"0c",	--2384
		x"0d",	--2385
		x"18",	--2386
		x"09",	--2387
		x"0c",	--2388
		x"04",	--2389
		x"0d",	--2390
		x"02",	--2391
		x"08",	--2392
		x"09",	--2393
		x"7e",	--2394
		x"1f",	--2395
		x"0e",	--2396
		x"0d",	--2397
		x"0e",	--2398
		x"0d",	--2399
		x"0e",	--2400
		x"81",	--2401
		x"04",	--2402
		x"81",	--2403
		x"06",	--2404
		x"3e",	--2405
		x"1e",	--2406
		x"0e",	--2407
		x"81",	--2408
		x"02",	--2409
		x"a4",	--2410
		x"12",	--2411
		x"0b",	--2412
		x"0a",	--2413
		x"7e",	--2414
		x"fb",	--2415
		x"ec",	--2416
		x"0b",	--2417
		x"0a",	--2418
		x"09",	--2419
		x"1f",	--2420
		x"17",	--2421
		x"3e",	--2422
		x"00",	--2423
		x"2c",	--2424
		x"3a",	--2425
		x"18",	--2426
		x"0b",	--2427
		x"39",	--2428
		x"0c",	--2429
		x"0d",	--2430
		x"4f",	--2431
		x"4f",	--2432
		x"17",	--2433
		x"3c",	--2434
		x"12",	--2435
		x"6e",	--2436
		x"0f",	--2437
		x"0a",	--2438
		x"0b",	--2439
		x"0f",	--2440
		x"39",	--2441
		x"3a",	--2442
		x"3b",	--2443
		x"30",	--2444
		x"3f",	--2445
		x"00",	--2446
		x"0f",	--2447
		x"3a",	--2448
		x"0b",	--2449
		x"39",	--2450
		x"18",	--2451
		x"0c",	--2452
		x"0d",	--2453
		x"4f",	--2454
		x"4f",	--2455
		x"e9",	--2456
		x"12",	--2457
		x"0d",	--2458
		x"0c",	--2459
		x"7f",	--2460
		x"fb",	--2461
		x"e3",	--2462
		x"3a",	--2463
		x"10",	--2464
		x"0b",	--2465
		x"39",	--2466
		x"10",	--2467
		x"ef",	--2468
		x"3a",	--2469
		x"20",	--2470
		x"0b",	--2471
		x"09",	--2472
		x"ea",	--2473
		x"0b",	--2474
		x"0a",	--2475
		x"09",	--2476
		x"08",	--2477
		x"07",	--2478
		x"0d",	--2479
		x"1e",	--2480
		x"04",	--2481
		x"1f",	--2482
		x"06",	--2483
		x"5a",	--2484
		x"01",	--2485
		x"6c",	--2486
		x"6c",	--2487
		x"70",	--2488
		x"6c",	--2489
		x"6a",	--2490
		x"6c",	--2491
		x"36",	--2492
		x"0e",	--2493
		x"32",	--2494
		x"1b",	--2495
		x"02",	--2496
		x"3b",	--2497
		x"82",	--2498
		x"6d",	--2499
		x"3b",	--2500
		x"80",	--2501
		x"5e",	--2502
		x"0c",	--2503
		x"0d",	--2504
		x"3c",	--2505
		x"7f",	--2506
		x"0d",	--2507
		x"3c",	--2508
		x"40",	--2509
		x"40",	--2510
		x"3e",	--2511
		x"3f",	--2512
		x"0f",	--2513
		x"0f",	--2514
		x"4a",	--2515
		x"0d",	--2516
		x"3d",	--2517
		x"7f",	--2518
		x"12",	--2519
		x"0f",	--2520
		x"0e",	--2521
		x"12",	--2522
		x"0f",	--2523
		x"0e",	--2524
		x"12",	--2525
		x"0f",	--2526
		x"0e",	--2527
		x"12",	--2528
		x"0f",	--2529
		x"0e",	--2530
		x"12",	--2531
		x"0f",	--2532
		x"0e",	--2533
		x"12",	--2534
		x"0f",	--2535
		x"0e",	--2536
		x"12",	--2537
		x"0f",	--2538
		x"0e",	--2539
		x"3e",	--2540
		x"3f",	--2541
		x"7f",	--2542
		x"4d",	--2543
		x"05",	--2544
		x"0f",	--2545
		x"cc",	--2546
		x"4d",	--2547
		x"0e",	--2548
		x"0f",	--2549
		x"4d",	--2550
		x"0d",	--2551
		x"0d",	--2552
		x"0d",	--2553
		x"0d",	--2554
		x"0d",	--2555
		x"0d",	--2556
		x"0d",	--2557
		x"0c",	--2558
		x"3c",	--2559
		x"7f",	--2560
		x"0c",	--2561
		x"4f",	--2562
		x"0f",	--2563
		x"0f",	--2564
		x"0f",	--2565
		x"0d",	--2566
		x"0d",	--2567
		x"0f",	--2568
		x"37",	--2569
		x"38",	--2570
		x"39",	--2571
		x"3a",	--2572
		x"3b",	--2573
		x"30",	--2574
		x"0d",	--2575
		x"be",	--2576
		x"0c",	--2577
		x"0d",	--2578
		x"3c",	--2579
		x"80",	--2580
		x"0d",	--2581
		x"0c",	--2582
		x"02",	--2583
		x"0d",	--2584
		x"b8",	--2585
		x"3e",	--2586
		x"40",	--2587
		x"0f",	--2588
		x"b4",	--2589
		x"12",	--2590
		x"0f",	--2591
		x"0e",	--2592
		x"0d",	--2593
		x"3d",	--2594
		x"80",	--2595
		x"b2",	--2596
		x"7d",	--2597
		x"0e",	--2598
		x"0f",	--2599
		x"cd",	--2600
		x"0e",	--2601
		x"3f",	--2602
		x"10",	--2603
		x"3e",	--2604
		x"3f",	--2605
		x"7f",	--2606
		x"7d",	--2607
		x"c5",	--2608
		x"37",	--2609
		x"82",	--2610
		x"07",	--2611
		x"37",	--2612
		x"1a",	--2613
		x"4f",	--2614
		x"0c",	--2615
		x"0d",	--2616
		x"4b",	--2617
		x"7b",	--2618
		x"1f",	--2619
		x"05",	--2620
		x"12",	--2621
		x"0d",	--2622
		x"0c",	--2623
		x"7b",	--2624
		x"fb",	--2625
		x"18",	--2626
		x"09",	--2627
		x"77",	--2628
		x"1f",	--2629
		x"04",	--2630
		x"08",	--2631
		x"09",	--2632
		x"77",	--2633
		x"fc",	--2634
		x"38",	--2635
		x"39",	--2636
		x"08",	--2637
		x"09",	--2638
		x"1e",	--2639
		x"0f",	--2640
		x"08",	--2641
		x"04",	--2642
		x"09",	--2643
		x"02",	--2644
		x"0e",	--2645
		x"0f",	--2646
		x"08",	--2647
		x"09",	--2648
		x"08",	--2649
		x"09",	--2650
		x"0e",	--2651
		x"0f",	--2652
		x"3e",	--2653
		x"7f",	--2654
		x"0f",	--2655
		x"3e",	--2656
		x"40",	--2657
		x"26",	--2658
		x"38",	--2659
		x"3f",	--2660
		x"09",	--2661
		x"0e",	--2662
		x"0f",	--2663
		x"12",	--2664
		x"0f",	--2665
		x"0e",	--2666
		x"12",	--2667
		x"0f",	--2668
		x"0e",	--2669
		x"12",	--2670
		x"0f",	--2671
		x"0e",	--2672
		x"12",	--2673
		x"0f",	--2674
		x"0e",	--2675
		x"12",	--2676
		x"0f",	--2677
		x"0e",	--2678
		x"12",	--2679
		x"0f",	--2680
		x"0e",	--2681
		x"12",	--2682
		x"0f",	--2683
		x"0e",	--2684
		x"3e",	--2685
		x"3f",	--2686
		x"7f",	--2687
		x"5d",	--2688
		x"39",	--2689
		x"00",	--2690
		x"72",	--2691
		x"4d",	--2692
		x"70",	--2693
		x"08",	--2694
		x"09",	--2695
		x"da",	--2696
		x"0f",	--2697
		x"d8",	--2698
		x"0e",	--2699
		x"0f",	--2700
		x"3e",	--2701
		x"80",	--2702
		x"0f",	--2703
		x"0e",	--2704
		x"04",	--2705
		x"38",	--2706
		x"40",	--2707
		x"09",	--2708
		x"d0",	--2709
		x"0f",	--2710
		x"ce",	--2711
		x"f9",	--2712
		x"0b",	--2713
		x"0a",	--2714
		x"2a",	--2715
		x"5b",	--2716
		x"02",	--2717
		x"3b",	--2718
		x"7f",	--2719
		x"1d",	--2720
		x"02",	--2721
		x"12",	--2722
		x"0d",	--2723
		x"12",	--2724
		x"0d",	--2725
		x"12",	--2726
		x"0d",	--2727
		x"12",	--2728
		x"0d",	--2729
		x"12",	--2730
		x"0d",	--2731
		x"12",	--2732
		x"0d",	--2733
		x"12",	--2734
		x"0d",	--2735
		x"4d",	--2736
		x"5f",	--2737
		x"03",	--2738
		x"3f",	--2739
		x"80",	--2740
		x"0f",	--2741
		x"0f",	--2742
		x"ce",	--2743
		x"01",	--2744
		x"0d",	--2745
		x"2d",	--2746
		x"0a",	--2747
		x"51",	--2748
		x"be",	--2749
		x"82",	--2750
		x"02",	--2751
		x"0c",	--2752
		x"0d",	--2753
		x"0c",	--2754
		x"0d",	--2755
		x"0c",	--2756
		x"0d",	--2757
		x"0c",	--2758
		x"0d",	--2759
		x"0c",	--2760
		x"0d",	--2761
		x"0c",	--2762
		x"0d",	--2763
		x"0c",	--2764
		x"0d",	--2765
		x"0c",	--2766
		x"0d",	--2767
		x"fe",	--2768
		x"03",	--2769
		x"00",	--2770
		x"3d",	--2771
		x"00",	--2772
		x"0b",	--2773
		x"3f",	--2774
		x"81",	--2775
		x"0c",	--2776
		x"0d",	--2777
		x"0a",	--2778
		x"3f",	--2779
		x"3d",	--2780
		x"00",	--2781
		x"f9",	--2782
		x"8e",	--2783
		x"02",	--2784
		x"8e",	--2785
		x"04",	--2786
		x"8e",	--2787
		x"06",	--2788
		x"3a",	--2789
		x"3b",	--2790
		x"30",	--2791
		x"3d",	--2792
		x"ff",	--2793
		x"2a",	--2794
		x"3d",	--2795
		x"81",	--2796
		x"8e",	--2797
		x"02",	--2798
		x"fe",	--2799
		x"03",	--2800
		x"00",	--2801
		x"0c",	--2802
		x"0d",	--2803
		x"0c",	--2804
		x"0d",	--2805
		x"0c",	--2806
		x"0d",	--2807
		x"0c",	--2808
		x"0d",	--2809
		x"0c",	--2810
		x"0d",	--2811
		x"0c",	--2812
		x"0d",	--2813
		x"0c",	--2814
		x"0d",	--2815
		x"0c",	--2816
		x"0d",	--2817
		x"0a",	--2818
		x"0b",	--2819
		x"0a",	--2820
		x"3b",	--2821
		x"00",	--2822
		x"8e",	--2823
		x"04",	--2824
		x"8e",	--2825
		x"06",	--2826
		x"3a",	--2827
		x"3b",	--2828
		x"30",	--2829
		x"0b",	--2830
		x"ad",	--2831
		x"ee",	--2832
		x"00",	--2833
		x"3a",	--2834
		x"3b",	--2835
		x"30",	--2836
		x"0a",	--2837
		x"0c",	--2838
		x"0c",	--2839
		x"0d",	--2840
		x"0c",	--2841
		x"3d",	--2842
		x"10",	--2843
		x"0c",	--2844
		x"02",	--2845
		x"0d",	--2846
		x"08",	--2847
		x"de",	--2848
		x"00",	--2849
		x"e4",	--2850
		x"0b",	--2851
		x"f2",	--2852
		x"ee",	--2853
		x"00",	--2854
		x"e3",	--2855
		x"ce",	--2856
		x"00",	--2857
		x"dc",	--2858
		x"0b",	--2859
		x"6d",	--2860
		x"6d",	--2861
		x"12",	--2862
		x"6c",	--2863
		x"6c",	--2864
		x"0f",	--2865
		x"6d",	--2866
		x"41",	--2867
		x"6c",	--2868
		x"11",	--2869
		x"6d",	--2870
		x"0d",	--2871
		x"6c",	--2872
		x"14",	--2873
		x"5d",	--2874
		x"01",	--2875
		x"5d",	--2876
		x"01",	--2877
		x"14",	--2878
		x"4d",	--2879
		x"09",	--2880
		x"1e",	--2881
		x"0f",	--2882
		x"3b",	--2883
		x"30",	--2884
		x"6c",	--2885
		x"28",	--2886
		x"ce",	--2887
		x"01",	--2888
		x"f7",	--2889
		x"3e",	--2890
		x"0f",	--2891
		x"3b",	--2892
		x"30",	--2893
		x"cf",	--2894
		x"01",	--2895
		x"f0",	--2896
		x"3e",	--2897
		x"f8",	--2898
		x"1b",	--2899
		x"02",	--2900
		x"1c",	--2901
		x"02",	--2902
		x"0c",	--2903
		x"e6",	--2904
		x"0b",	--2905
		x"16",	--2906
		x"1b",	--2907
		x"04",	--2908
		x"1f",	--2909
		x"06",	--2910
		x"1c",	--2911
		x"04",	--2912
		x"1e",	--2913
		x"06",	--2914
		x"0e",	--2915
		x"da",	--2916
		x"0f",	--2917
		x"02",	--2918
		x"0c",	--2919
		x"d6",	--2920
		x"0f",	--2921
		x"06",	--2922
		x"0e",	--2923
		x"02",	--2924
		x"0b",	--2925
		x"02",	--2926
		x"0e",	--2927
		x"d1",	--2928
		x"4d",	--2929
		x"ce",	--2930
		x"3e",	--2931
		x"d6",	--2932
		x"6c",	--2933
		x"d7",	--2934
		x"5e",	--2935
		x"01",	--2936
		x"5f",	--2937
		x"01",	--2938
		x"0e",	--2939
		x"c5",	--2940
		x"0d",	--2941
		x"0f",	--2942
		x"04",	--2943
		x"3d",	--2944
		x"03",	--2945
		x"3f",	--2946
		x"1f",	--2947
		x"0e",	--2948
		x"03",	--2949
		x"5d",	--2950
		x"3e",	--2951
		x"1e",	--2952
		x"0d",	--2953
		x"b0",	--2954
		x"80",	--2955
		x"3d",	--2956
		x"6d",	--2957
		x"02",	--2958
		x"3e",	--2959
		x"1e",	--2960
		x"5d",	--2961
		x"02",	--2962
		x"3f",	--2963
		x"1f",	--2964
		x"30",	--2965
		x"b0",	--2966
		x"fa",	--2967
		x"0f",	--2968
		x"30",	--2969
		x"0b",	--2970
		x"0b",	--2971
		x"0f",	--2972
		x"06",	--2973
		x"3b",	--2974
		x"03",	--2975
		x"3e",	--2976
		x"3f",	--2977
		x"1e",	--2978
		x"0f",	--2979
		x"0d",	--2980
		x"05",	--2981
		x"5b",	--2982
		x"3c",	--2983
		x"3d",	--2984
		x"1c",	--2985
		x"0d",	--2986
		x"b0",	--2987
		x"a2",	--2988
		x"6b",	--2989
		x"04",	--2990
		x"3c",	--2991
		x"3d",	--2992
		x"1c",	--2993
		x"0d",	--2994
		x"5b",	--2995
		x"04",	--2996
		x"3e",	--2997
		x"3f",	--2998
		x"1e",	--2999
		x"0f",	--3000
		x"3b",	--3001
		x"30",	--3002
		x"b0",	--3003
		x"34",	--3004
		x"0e",	--3005
		x"0f",	--3006
		x"30",	--3007
		x"7c",	--3008
		x"10",	--3009
		x"0d",	--3010
		x"0e",	--3011
		x"0f",	--3012
		x"0e",	--3013
		x"0e",	--3014
		x"02",	--3015
		x"0e",	--3016
		x"1f",	--3017
		x"1c",	--3018
		x"f8",	--3019
		x"30",	--3020
		x"b0",	--3021
		x"80",	--3022
		x"0f",	--3023
		x"30",	--3024
		x"0b",	--3025
		x"0a",	--3026
		x"09",	--3027
		x"79",	--3028
		x"20",	--3029
		x"0a",	--3030
		x"0b",	--3031
		x"0c",	--3032
		x"0d",	--3033
		x"0e",	--3034
		x"0f",	--3035
		x"0c",	--3036
		x"0d",	--3037
		x"0d",	--3038
		x"06",	--3039
		x"02",	--3040
		x"0c",	--3041
		x"03",	--3042
		x"0c",	--3043
		x"0d",	--3044
		x"1e",	--3045
		x"19",	--3046
		x"f2",	--3047
		x"39",	--3048
		x"3a",	--3049
		x"3b",	--3050
		x"30",	--3051
		x"b0",	--3052
		x"a2",	--3053
		x"0e",	--3054
		x"0f",	--3055
		x"30",	--3056
		x"00",	--3057
		x"32",	--3058
		x"f0",	--3059
		x"fd",	--3060
		x"57",	--3061
		x"69",	--3062
		x"69",	--3063
		x"67",	--3064
		x"66",	--3065
		x"72",	--3066
		x"61",	--3067
		x"6e",	--3068
		x"77",	--3069
		x"2e",	--3070
		x"69",	--3071
		x"20",	--3072
		x"69",	--3073
		x"65",	--3074
		x"0a",	--3075
		x"57",	--3076
		x"20",	--3077
		x"68",	--3078
		x"75",	--3079
		x"64",	--3080
		x"6e",	--3081
		x"74",	--3082
		x"73",	--3083
		x"65",	--3084
		x"74",	--3085
		x"61",	--3086
		x"0d",	--3087
		x"00",	--3088
		x"6f",	--3089
		x"72",	--3090
		x"63",	--3091
		x"20",	--3092
		x"73",	--3093
		x"67",	--3094
		x"3a",	--3095
		x"0a",	--3096
		x"09",	--3097
		x"63",	--3098
		x"4c",	--3099
		x"46",	--3100
		x"20",	--3101
		x"49",	--3102
		x"48",	--3103
		x"0d",	--3104
		x"00",	--3105
		x"6f",	--3106
		x"65",	--3107
		x"68",	--3108
		x"6e",	--3109
		x"20",	--3110
		x"65",	--3111
		x"74",	--3112
		x"74",	--3113
		x"72",	--3114
		x"69",	--3115
		x"6c",	--3116
		x"20",	--3117
		x"72",	--3118
		x"6e",	--3119
		x"0d",	--3120
		x"00",	--3121
		x"0a",	--3122
		x"3d",	--3123
		x"3d",	--3124
		x"3d",	--3125
		x"4d",	--3126
		x"72",	--3127
		x"65",	--3128
		x"20",	--3129
		x"43",	--3130
		x"20",	--3131
		x"3d",	--3132
		x"3d",	--3133
		x"3d",	--3134
		x"0a",	--3135
		x"77",	--3136
		x"69",	--3137
		x"65",	--3138
		x"72",	--3139
		x"61",	--3140
		x"00",	--3141
		x"77",	--3142
		x"00",	--3143
		x"6f",	--3144
		x"74",	--3145
		x"6f",	--3146
		x"64",	--3147
		x"72",	--3148
		x"3e",	--3149
		x"00",	--3150
		x"0a",	--3151
		x"3a",	--3152
		x"73",	--3153
		x"0a",	--3154
		x"08",	--3155
		x"08",	--3156
		x"25",	--3157
		x"00",	--3158
		x"72",	--3159
		x"74",	--3160
		x"0a",	--3161
		x"00",	--3162
		x"6f",	--3163
		x"72",	--3164
		x"63",	--3165
		x"20",	--3166
		x"73",	--3167
		x"67",	--3168
		x"3a",	--3169
		x"0a",	--3170
		x"09",	--3171
		x"63",	--3172
		x"52",	--3173
		x"47",	--3174
		x"53",	--3175
		x"45",	--3176
		x"20",	--3177
		x"41",	--3178
		x"55",	--3179
		x"0d",	--3180
		x"00",	--3181
		x"6f",	--3182
		x"65",	--3183
		x"68",	--3184
		x"6e",	--3185
		x"20",	--3186
		x"65",	--3187
		x"74",	--3188
		x"74",	--3189
		x"72",	--3190
		x"69",	--3191
		x"6c",	--3192
		x"20",	--3193
		x"72",	--3194
		x"6e",	--3195
		x"0d",	--3196
		x"00",	--3197
		x"3d",	--3198
		x"64",	--3199
		x"76",	--3200
		x"25",	--3201
		x"0d",	--3202
		x"00",	--3203
		x"65",	--3204
		x"64",	--3205
		x"0d",	--3206
		x"09",	--3207
		x"63",	--3208
		x"52",	--3209
		x"47",	--3210
		x"53",	--3211
		x"45",	--3212
		x"0d",	--3213
		x"00",	--3214
		x"63",	--3215
		x"69",	--3216
		x"20",	--3217
		x"6f",	--3218
		x"20",	--3219
		x"20",	--3220
		x"75",	--3221
		x"62",	--3222
		x"72",	--3223
		x"0a",	--3224
		x"25",	--3225
		x"20",	--3226
		x"73",	--3227
		x"0a",	--3228
		x"25",	--3229
		x"3a",	--3230
		x"6e",	--3231
		x"20",	--3232
		x"75",	--3233
		x"68",	--3234
		x"63",	--3235
		x"6d",	--3236
		x"61",	--3237
		x"64",	--3238
		x"0a",	--3239
		x"84",	--3240
		x"b2",	--3241
		x"b2",	--3242
		x"b2",	--3243
		x"b2",	--3244
		x"b2",	--3245
		x"b2",	--3246
		x"b2",	--3247
		x"b2",	--3248
		x"b2",	--3249
		x"b2",	--3250
		x"b2",	--3251
		x"b2",	--3252
		x"b2",	--3253
		x"b2",	--3254
		x"b2",	--3255
		x"b2",	--3256
		x"b2",	--3257
		x"b2",	--3258
		x"b2",	--3259
		x"b2",	--3260
		x"b2",	--3261
		x"b2",	--3262
		x"b2",	--3263
		x"b2",	--3264
		x"b2",	--3265
		x"b2",	--3266
		x"b2",	--3267
		x"b2",	--3268
		x"76",	--3269
		x"b2",	--3270
		x"b2",	--3271
		x"b2",	--3272
		x"b2",	--3273
		x"b2",	--3274
		x"b2",	--3275
		x"b2",	--3276
		x"b2",	--3277
		x"b2",	--3278
		x"b2",	--3279
		x"b2",	--3280
		x"b2",	--3281
		x"b2",	--3282
		x"b2",	--3283
		x"b2",	--3284
		x"b2",	--3285
		x"b2",	--3286
		x"b2",	--3287
		x"b2",	--3288
		x"b2",	--3289
		x"b2",	--3290
		x"b2",	--3291
		x"b2",	--3292
		x"b2",	--3293
		x"b2",	--3294
		x"b2",	--3295
		x"b2",	--3296
		x"b2",	--3297
		x"b2",	--3298
		x"b2",	--3299
		x"b2",	--3300
		x"68",	--3301
		x"5a",	--3302
		x"4c",	--3303
		x"b2",	--3304
		x"b2",	--3305
		x"b2",	--3306
		x"b2",	--3307
		x"b2",	--3308
		x"b2",	--3309
		x"b2",	--3310
		x"34",	--3311
		x"b2",	--3312
		x"22",	--3313
		x"b2",	--3314
		x"b2",	--3315
		x"b2",	--3316
		x"b2",	--3317
		x"06",	--3318
		x"b2",	--3319
		x"b2",	--3320
		x"b2",	--3321
		x"f8",	--3322
		x"e6",	--3323
		x"30",	--3324
		x"32",	--3325
		x"34",	--3326
		x"36",	--3327
		x"38",	--3328
		x"61",	--3329
		x"63",	--3330
		x"65",	--3331
		x"00",	--3332
		x"00",	--3333
		x"00",	--3334
		x"00",	--3335
		x"00",	--3336
		x"00",	--3337
		x"02",	--3338
		x"03",	--3339
		x"03",	--3340
		x"04",	--3341
		x"04",	--3342
		x"04",	--3343
		x"04",	--3344
		x"05",	--3345
		x"05",	--3346
		x"05",	--3347
		x"05",	--3348
		x"05",	--3349
		x"05",	--3350
		x"05",	--3351
		x"05",	--3352
		x"06",	--3353
		x"06",	--3354
		x"06",	--3355
		x"06",	--3356
		x"06",	--3357
		x"06",	--3358
		x"06",	--3359
		x"06",	--3360
		x"06",	--3361
		x"06",	--3362
		x"06",	--3363
		x"06",	--3364
		x"06",	--3365
		x"06",	--3366
		x"06",	--3367
		x"06",	--3368
		x"07",	--3369
		x"07",	--3370
		x"07",	--3371
		x"07",	--3372
		x"07",	--3373
		x"07",	--3374
		x"07",	--3375
		x"07",	--3376
		x"07",	--3377
		x"07",	--3378
		x"07",	--3379
		x"07",	--3380
		x"07",	--3381
		x"07",	--3382
		x"07",	--3383
		x"07",	--3384
		x"07",	--3385
		x"07",	--3386
		x"07",	--3387
		x"07",	--3388
		x"07",	--3389
		x"07",	--3390
		x"07",	--3391
		x"07",	--3392
		x"07",	--3393
		x"07",	--3394
		x"07",	--3395
		x"07",	--3396
		x"07",	--3397
		x"07",	--3398
		x"07",	--3399
		x"07",	--3400
		x"08",	--3401
		x"08",	--3402
		x"08",	--3403
		x"08",	--3404
		x"08",	--3405
		x"08",	--3406
		x"08",	--3407
		x"08",	--3408
		x"08",	--3409
		x"08",	--3410
		x"08",	--3411
		x"08",	--3412
		x"08",	--3413
		x"08",	--3414
		x"08",	--3415
		x"08",	--3416
		x"08",	--3417
		x"08",	--3418
		x"08",	--3419
		x"08",	--3420
		x"08",	--3421
		x"08",	--3422
		x"08",	--3423
		x"08",	--3424
		x"08",	--3425
		x"08",	--3426
		x"08",	--3427
		x"08",	--3428
		x"08",	--3429
		x"08",	--3430
		x"08",	--3431
		x"08",	--3432
		x"08",	--3433
		x"08",	--3434
		x"08",	--3435
		x"08",	--3436
		x"08",	--3437
		x"08",	--3438
		x"08",	--3439
		x"08",	--3440
		x"08",	--3441
		x"08",	--3442
		x"08",	--3443
		x"08",	--3444
		x"08",	--3445
		x"08",	--3446
		x"08",	--3447
		x"08",	--3448
		x"08",	--3449
		x"08",	--3450
		x"08",	--3451
		x"08",	--3452
		x"08",	--3453
		x"08",	--3454
		x"08",	--3455
		x"08",	--3456
		x"08",	--3457
		x"08",	--3458
		x"08",	--3459
		x"08",	--3460
		x"08",	--3461
		x"08",	--3462
		x"08",	--3463
		x"08",	--3464
		x"68",	--3465
		x"6c",	--3466
		x"00",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"b8",	--4080
		x"b8",	--4081
		x"b8",	--4082
		x"b8",	--4083
		x"b8",	--4084
		x"b8",	--4085
		x"b8",	--4086
		x"8e",	--4087
		x"b8",	--4088
		x"b8",	--4089
		x"b8",	--4090
		x"b8",	--4091
		x"b8",	--4092
		x"b8",	--4093
		x"b8",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"03",	--5
		x"40",	--6
		x"06",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"03",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"fb",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"01",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"03",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"25",	--41
		x"43",	--42
		x"12",	--43
		x"e9",	--44
		x"12",	--45
		x"e6",	--46
		x"43",	--47
		x"00",	--48
		x"12",	--49
		x"f8",	--50
		x"12",	--51
		x"e8",	--52
		x"53",	--53
		x"40",	--54
		x"f8",	--55
		x"40",	--56
		x"e2",	--57
		x"40",	--58
		x"00",	--59
		x"12",	--60
		x"e6",	--61
		x"40",	--62
		x"f8",	--63
		x"40",	--64
		x"e3",	--65
		x"40",	--66
		x"00",	--67
		x"12",	--68
		x"e6",	--69
		x"40",	--70
		x"f8",	--71
		x"40",	--72
		x"e1",	--73
		x"40",	--74
		x"00",	--75
		x"12",	--76
		x"e6",	--77
		x"40",	--78
		x"f8",	--79
		x"40",	--80
		x"e1",	--81
		x"40",	--82
		x"00",	--83
		x"12",	--84
		x"e6",	--85
		x"43",	--86
		x"12",	--87
		x"e5",	--88
		x"43",	--89
		x"40",	--90
		x"4e",	--91
		x"40",	--92
		x"01",	--93
		x"41",	--94
		x"50",	--95
		x"00",	--96
		x"12",	--97
		x"e4",	--98
		x"41",	--99
		x"50",	--100
		x"00",	--101
		x"12",	--102
		x"e5",	--103
		x"43",	--104
		x"40",	--105
		x"4e",	--106
		x"40",	--107
		x"01",	--108
		x"41",	--109
		x"12",	--110
		x"e4",	--111
		x"41",	--112
		x"12",	--113
		x"e5",	--114
		x"41",	--115
		x"41",	--116
		x"50",	--117
		x"00",	--118
		x"12",	--119
		x"e1",	--120
		x"40",	--121
		x"ff",	--122
		x"00",	--123
		x"d2",	--124
		x"43",	--125
		x"12",	--126
		x"f8",	--127
		x"12",	--128
		x"e8",	--129
		x"53",	--130
		x"43",	--131
		x"d0",	--132
		x"00",	--133
		x"53",	--134
		x"90",	--135
		x"00",	--136
		x"24",	--137
		x"43",	--138
		x"4b",	--139
		x"f0",	--140
		x"00",	--141
		x"24",	--142
		x"5f",	--143
		x"53",	--144
		x"23",	--145
		x"4f",	--146
		x"3c",	--147
		x"43",	--148
		x"43",	--149
		x"4f",	--150
		x"00",	--151
		x"12",	--152
		x"e9",	--153
		x"93",	--154
		x"27",	--155
		x"12",	--156
		x"ea",	--157
		x"92",	--158
		x"24",	--159
		x"90",	--160
		x"00",	--161
		x"20",	--162
		x"12",	--163
		x"f8",	--164
		x"12",	--165
		x"e8",	--166
		x"53",	--167
		x"40",	--168
		x"00",	--169
		x"51",	--170
		x"5f",	--171
		x"43",	--172
		x"00",	--173
		x"12",	--174
		x"12",	--175
		x"f8",	--176
		x"12",	--177
		x"e8",	--178
		x"52",	--179
		x"41",	--180
		x"50",	--181
		x"00",	--182
		x"41",	--183
		x"00",	--184
		x"12",	--185
		x"e6",	--186
		x"3f",	--187
		x"93",	--188
		x"27",	--189
		x"53",	--190
		x"12",	--191
		x"f8",	--192
		x"12",	--193
		x"e8",	--194
		x"53",	--195
		x"3f",	--196
		x"90",	--197
		x"00",	--198
		x"2f",	--199
		x"4f",	--200
		x"11",	--201
		x"12",	--202
		x"12",	--203
		x"f8",	--204
		x"4f",	--205
		x"00",	--206
		x"12",	--207
		x"e8",	--208
		x"52",	--209
		x"40",	--210
		x"00",	--211
		x"51",	--212
		x"5a",	--213
		x"41",	--214
		x"00",	--215
		x"4f",	--216
		x"00",	--217
		x"53",	--218
		x"3f",	--219
		x"40",	--220
		x"f7",	--221
		x"40",	--222
		x"e0",	--223
		x"01",	--224
		x"42",	--225
		x"01",	--226
		x"40",	--227
		x"02",	--228
		x"01",	--229
		x"12",	--230
		x"f7",	--231
		x"12",	--232
		x"e8",	--233
		x"43",	--234
		x"01",	--235
		x"40",	--236
		x"f8",	--237
		x"00",	--238
		x"12",	--239
		x"e8",	--240
		x"53",	--241
		x"43",	--242
		x"41",	--243
		x"4f",	--244
		x"02",	--245
		x"4e",	--246
		x"02",	--247
		x"41",	--248
		x"82",	--249
		x"90",	--250
		x"00",	--251
		x"00",	--252
		x"20",	--253
		x"93",	--254
		x"00",	--255
		x"24",	--256
		x"41",	--257
		x"4f",	--258
		x"53",	--259
		x"41",	--260
		x"52",	--261
		x"12",	--262
		x"e3",	--263
		x"93",	--264
		x"00",	--265
		x"24",	--266
		x"41",	--267
		x"4f",	--268
		x"41",	--269
		x"53",	--270
		x"12",	--271
		x"e3",	--272
		x"93",	--273
		x"00",	--274
		x"24",	--275
		x"41",	--276
		x"00",	--277
		x"43",	--278
		x"12",	--279
		x"f2",	--280
		x"43",	--281
		x"40",	--282
		x"42",	--283
		x"12",	--284
		x"ef",	--285
		x"4e",	--286
		x"4f",	--287
		x"42",	--288
		x"02",	--289
		x"12",	--290
		x"e5",	--291
		x"41",	--292
		x"00",	--293
		x"43",	--294
		x"12",	--295
		x"f2",	--296
		x"43",	--297
		x"40",	--298
		x"42",	--299
		x"12",	--300
		x"ef",	--301
		x"4e",	--302
		x"4f",	--303
		x"42",	--304
		x"02",	--305
		x"12",	--306
		x"e5",	--307
		x"43",	--308
		x"52",	--309
		x"41",	--310
		x"12",	--311
		x"f8",	--312
		x"4f",	--313
		x"00",	--314
		x"12",	--315
		x"e8",	--316
		x"41",	--317
		x"00",	--318
		x"4f",	--319
		x"11",	--320
		x"4f",	--321
		x"00",	--322
		x"12",	--323
		x"f8",	--324
		x"12",	--325
		x"e8",	--326
		x"52",	--327
		x"43",	--328
		x"52",	--329
		x"41",	--330
		x"12",	--331
		x"f8",	--332
		x"12",	--333
		x"e8",	--334
		x"53",	--335
		x"43",	--336
		x"3f",	--337
		x"12",	--338
		x"50",	--339
		x"ff",	--340
		x"4f",	--341
		x"12",	--342
		x"f8",	--343
		x"12",	--344
		x"e8",	--345
		x"53",	--346
		x"90",	--347
		x"00",	--348
		x"00",	--349
		x"20",	--350
		x"93",	--351
		x"00",	--352
		x"24",	--353
		x"41",	--354
		x"4b",	--355
		x"53",	--356
		x"41",	--357
		x"52",	--358
		x"12",	--359
		x"e3",	--360
		x"93",	--361
		x"00",	--362
		x"24",	--363
		x"41",	--364
		x"4f",	--365
		x"41",	--366
		x"53",	--367
		x"12",	--368
		x"e3",	--369
		x"93",	--370
		x"00",	--371
		x"24",	--372
		x"12",	--373
		x"00",	--374
		x"12",	--375
		x"00",	--376
		x"12",	--377
		x"f8",	--378
		x"12",	--379
		x"e8",	--380
		x"50",	--381
		x"00",	--382
		x"41",	--383
		x"00",	--384
		x"41",	--385
		x"00",	--386
		x"00",	--387
		x"43",	--388
		x"50",	--389
		x"00",	--390
		x"41",	--391
		x"41",	--392
		x"12",	--393
		x"f8",	--394
		x"12",	--395
		x"e8",	--396
		x"4b",	--397
		x"11",	--398
		x"4f",	--399
		x"00",	--400
		x"12",	--401
		x"f8",	--402
		x"12",	--403
		x"e8",	--404
		x"52",	--405
		x"43",	--406
		x"50",	--407
		x"00",	--408
		x"41",	--409
		x"41",	--410
		x"12",	--411
		x"f8",	--412
		x"12",	--413
		x"e8",	--414
		x"53",	--415
		x"43",	--416
		x"3f",	--417
		x"12",	--418
		x"82",	--419
		x"4f",	--420
		x"12",	--421
		x"f9",	--422
		x"12",	--423
		x"e8",	--424
		x"53",	--425
		x"90",	--426
		x"00",	--427
		x"00",	--428
		x"20",	--429
		x"93",	--430
		x"00",	--431
		x"24",	--432
		x"41",	--433
		x"4b",	--434
		x"53",	--435
		x"41",	--436
		x"53",	--437
		x"12",	--438
		x"e3",	--439
		x"93",	--440
		x"00",	--441
		x"24",	--442
		x"41",	--443
		x"00",	--444
		x"12",	--445
		x"12",	--446
		x"12",	--447
		x"f8",	--448
		x"12",	--449
		x"e8",	--450
		x"50",	--451
		x"00",	--452
		x"43",	--453
		x"52",	--454
		x"41",	--455
		x"41",	--456
		x"12",	--457
		x"f8",	--458
		x"12",	--459
		x"e8",	--460
		x"4b",	--461
		x"11",	--462
		x"4f",	--463
		x"00",	--464
		x"12",	--465
		x"f9",	--466
		x"12",	--467
		x"e8",	--468
		x"52",	--469
		x"43",	--470
		x"52",	--471
		x"41",	--472
		x"41",	--473
		x"12",	--474
		x"f8",	--475
		x"12",	--476
		x"e8",	--477
		x"53",	--478
		x"43",	--479
		x"3f",	--480
		x"12",	--481
		x"12",	--482
		x"12",	--483
		x"12",	--484
		x"12",	--485
		x"43",	--486
		x"00",	--487
		x"43",	--488
		x"00",	--489
		x"4e",	--490
		x"93",	--491
		x"24",	--492
		x"4e",	--493
		x"53",	--494
		x"4e",	--495
		x"43",	--496
		x"43",	--497
		x"43",	--498
		x"3c",	--499
		x"90",	--500
		x"00",	--501
		x"2c",	--502
		x"4f",	--503
		x"5c",	--504
		x"5c",	--505
		x"5c",	--506
		x"5c",	--507
		x"4c",	--508
		x"00",	--509
		x"50",	--510
		x"ff",	--511
		x"48",	--512
		x"11",	--513
		x"5a",	--514
		x"4c",	--515
		x"00",	--516
		x"43",	--517
		x"53",	--518
		x"49",	--519
		x"4b",	--520
		x"4b",	--521
		x"93",	--522
		x"24",	--523
		x"90",	--524
		x"00",	--525
		x"24",	--526
		x"90",	--527
		x"00",	--528
		x"24",	--529
		x"4c",	--530
		x"50",	--531
		x"ff",	--532
		x"93",	--533
		x"23",	--534
		x"90",	--535
		x"00",	--536
		x"2c",	--537
		x"4f",	--538
		x"5a",	--539
		x"4a",	--540
		x"5c",	--541
		x"5c",	--542
		x"5a",	--543
		x"4c",	--544
		x"00",	--545
		x"50",	--546
		x"ff",	--547
		x"48",	--548
		x"11",	--549
		x"58",	--550
		x"4c",	--551
		x"00",	--552
		x"3f",	--553
		x"43",	--554
		x"3f",	--555
		x"4c",	--556
		x"50",	--557
		x"ff",	--558
		x"90",	--559
		x"00",	--560
		x"2c",	--561
		x"4f",	--562
		x"5c",	--563
		x"5c",	--564
		x"5c",	--565
		x"5c",	--566
		x"4c",	--567
		x"00",	--568
		x"50",	--569
		x"ff",	--570
		x"3f",	--571
		x"4c",	--572
		x"50",	--573
		x"ff",	--574
		x"90",	--575
		x"00",	--576
		x"2c",	--577
		x"4f",	--578
		x"5c",	--579
		x"5c",	--580
		x"5c",	--581
		x"5c",	--582
		x"4c",	--583
		x"00",	--584
		x"50",	--585
		x"ff",	--586
		x"3f",	--587
		x"43",	--588
		x"00",	--589
		x"43",	--590
		x"41",	--591
		x"41",	--592
		x"41",	--593
		x"41",	--594
		x"41",	--595
		x"41",	--596
		x"43",	--597
		x"00",	--598
		x"4a",	--599
		x"53",	--600
		x"5e",	--601
		x"41",	--602
		x"41",	--603
		x"41",	--604
		x"41",	--605
		x"41",	--606
		x"41",	--607
		x"11",	--608
		x"12",	--609
		x"12",	--610
		x"f9",	--611
		x"12",	--612
		x"e8",	--613
		x"52",	--614
		x"43",	--615
		x"41",	--616
		x"41",	--617
		x"41",	--618
		x"41",	--619
		x"41",	--620
		x"41",	--621
		x"12",	--622
		x"12",	--623
		x"4e",	--624
		x"4c",	--625
		x"4e",	--626
		x"00",	--627
		x"4d",	--628
		x"00",	--629
		x"4c",	--630
		x"00",	--631
		x"4d",	--632
		x"43",	--633
		x"40",	--634
		x"36",	--635
		x"40",	--636
		x"01",	--637
		x"12",	--638
		x"f7",	--639
		x"4e",	--640
		x"00",	--641
		x"12",	--642
		x"c2",	--643
		x"43",	--644
		x"4a",	--645
		x"01",	--646
		x"40",	--647
		x"00",	--648
		x"01",	--649
		x"42",	--650
		x"01",	--651
		x"00",	--652
		x"41",	--653
		x"43",	--654
		x"41",	--655
		x"41",	--656
		x"41",	--657
		x"12",	--658
		x"12",	--659
		x"12",	--660
		x"43",	--661
		x"00",	--662
		x"40",	--663
		x"3f",	--664
		x"00",	--665
		x"4f",	--666
		x"4b",	--667
		x"00",	--668
		x"43",	--669
		x"12",	--670
		x"f2",	--671
		x"43",	--672
		x"40",	--673
		x"3f",	--674
		x"12",	--675
		x"ed",	--676
		x"4e",	--677
		x"4f",	--678
		x"4b",	--679
		x"00",	--680
		x"43",	--681
		x"12",	--682
		x"f2",	--683
		x"4e",	--684
		x"4f",	--685
		x"48",	--686
		x"49",	--687
		x"12",	--688
		x"ed",	--689
		x"12",	--690
		x"ea",	--691
		x"4e",	--692
		x"00",	--693
		x"43",	--694
		x"00",	--695
		x"41",	--696
		x"41",	--697
		x"41",	--698
		x"41",	--699
		x"12",	--700
		x"12",	--701
		x"12",	--702
		x"4d",	--703
		x"4e",	--704
		x"4d",	--705
		x"00",	--706
		x"4e",	--707
		x"00",	--708
		x"4f",	--709
		x"49",	--710
		x"00",	--711
		x"43",	--712
		x"12",	--713
		x"f2",	--714
		x"4e",	--715
		x"4f",	--716
		x"4a",	--717
		x"4b",	--718
		x"12",	--719
		x"ed",	--720
		x"4e",	--721
		x"4f",	--722
		x"49",	--723
		x"00",	--724
		x"43",	--725
		x"12",	--726
		x"f2",	--727
		x"4e",	--728
		x"4f",	--729
		x"4a",	--730
		x"4b",	--731
		x"12",	--732
		x"ed",	--733
		x"12",	--734
		x"ea",	--735
		x"4e",	--736
		x"00",	--737
		x"41",	--738
		x"41",	--739
		x"41",	--740
		x"41",	--741
		x"12",	--742
		x"12",	--743
		x"93",	--744
		x"02",	--745
		x"38",	--746
		x"40",	--747
		x"02",	--748
		x"43",	--749
		x"12",	--750
		x"4b",	--751
		x"ff",	--752
		x"11",	--753
		x"12",	--754
		x"12",	--755
		x"f9",	--756
		x"12",	--757
		x"e8",	--758
		x"50",	--759
		x"00",	--760
		x"53",	--761
		x"50",	--762
		x"00",	--763
		x"92",	--764
		x"02",	--765
		x"3b",	--766
		x"43",	--767
		x"41",	--768
		x"41",	--769
		x"41",	--770
		x"42",	--771
		x"02",	--772
		x"90",	--773
		x"00",	--774
		x"34",	--775
		x"4e",	--776
		x"5f",	--777
		x"5e",	--778
		x"5f",	--779
		x"50",	--780
		x"02",	--781
		x"40",	--782
		x"00",	--783
		x"00",	--784
		x"40",	--785
		x"e5",	--786
		x"00",	--787
		x"40",	--788
		x"02",	--789
		x"00",	--790
		x"53",	--791
		x"4e",	--792
		x"02",	--793
		x"41",	--794
		x"12",	--795
		x"42",	--796
		x"02",	--797
		x"90",	--798
		x"00",	--799
		x"34",	--800
		x"4b",	--801
		x"5c",	--802
		x"5b",	--803
		x"5c",	--804
		x"50",	--805
		x"02",	--806
		x"4f",	--807
		x"00",	--808
		x"4e",	--809
		x"00",	--810
		x"4d",	--811
		x"00",	--812
		x"53",	--813
		x"4b",	--814
		x"02",	--815
		x"43",	--816
		x"41",	--817
		x"41",	--818
		x"43",	--819
		x"3f",	--820
		x"12",	--821
		x"42",	--822
		x"02",	--823
		x"93",	--824
		x"38",	--825
		x"92",	--826
		x"02",	--827
		x"24",	--828
		x"40",	--829
		x"02",	--830
		x"43",	--831
		x"3c",	--832
		x"50",	--833
		x"00",	--834
		x"9f",	--835
		x"ff",	--836
		x"24",	--837
		x"53",	--838
		x"9b",	--839
		x"23",	--840
		x"12",	--841
		x"f9",	--842
		x"12",	--843
		x"e8",	--844
		x"53",	--845
		x"43",	--846
		x"41",	--847
		x"41",	--848
		x"43",	--849
		x"4c",	--850
		x"5d",	--851
		x"5d",	--852
		x"5c",	--853
		x"50",	--854
		x"02",	--855
		x"4e",	--856
		x"12",	--857
		x"00",	--858
		x"41",	--859
		x"41",	--860
		x"42",	--861
		x"00",	--862
		x"f2",	--863
		x"23",	--864
		x"4f",	--865
		x"00",	--866
		x"43",	--867
		x"41",	--868
		x"f0",	--869
		x"00",	--870
		x"4f",	--871
		x"f9",	--872
		x"11",	--873
		x"12",	--874
		x"e6",	--875
		x"41",	--876
		x"12",	--877
		x"4f",	--878
		x"4f",	--879
		x"11",	--880
		x"11",	--881
		x"11",	--882
		x"11",	--883
		x"4e",	--884
		x"12",	--885
		x"e6",	--886
		x"4b",	--887
		x"12",	--888
		x"e6",	--889
		x"41",	--890
		x"41",	--891
		x"12",	--892
		x"12",	--893
		x"4f",	--894
		x"40",	--895
		x"00",	--896
		x"4a",	--897
		x"4b",	--898
		x"f0",	--899
		x"00",	--900
		x"24",	--901
		x"11",	--902
		x"53",	--903
		x"23",	--904
		x"f3",	--905
		x"24",	--906
		x"40",	--907
		x"00",	--908
		x"12",	--909
		x"e6",	--910
		x"53",	--911
		x"93",	--912
		x"23",	--913
		x"41",	--914
		x"41",	--915
		x"41",	--916
		x"40",	--917
		x"00",	--918
		x"3f",	--919
		x"12",	--920
		x"4f",	--921
		x"4f",	--922
		x"10",	--923
		x"11",	--924
		x"4e",	--925
		x"12",	--926
		x"e6",	--927
		x"4b",	--928
		x"12",	--929
		x"e6",	--930
		x"41",	--931
		x"41",	--932
		x"12",	--933
		x"12",	--934
		x"4e",	--935
		x"4f",	--936
		x"4f",	--937
		x"10",	--938
		x"11",	--939
		x"4d",	--940
		x"12",	--941
		x"e6",	--942
		x"4b",	--943
		x"12",	--944
		x"e6",	--945
		x"4b",	--946
		x"4a",	--947
		x"10",	--948
		x"10",	--949
		x"ec",	--950
		x"ec",	--951
		x"4d",	--952
		x"12",	--953
		x"e6",	--954
		x"4a",	--955
		x"12",	--956
		x"e6",	--957
		x"41",	--958
		x"41",	--959
		x"41",	--960
		x"12",	--961
		x"12",	--962
		x"12",	--963
		x"4f",	--964
		x"93",	--965
		x"24",	--966
		x"4e",	--967
		x"53",	--968
		x"43",	--969
		x"4a",	--970
		x"5b",	--971
		x"4d",	--972
		x"11",	--973
		x"12",	--974
		x"e6",	--975
		x"99",	--976
		x"24",	--977
		x"53",	--978
		x"b0",	--979
		x"00",	--980
		x"20",	--981
		x"40",	--982
		x"00",	--983
		x"12",	--984
		x"e6",	--985
		x"3f",	--986
		x"40",	--987
		x"00",	--988
		x"12",	--989
		x"e6",	--990
		x"3f",	--991
		x"41",	--992
		x"41",	--993
		x"41",	--994
		x"41",	--995
		x"12",	--996
		x"12",	--997
		x"12",	--998
		x"4f",	--999
		x"93",	--1000
		x"24",	--1001
		x"4e",	--1002
		x"53",	--1003
		x"43",	--1004
		x"4a",	--1005
		x"11",	--1006
		x"12",	--1007
		x"e6",	--1008
		x"99",	--1009
		x"24",	--1010
		x"53",	--1011
		x"b0",	--1012
		x"00",	--1013
		x"23",	--1014
		x"40",	--1015
		x"00",	--1016
		x"12",	--1017
		x"e6",	--1018
		x"4a",	--1019
		x"11",	--1020
		x"12",	--1021
		x"e6",	--1022
		x"99",	--1023
		x"23",	--1024
		x"41",	--1025
		x"41",	--1026
		x"41",	--1027
		x"41",	--1028
		x"12",	--1029
		x"12",	--1030
		x"12",	--1031
		x"50",	--1032
		x"ff",	--1033
		x"4f",	--1034
		x"93",	--1035
		x"38",	--1036
		x"90",	--1037
		x"00",	--1038
		x"38",	--1039
		x"43",	--1040
		x"41",	--1041
		x"59",	--1042
		x"40",	--1043
		x"00",	--1044
		x"4b",	--1045
		x"12",	--1046
		x"f7",	--1047
		x"50",	--1048
		x"00",	--1049
		x"4f",	--1050
		x"00",	--1051
		x"53",	--1052
		x"40",	--1053
		x"00",	--1054
		x"4b",	--1055
		x"12",	--1056
		x"f6",	--1057
		x"4f",	--1058
		x"90",	--1059
		x"00",	--1060
		x"37",	--1061
		x"49",	--1062
		x"53",	--1063
		x"51",	--1064
		x"40",	--1065
		x"00",	--1066
		x"4b",	--1067
		x"12",	--1068
		x"f7",	--1069
		x"50",	--1070
		x"00",	--1071
		x"4f",	--1072
		x"00",	--1073
		x"53",	--1074
		x"41",	--1075
		x"5a",	--1076
		x"4f",	--1077
		x"11",	--1078
		x"12",	--1079
		x"e6",	--1080
		x"93",	--1081
		x"23",	--1082
		x"50",	--1083
		x"00",	--1084
		x"41",	--1085
		x"41",	--1086
		x"41",	--1087
		x"41",	--1088
		x"40",	--1089
		x"00",	--1090
		x"12",	--1091
		x"e6",	--1092
		x"e3",	--1093
		x"53",	--1094
		x"3f",	--1095
		x"43",	--1096
		x"43",	--1097
		x"3f",	--1098
		x"12",	--1099
		x"12",	--1100
		x"12",	--1101
		x"41",	--1102
		x"52",	--1103
		x"4b",	--1104
		x"49",	--1105
		x"93",	--1106
		x"20",	--1107
		x"3c",	--1108
		x"11",	--1109
		x"12",	--1110
		x"e6",	--1111
		x"49",	--1112
		x"4a",	--1113
		x"53",	--1114
		x"4a",	--1115
		x"00",	--1116
		x"93",	--1117
		x"24",	--1118
		x"90",	--1119
		x"00",	--1120
		x"23",	--1121
		x"49",	--1122
		x"53",	--1123
		x"49",	--1124
		x"00",	--1125
		x"50",	--1126
		x"ff",	--1127
		x"90",	--1128
		x"00",	--1129
		x"2f",	--1130
		x"4f",	--1131
		x"5f",	--1132
		x"4f",	--1133
		x"f9",	--1134
		x"41",	--1135
		x"41",	--1136
		x"41",	--1137
		x"41",	--1138
		x"4b",	--1139
		x"52",	--1140
		x"4b",	--1141
		x"00",	--1142
		x"4b",	--1143
		x"12",	--1144
		x"e7",	--1145
		x"49",	--1146
		x"3f",	--1147
		x"4b",	--1148
		x"53",	--1149
		x"4b",	--1150
		x"12",	--1151
		x"e7",	--1152
		x"49",	--1153
		x"3f",	--1154
		x"4b",	--1155
		x"53",	--1156
		x"4f",	--1157
		x"49",	--1158
		x"93",	--1159
		x"27",	--1160
		x"53",	--1161
		x"11",	--1162
		x"12",	--1163
		x"e6",	--1164
		x"49",	--1165
		x"93",	--1166
		x"23",	--1167
		x"3f",	--1168
		x"4b",	--1169
		x"52",	--1170
		x"4b",	--1171
		x"00",	--1172
		x"4b",	--1173
		x"12",	--1174
		x"e7",	--1175
		x"49",	--1176
		x"3f",	--1177
		x"4b",	--1178
		x"53",	--1179
		x"4b",	--1180
		x"4e",	--1181
		x"10",	--1182
		x"11",	--1183
		x"10",	--1184
		x"11",	--1185
		x"12",	--1186
		x"e7",	--1187
		x"49",	--1188
		x"3f",	--1189
		x"4b",	--1190
		x"53",	--1191
		x"4b",	--1192
		x"12",	--1193
		x"e8",	--1194
		x"49",	--1195
		x"3f",	--1196
		x"4b",	--1197
		x"53",	--1198
		x"4b",	--1199
		x"12",	--1200
		x"e6",	--1201
		x"49",	--1202
		x"3f",	--1203
		x"4b",	--1204
		x"53",	--1205
		x"4b",	--1206
		x"12",	--1207
		x"e6",	--1208
		x"49",	--1209
		x"3f",	--1210
		x"4b",	--1211
		x"53",	--1212
		x"4b",	--1213
		x"12",	--1214
		x"e6",	--1215
		x"49",	--1216
		x"3f",	--1217
		x"40",	--1218
		x"00",	--1219
		x"12",	--1220
		x"e6",	--1221
		x"3f",	--1222
		x"12",	--1223
		x"12",	--1224
		x"42",	--1225
		x"02",	--1226
		x"42",	--1227
		x"00",	--1228
		x"03",	--1229
		x"42",	--1230
		x"02",	--1231
		x"90",	--1232
		x"00",	--1233
		x"34",	--1234
		x"53",	--1235
		x"02",	--1236
		x"42",	--1237
		x"02",	--1238
		x"42",	--1239
		x"02",	--1240
		x"9f",	--1241
		x"20",	--1242
		x"53",	--1243
		x"02",	--1244
		x"40",	--1245
		x"00",	--1246
		x"00",	--1247
		x"c0",	--1248
		x"00",	--1249
		x"00",	--1250
		x"41",	--1251
		x"41",	--1252
		x"c0",	--1253
		x"00",	--1254
		x"00",	--1255
		x"13",	--1256
		x"43",	--1257
		x"02",	--1258
		x"3f",	--1259
		x"40",	--1260
		x"09",	--1261
		x"00",	--1262
		x"40",	--1263
		x"00",	--1264
		x"00",	--1265
		x"41",	--1266
		x"42",	--1267
		x"02",	--1268
		x"42",	--1269
		x"02",	--1270
		x"9f",	--1271
		x"38",	--1272
		x"42",	--1273
		x"02",	--1274
		x"82",	--1275
		x"02",	--1276
		x"41",	--1277
		x"42",	--1278
		x"02",	--1279
		x"42",	--1280
		x"02",	--1281
		x"40",	--1282
		x"00",	--1283
		x"8d",	--1284
		x"8e",	--1285
		x"41",	--1286
		x"42",	--1287
		x"02",	--1288
		x"4f",	--1289
		x"03",	--1290
		x"42",	--1291
		x"02",	--1292
		x"42",	--1293
		x"02",	--1294
		x"9e",	--1295
		x"24",	--1296
		x"42",	--1297
		x"02",	--1298
		x"90",	--1299
		x"00",	--1300
		x"38",	--1301
		x"43",	--1302
		x"02",	--1303
		x"41",	--1304
		x"53",	--1305
		x"02",	--1306
		x"41",	--1307
		x"43",	--1308
		x"41",	--1309
		x"12",	--1310
		x"12",	--1311
		x"4e",	--1312
		x"4f",	--1313
		x"43",	--1314
		x"40",	--1315
		x"4f",	--1316
		x"12",	--1317
		x"f1",	--1318
		x"93",	--1319
		x"34",	--1320
		x"4a",	--1321
		x"4b",	--1322
		x"12",	--1323
		x"f1",	--1324
		x"41",	--1325
		x"41",	--1326
		x"41",	--1327
		x"43",	--1328
		x"40",	--1329
		x"4f",	--1330
		x"4a",	--1331
		x"4b",	--1332
		x"12",	--1333
		x"ed",	--1334
		x"12",	--1335
		x"f1",	--1336
		x"53",	--1337
		x"60",	--1338
		x"80",	--1339
		x"41",	--1340
		x"41",	--1341
		x"41",	--1342
		x"12",	--1343
		x"12",	--1344
		x"12",	--1345
		x"12",	--1346
		x"12",	--1347
		x"12",	--1348
		x"12",	--1349
		x"12",	--1350
		x"50",	--1351
		x"ff",	--1352
		x"4d",	--1353
		x"4f",	--1354
		x"93",	--1355
		x"28",	--1356
		x"4e",	--1357
		x"93",	--1358
		x"28",	--1359
		x"92",	--1360
		x"20",	--1361
		x"40",	--1362
		x"ec",	--1363
		x"92",	--1364
		x"24",	--1365
		x"93",	--1366
		x"24",	--1367
		x"93",	--1368
		x"24",	--1369
		x"4f",	--1370
		x"00",	--1371
		x"00",	--1372
		x"4e",	--1373
		x"00",	--1374
		x"4f",	--1375
		x"00",	--1376
		x"4f",	--1377
		x"00",	--1378
		x"4e",	--1379
		x"00",	--1380
		x"4e",	--1381
		x"00",	--1382
		x"41",	--1383
		x"8b",	--1384
		x"4c",	--1385
		x"93",	--1386
		x"38",	--1387
		x"90",	--1388
		x"00",	--1389
		x"34",	--1390
		x"93",	--1391
		x"38",	--1392
		x"46",	--1393
		x"00",	--1394
		x"47",	--1395
		x"00",	--1396
		x"49",	--1397
		x"f0",	--1398
		x"00",	--1399
		x"24",	--1400
		x"46",	--1401
		x"47",	--1402
		x"c3",	--1403
		x"10",	--1404
		x"10",	--1405
		x"53",	--1406
		x"23",	--1407
		x"4a",	--1408
		x"00",	--1409
		x"4b",	--1410
		x"00",	--1411
		x"43",	--1412
		x"43",	--1413
		x"f0",	--1414
		x"00",	--1415
		x"24",	--1416
		x"5c",	--1417
		x"6d",	--1418
		x"53",	--1419
		x"23",	--1420
		x"53",	--1421
		x"63",	--1422
		x"f6",	--1423
		x"f7",	--1424
		x"43",	--1425
		x"43",	--1426
		x"93",	--1427
		x"20",	--1428
		x"93",	--1429
		x"24",	--1430
		x"41",	--1431
		x"00",	--1432
		x"41",	--1433
		x"00",	--1434
		x"da",	--1435
		x"db",	--1436
		x"4f",	--1437
		x"00",	--1438
		x"9e",	--1439
		x"00",	--1440
		x"20",	--1441
		x"4f",	--1442
		x"00",	--1443
		x"41",	--1444
		x"00",	--1445
		x"46",	--1446
		x"47",	--1447
		x"54",	--1448
		x"65",	--1449
		x"4e",	--1450
		x"00",	--1451
		x"4f",	--1452
		x"00",	--1453
		x"40",	--1454
		x"00",	--1455
		x"00",	--1456
		x"93",	--1457
		x"38",	--1458
		x"48",	--1459
		x"50",	--1460
		x"00",	--1461
		x"41",	--1462
		x"41",	--1463
		x"41",	--1464
		x"41",	--1465
		x"41",	--1466
		x"41",	--1467
		x"41",	--1468
		x"41",	--1469
		x"41",	--1470
		x"91",	--1471
		x"38",	--1472
		x"4b",	--1473
		x"00",	--1474
		x"43",	--1475
		x"43",	--1476
		x"4f",	--1477
		x"00",	--1478
		x"9e",	--1479
		x"00",	--1480
		x"27",	--1481
		x"93",	--1482
		x"24",	--1483
		x"46",	--1484
		x"47",	--1485
		x"84",	--1486
		x"75",	--1487
		x"93",	--1488
		x"38",	--1489
		x"43",	--1490
		x"00",	--1491
		x"41",	--1492
		x"00",	--1493
		x"4e",	--1494
		x"00",	--1495
		x"4f",	--1496
		x"00",	--1497
		x"4e",	--1498
		x"4f",	--1499
		x"53",	--1500
		x"63",	--1501
		x"90",	--1502
		x"3f",	--1503
		x"28",	--1504
		x"90",	--1505
		x"40",	--1506
		x"2c",	--1507
		x"93",	--1508
		x"2c",	--1509
		x"48",	--1510
		x"00",	--1511
		x"53",	--1512
		x"5e",	--1513
		x"6f",	--1514
		x"4b",	--1515
		x"53",	--1516
		x"4e",	--1517
		x"4f",	--1518
		x"53",	--1519
		x"63",	--1520
		x"90",	--1521
		x"3f",	--1522
		x"2b",	--1523
		x"24",	--1524
		x"4e",	--1525
		x"00",	--1526
		x"4f",	--1527
		x"00",	--1528
		x"4a",	--1529
		x"00",	--1530
		x"40",	--1531
		x"00",	--1532
		x"00",	--1533
		x"93",	--1534
		x"37",	--1535
		x"4e",	--1536
		x"4f",	--1537
		x"f3",	--1538
		x"f3",	--1539
		x"c3",	--1540
		x"10",	--1541
		x"10",	--1542
		x"4c",	--1543
		x"4d",	--1544
		x"de",	--1545
		x"df",	--1546
		x"4a",	--1547
		x"00",	--1548
		x"4b",	--1549
		x"00",	--1550
		x"53",	--1551
		x"00",	--1552
		x"48",	--1553
		x"3f",	--1554
		x"93",	--1555
		x"23",	--1556
		x"4f",	--1557
		x"00",	--1558
		x"4f",	--1559
		x"00",	--1560
		x"00",	--1561
		x"4f",	--1562
		x"00",	--1563
		x"00",	--1564
		x"4f",	--1565
		x"00",	--1566
		x"00",	--1567
		x"4e",	--1568
		x"00",	--1569
		x"ff",	--1570
		x"00",	--1571
		x"4e",	--1572
		x"00",	--1573
		x"4d",	--1574
		x"3f",	--1575
		x"43",	--1576
		x"43",	--1577
		x"3f",	--1578
		x"e3",	--1579
		x"53",	--1580
		x"90",	--1581
		x"00",	--1582
		x"37",	--1583
		x"3f",	--1584
		x"93",	--1585
		x"2b",	--1586
		x"3f",	--1587
		x"44",	--1588
		x"45",	--1589
		x"86",	--1590
		x"77",	--1591
		x"3f",	--1592
		x"4e",	--1593
		x"3f",	--1594
		x"43",	--1595
		x"00",	--1596
		x"41",	--1597
		x"00",	--1598
		x"e3",	--1599
		x"e3",	--1600
		x"53",	--1601
		x"63",	--1602
		x"4e",	--1603
		x"00",	--1604
		x"4f",	--1605
		x"00",	--1606
		x"3f",	--1607
		x"93",	--1608
		x"27",	--1609
		x"59",	--1610
		x"00",	--1611
		x"44",	--1612
		x"00",	--1613
		x"45",	--1614
		x"00",	--1615
		x"49",	--1616
		x"f0",	--1617
		x"00",	--1618
		x"24",	--1619
		x"4d",	--1620
		x"44",	--1621
		x"45",	--1622
		x"c3",	--1623
		x"10",	--1624
		x"10",	--1625
		x"53",	--1626
		x"23",	--1627
		x"4c",	--1628
		x"00",	--1629
		x"4d",	--1630
		x"00",	--1631
		x"43",	--1632
		x"43",	--1633
		x"f0",	--1634
		x"00",	--1635
		x"24",	--1636
		x"5c",	--1637
		x"6d",	--1638
		x"53",	--1639
		x"23",	--1640
		x"53",	--1641
		x"63",	--1642
		x"f4",	--1643
		x"f5",	--1644
		x"43",	--1645
		x"43",	--1646
		x"93",	--1647
		x"20",	--1648
		x"93",	--1649
		x"20",	--1650
		x"43",	--1651
		x"43",	--1652
		x"41",	--1653
		x"00",	--1654
		x"41",	--1655
		x"00",	--1656
		x"da",	--1657
		x"db",	--1658
		x"3f",	--1659
		x"43",	--1660
		x"43",	--1661
		x"3f",	--1662
		x"92",	--1663
		x"23",	--1664
		x"9e",	--1665
		x"00",	--1666
		x"00",	--1667
		x"27",	--1668
		x"40",	--1669
		x"fa",	--1670
		x"3f",	--1671
		x"50",	--1672
		x"ff",	--1673
		x"4e",	--1674
		x"00",	--1675
		x"4f",	--1676
		x"00",	--1677
		x"4c",	--1678
		x"00",	--1679
		x"4d",	--1680
		x"00",	--1681
		x"41",	--1682
		x"50",	--1683
		x"00",	--1684
		x"41",	--1685
		x"52",	--1686
		x"12",	--1687
		x"f5",	--1688
		x"41",	--1689
		x"50",	--1690
		x"00",	--1691
		x"41",	--1692
		x"12",	--1693
		x"f5",	--1694
		x"41",	--1695
		x"52",	--1696
		x"41",	--1697
		x"50",	--1698
		x"00",	--1699
		x"41",	--1700
		x"50",	--1701
		x"00",	--1702
		x"12",	--1703
		x"ea",	--1704
		x"12",	--1705
		x"f3",	--1706
		x"50",	--1707
		x"00",	--1708
		x"41",	--1709
		x"50",	--1710
		x"ff",	--1711
		x"4e",	--1712
		x"00",	--1713
		x"4f",	--1714
		x"00",	--1715
		x"4c",	--1716
		x"00",	--1717
		x"4d",	--1718
		x"00",	--1719
		x"41",	--1720
		x"50",	--1721
		x"00",	--1722
		x"41",	--1723
		x"52",	--1724
		x"12",	--1725
		x"f5",	--1726
		x"41",	--1727
		x"50",	--1728
		x"00",	--1729
		x"41",	--1730
		x"12",	--1731
		x"f5",	--1732
		x"e3",	--1733
		x"00",	--1734
		x"41",	--1735
		x"52",	--1736
		x"41",	--1737
		x"50",	--1738
		x"00",	--1739
		x"41",	--1740
		x"50",	--1741
		x"00",	--1742
		x"12",	--1743
		x"ea",	--1744
		x"12",	--1745
		x"f3",	--1746
		x"50",	--1747
		x"00",	--1748
		x"41",	--1749
		x"12",	--1750
		x"12",	--1751
		x"12",	--1752
		x"12",	--1753
		x"12",	--1754
		x"12",	--1755
		x"12",	--1756
		x"12",	--1757
		x"50",	--1758
		x"ff",	--1759
		x"4e",	--1760
		x"00",	--1761
		x"4f",	--1762
		x"00",	--1763
		x"4c",	--1764
		x"00",	--1765
		x"4d",	--1766
		x"00",	--1767
		x"41",	--1768
		x"50",	--1769
		x"00",	--1770
		x"41",	--1771
		x"52",	--1772
		x"12",	--1773
		x"f5",	--1774
		x"41",	--1775
		x"50",	--1776
		x"00",	--1777
		x"41",	--1778
		x"12",	--1779
		x"f5",	--1780
		x"41",	--1781
		x"00",	--1782
		x"93",	--1783
		x"28",	--1784
		x"41",	--1785
		x"00",	--1786
		x"93",	--1787
		x"28",	--1788
		x"92",	--1789
		x"24",	--1790
		x"92",	--1791
		x"24",	--1792
		x"93",	--1793
		x"24",	--1794
		x"93",	--1795
		x"24",	--1796
		x"41",	--1797
		x"00",	--1798
		x"41",	--1799
		x"00",	--1800
		x"41",	--1801
		x"00",	--1802
		x"41",	--1803
		x"00",	--1804
		x"40",	--1805
		x"00",	--1806
		x"43",	--1807
		x"43",	--1808
		x"43",	--1809
		x"43",	--1810
		x"43",	--1811
		x"00",	--1812
		x"43",	--1813
		x"00",	--1814
		x"43",	--1815
		x"43",	--1816
		x"4c",	--1817
		x"00",	--1818
		x"3c",	--1819
		x"58",	--1820
		x"69",	--1821
		x"c3",	--1822
		x"10",	--1823
		x"10",	--1824
		x"53",	--1825
		x"00",	--1826
		x"24",	--1827
		x"b3",	--1828
		x"24",	--1829
		x"58",	--1830
		x"69",	--1831
		x"56",	--1832
		x"67",	--1833
		x"43",	--1834
		x"43",	--1835
		x"99",	--1836
		x"28",	--1837
		x"24",	--1838
		x"43",	--1839
		x"43",	--1840
		x"5c",	--1841
		x"6d",	--1842
		x"56",	--1843
		x"67",	--1844
		x"93",	--1845
		x"37",	--1846
		x"d3",	--1847
		x"d3",	--1848
		x"3f",	--1849
		x"98",	--1850
		x"2b",	--1851
		x"3f",	--1852
		x"4a",	--1853
		x"00",	--1854
		x"4b",	--1855
		x"00",	--1856
		x"4f",	--1857
		x"41",	--1858
		x"00",	--1859
		x"51",	--1860
		x"00",	--1861
		x"4a",	--1862
		x"53",	--1863
		x"46",	--1864
		x"00",	--1865
		x"43",	--1866
		x"91",	--1867
		x"00",	--1868
		x"00",	--1869
		x"24",	--1870
		x"4d",	--1871
		x"00",	--1872
		x"93",	--1873
		x"38",	--1874
		x"90",	--1875
		x"40",	--1876
		x"2c",	--1877
		x"41",	--1878
		x"00",	--1879
		x"53",	--1880
		x"41",	--1881
		x"00",	--1882
		x"41",	--1883
		x"00",	--1884
		x"4d",	--1885
		x"5e",	--1886
		x"6f",	--1887
		x"93",	--1888
		x"38",	--1889
		x"5a",	--1890
		x"6b",	--1891
		x"53",	--1892
		x"90",	--1893
		x"40",	--1894
		x"2b",	--1895
		x"4a",	--1896
		x"00",	--1897
		x"4b",	--1898
		x"00",	--1899
		x"4c",	--1900
		x"00",	--1901
		x"4e",	--1902
		x"4f",	--1903
		x"f0",	--1904
		x"00",	--1905
		x"f3",	--1906
		x"90",	--1907
		x"00",	--1908
		x"24",	--1909
		x"4e",	--1910
		x"00",	--1911
		x"4f",	--1912
		x"00",	--1913
		x"40",	--1914
		x"00",	--1915
		x"00",	--1916
		x"41",	--1917
		x"52",	--1918
		x"12",	--1919
		x"f3",	--1920
		x"50",	--1921
		x"00",	--1922
		x"41",	--1923
		x"41",	--1924
		x"41",	--1925
		x"41",	--1926
		x"41",	--1927
		x"41",	--1928
		x"41",	--1929
		x"41",	--1930
		x"41",	--1931
		x"d3",	--1932
		x"d3",	--1933
		x"3f",	--1934
		x"50",	--1935
		x"00",	--1936
		x"4a",	--1937
		x"b3",	--1938
		x"24",	--1939
		x"41",	--1940
		x"00",	--1941
		x"41",	--1942
		x"00",	--1943
		x"c3",	--1944
		x"10",	--1945
		x"10",	--1946
		x"4c",	--1947
		x"4d",	--1948
		x"d3",	--1949
		x"d0",	--1950
		x"80",	--1951
		x"46",	--1952
		x"00",	--1953
		x"47",	--1954
		x"00",	--1955
		x"c3",	--1956
		x"10",	--1957
		x"10",	--1958
		x"53",	--1959
		x"93",	--1960
		x"3b",	--1961
		x"48",	--1962
		x"00",	--1963
		x"3f",	--1964
		x"93",	--1965
		x"24",	--1966
		x"43",	--1967
		x"91",	--1968
		x"00",	--1969
		x"00",	--1970
		x"24",	--1971
		x"4f",	--1972
		x"00",	--1973
		x"41",	--1974
		x"50",	--1975
		x"00",	--1976
		x"3f",	--1977
		x"93",	--1978
		x"23",	--1979
		x"4e",	--1980
		x"4f",	--1981
		x"f0",	--1982
		x"00",	--1983
		x"f3",	--1984
		x"93",	--1985
		x"23",	--1986
		x"93",	--1987
		x"23",	--1988
		x"93",	--1989
		x"00",	--1990
		x"20",	--1991
		x"93",	--1992
		x"00",	--1993
		x"27",	--1994
		x"50",	--1995
		x"00",	--1996
		x"63",	--1997
		x"f0",	--1998
		x"ff",	--1999
		x"f3",	--2000
		x"3f",	--2001
		x"43",	--2002
		x"3f",	--2003
		x"43",	--2004
		x"3f",	--2005
		x"43",	--2006
		x"91",	--2007
		x"00",	--2008
		x"00",	--2009
		x"24",	--2010
		x"4f",	--2011
		x"00",	--2012
		x"41",	--2013
		x"50",	--2014
		x"00",	--2015
		x"3f",	--2016
		x"43",	--2017
		x"3f",	--2018
		x"93",	--2019
		x"23",	--2020
		x"40",	--2021
		x"fa",	--2022
		x"3f",	--2023
		x"12",	--2024
		x"12",	--2025
		x"12",	--2026
		x"12",	--2027
		x"12",	--2028
		x"50",	--2029
		x"ff",	--2030
		x"4e",	--2031
		x"00",	--2032
		x"4f",	--2033
		x"00",	--2034
		x"4c",	--2035
		x"00",	--2036
		x"4d",	--2037
		x"00",	--2038
		x"41",	--2039
		x"50",	--2040
		x"00",	--2041
		x"41",	--2042
		x"52",	--2043
		x"12",	--2044
		x"f5",	--2045
		x"41",	--2046
		x"52",	--2047
		x"41",	--2048
		x"12",	--2049
		x"f5",	--2050
		x"41",	--2051
		x"00",	--2052
		x"93",	--2053
		x"28",	--2054
		x"41",	--2055
		x"00",	--2056
		x"93",	--2057
		x"28",	--2058
		x"e1",	--2059
		x"00",	--2060
		x"00",	--2061
		x"92",	--2062
		x"24",	--2063
		x"93",	--2064
		x"24",	--2065
		x"92",	--2066
		x"24",	--2067
		x"93",	--2068
		x"24",	--2069
		x"41",	--2070
		x"00",	--2071
		x"81",	--2072
		x"00",	--2073
		x"4d",	--2074
		x"00",	--2075
		x"41",	--2076
		x"00",	--2077
		x"41",	--2078
		x"00",	--2079
		x"41",	--2080
		x"00",	--2081
		x"41",	--2082
		x"00",	--2083
		x"99",	--2084
		x"2c",	--2085
		x"5e",	--2086
		x"6f",	--2087
		x"53",	--2088
		x"4d",	--2089
		x"00",	--2090
		x"40",	--2091
		x"00",	--2092
		x"43",	--2093
		x"40",	--2094
		x"40",	--2095
		x"43",	--2096
		x"43",	--2097
		x"3c",	--2098
		x"dc",	--2099
		x"dd",	--2100
		x"88",	--2101
		x"79",	--2102
		x"c3",	--2103
		x"10",	--2104
		x"10",	--2105
		x"5e",	--2106
		x"6f",	--2107
		x"53",	--2108
		x"24",	--2109
		x"99",	--2110
		x"2b",	--2111
		x"23",	--2112
		x"98",	--2113
		x"2b",	--2114
		x"3f",	--2115
		x"9f",	--2116
		x"2b",	--2117
		x"98",	--2118
		x"2f",	--2119
		x"3f",	--2120
		x"4a",	--2121
		x"4b",	--2122
		x"f0",	--2123
		x"00",	--2124
		x"f3",	--2125
		x"90",	--2126
		x"00",	--2127
		x"24",	--2128
		x"4a",	--2129
		x"00",	--2130
		x"4b",	--2131
		x"00",	--2132
		x"41",	--2133
		x"50",	--2134
		x"00",	--2135
		x"12",	--2136
		x"f3",	--2137
		x"50",	--2138
		x"00",	--2139
		x"41",	--2140
		x"41",	--2141
		x"41",	--2142
		x"41",	--2143
		x"41",	--2144
		x"41",	--2145
		x"42",	--2146
		x"00",	--2147
		x"41",	--2148
		x"50",	--2149
		x"00",	--2150
		x"3f",	--2151
		x"9e",	--2152
		x"23",	--2153
		x"40",	--2154
		x"fa",	--2155
		x"3f",	--2156
		x"93",	--2157
		x"23",	--2158
		x"4a",	--2159
		x"4b",	--2160
		x"f0",	--2161
		x"00",	--2162
		x"f3",	--2163
		x"93",	--2164
		x"23",	--2165
		x"93",	--2166
		x"23",	--2167
		x"93",	--2168
		x"20",	--2169
		x"93",	--2170
		x"27",	--2171
		x"50",	--2172
		x"00",	--2173
		x"63",	--2174
		x"f0",	--2175
		x"ff",	--2176
		x"f3",	--2177
		x"3f",	--2178
		x"43",	--2179
		x"00",	--2180
		x"43",	--2181
		x"00",	--2182
		x"43",	--2183
		x"00",	--2184
		x"41",	--2185
		x"50",	--2186
		x"00",	--2187
		x"3f",	--2188
		x"41",	--2189
		x"52",	--2190
		x"3f",	--2191
		x"50",	--2192
		x"ff",	--2193
		x"4e",	--2194
		x"00",	--2195
		x"4f",	--2196
		x"00",	--2197
		x"4c",	--2198
		x"00",	--2199
		x"4d",	--2200
		x"00",	--2201
		x"41",	--2202
		x"50",	--2203
		x"00",	--2204
		x"41",	--2205
		x"52",	--2206
		x"12",	--2207
		x"f5",	--2208
		x"41",	--2209
		x"52",	--2210
		x"41",	--2211
		x"12",	--2212
		x"f5",	--2213
		x"93",	--2214
		x"00",	--2215
		x"28",	--2216
		x"93",	--2217
		x"00",	--2218
		x"28",	--2219
		x"41",	--2220
		x"52",	--2221
		x"41",	--2222
		x"50",	--2223
		x"00",	--2224
		x"12",	--2225
		x"f6",	--2226
		x"50",	--2227
		x"00",	--2228
		x"41",	--2229
		x"43",	--2230
		x"3f",	--2231
		x"50",	--2232
		x"ff",	--2233
		x"4e",	--2234
		x"00",	--2235
		x"4f",	--2236
		x"00",	--2237
		x"41",	--2238
		x"52",	--2239
		x"41",	--2240
		x"12",	--2241
		x"f5",	--2242
		x"41",	--2243
		x"00",	--2244
		x"93",	--2245
		x"24",	--2246
		x"28",	--2247
		x"92",	--2248
		x"24",	--2249
		x"41",	--2250
		x"00",	--2251
		x"93",	--2252
		x"38",	--2253
		x"90",	--2254
		x"00",	--2255
		x"38",	--2256
		x"93",	--2257
		x"00",	--2258
		x"20",	--2259
		x"43",	--2260
		x"40",	--2261
		x"7f",	--2262
		x"50",	--2263
		x"00",	--2264
		x"41",	--2265
		x"41",	--2266
		x"00",	--2267
		x"41",	--2268
		x"00",	--2269
		x"40",	--2270
		x"00",	--2271
		x"8d",	--2272
		x"4c",	--2273
		x"f0",	--2274
		x"00",	--2275
		x"20",	--2276
		x"93",	--2277
		x"00",	--2278
		x"27",	--2279
		x"e3",	--2280
		x"e3",	--2281
		x"53",	--2282
		x"63",	--2283
		x"50",	--2284
		x"00",	--2285
		x"41",	--2286
		x"43",	--2287
		x"43",	--2288
		x"50",	--2289
		x"00",	--2290
		x"41",	--2291
		x"c3",	--2292
		x"10",	--2293
		x"10",	--2294
		x"53",	--2295
		x"23",	--2296
		x"3f",	--2297
		x"43",	--2298
		x"40",	--2299
		x"80",	--2300
		x"50",	--2301
		x"00",	--2302
		x"41",	--2303
		x"12",	--2304
		x"12",	--2305
		x"12",	--2306
		x"12",	--2307
		x"82",	--2308
		x"4e",	--2309
		x"4f",	--2310
		x"43",	--2311
		x"00",	--2312
		x"93",	--2313
		x"20",	--2314
		x"93",	--2315
		x"20",	--2316
		x"43",	--2317
		x"00",	--2318
		x"41",	--2319
		x"12",	--2320
		x"f3",	--2321
		x"52",	--2322
		x"41",	--2323
		x"41",	--2324
		x"41",	--2325
		x"41",	--2326
		x"41",	--2327
		x"40",	--2328
		x"00",	--2329
		x"00",	--2330
		x"40",	--2331
		x"00",	--2332
		x"00",	--2333
		x"4a",	--2334
		x"00",	--2335
		x"4b",	--2336
		x"00",	--2337
		x"4a",	--2338
		x"4b",	--2339
		x"12",	--2340
		x"f2",	--2341
		x"53",	--2342
		x"93",	--2343
		x"38",	--2344
		x"27",	--2345
		x"4a",	--2346
		x"00",	--2347
		x"4b",	--2348
		x"00",	--2349
		x"4f",	--2350
		x"f0",	--2351
		x"00",	--2352
		x"20",	--2353
		x"40",	--2354
		x"00",	--2355
		x"8f",	--2356
		x"4e",	--2357
		x"00",	--2358
		x"3f",	--2359
		x"51",	--2360
		x"00",	--2361
		x"00",	--2362
		x"61",	--2363
		x"00",	--2364
		x"00",	--2365
		x"53",	--2366
		x"23",	--2367
		x"3f",	--2368
		x"4f",	--2369
		x"e3",	--2370
		x"53",	--2371
		x"43",	--2372
		x"43",	--2373
		x"4e",	--2374
		x"f0",	--2375
		x"00",	--2376
		x"24",	--2377
		x"5c",	--2378
		x"6d",	--2379
		x"53",	--2380
		x"23",	--2381
		x"53",	--2382
		x"63",	--2383
		x"fa",	--2384
		x"fb",	--2385
		x"43",	--2386
		x"43",	--2387
		x"93",	--2388
		x"20",	--2389
		x"93",	--2390
		x"20",	--2391
		x"43",	--2392
		x"43",	--2393
		x"f0",	--2394
		x"00",	--2395
		x"20",	--2396
		x"48",	--2397
		x"49",	--2398
		x"da",	--2399
		x"db",	--2400
		x"4d",	--2401
		x"00",	--2402
		x"4e",	--2403
		x"00",	--2404
		x"40",	--2405
		x"00",	--2406
		x"8f",	--2407
		x"4e",	--2408
		x"00",	--2409
		x"3f",	--2410
		x"c3",	--2411
		x"10",	--2412
		x"10",	--2413
		x"53",	--2414
		x"23",	--2415
		x"3f",	--2416
		x"12",	--2417
		x"12",	--2418
		x"12",	--2419
		x"93",	--2420
		x"2c",	--2421
		x"90",	--2422
		x"01",	--2423
		x"28",	--2424
		x"40",	--2425
		x"00",	--2426
		x"43",	--2427
		x"42",	--2428
		x"4e",	--2429
		x"4f",	--2430
		x"49",	--2431
		x"93",	--2432
		x"20",	--2433
		x"50",	--2434
		x"fa",	--2435
		x"4c",	--2436
		x"43",	--2437
		x"8e",	--2438
		x"7f",	--2439
		x"4a",	--2440
		x"41",	--2441
		x"41",	--2442
		x"41",	--2443
		x"41",	--2444
		x"90",	--2445
		x"01",	--2446
		x"28",	--2447
		x"42",	--2448
		x"43",	--2449
		x"40",	--2450
		x"00",	--2451
		x"4e",	--2452
		x"4f",	--2453
		x"49",	--2454
		x"93",	--2455
		x"27",	--2456
		x"c3",	--2457
		x"10",	--2458
		x"10",	--2459
		x"53",	--2460
		x"23",	--2461
		x"3f",	--2462
		x"40",	--2463
		x"00",	--2464
		x"43",	--2465
		x"40",	--2466
		x"00",	--2467
		x"3f",	--2468
		x"40",	--2469
		x"00",	--2470
		x"43",	--2471
		x"43",	--2472
		x"3f",	--2473
		x"12",	--2474
		x"12",	--2475
		x"12",	--2476
		x"12",	--2477
		x"12",	--2478
		x"4f",	--2479
		x"4f",	--2480
		x"00",	--2481
		x"4f",	--2482
		x"00",	--2483
		x"4d",	--2484
		x"00",	--2485
		x"4d",	--2486
		x"93",	--2487
		x"28",	--2488
		x"92",	--2489
		x"24",	--2490
		x"93",	--2491
		x"24",	--2492
		x"93",	--2493
		x"24",	--2494
		x"4d",	--2495
		x"00",	--2496
		x"90",	--2497
		x"ff",	--2498
		x"38",	--2499
		x"90",	--2500
		x"00",	--2501
		x"34",	--2502
		x"4e",	--2503
		x"4f",	--2504
		x"f0",	--2505
		x"00",	--2506
		x"f3",	--2507
		x"90",	--2508
		x"00",	--2509
		x"24",	--2510
		x"50",	--2511
		x"00",	--2512
		x"63",	--2513
		x"93",	--2514
		x"38",	--2515
		x"4b",	--2516
		x"50",	--2517
		x"00",	--2518
		x"c3",	--2519
		x"10",	--2520
		x"10",	--2521
		x"c3",	--2522
		x"10",	--2523
		x"10",	--2524
		x"c3",	--2525
		x"10",	--2526
		x"10",	--2527
		x"c3",	--2528
		x"10",	--2529
		x"10",	--2530
		x"c3",	--2531
		x"10",	--2532
		x"10",	--2533
		x"c3",	--2534
		x"10",	--2535
		x"10",	--2536
		x"c3",	--2537
		x"10",	--2538
		x"10",	--2539
		x"f3",	--2540
		x"f0",	--2541
		x"00",	--2542
		x"4d",	--2543
		x"3c",	--2544
		x"93",	--2545
		x"23",	--2546
		x"43",	--2547
		x"43",	--2548
		x"43",	--2549
		x"4d",	--2550
		x"5d",	--2551
		x"5d",	--2552
		x"5d",	--2553
		x"5d",	--2554
		x"5d",	--2555
		x"5d",	--2556
		x"5d",	--2557
		x"4f",	--2558
		x"f0",	--2559
		x"00",	--2560
		x"dd",	--2561
		x"4a",	--2562
		x"11",	--2563
		x"43",	--2564
		x"10",	--2565
		x"4c",	--2566
		x"df",	--2567
		x"4d",	--2568
		x"41",	--2569
		x"41",	--2570
		x"41",	--2571
		x"41",	--2572
		x"41",	--2573
		x"41",	--2574
		x"93",	--2575
		x"23",	--2576
		x"4e",	--2577
		x"4f",	--2578
		x"f0",	--2579
		x"00",	--2580
		x"f3",	--2581
		x"93",	--2582
		x"20",	--2583
		x"93",	--2584
		x"27",	--2585
		x"50",	--2586
		x"00",	--2587
		x"63",	--2588
		x"3f",	--2589
		x"c3",	--2590
		x"10",	--2591
		x"10",	--2592
		x"4b",	--2593
		x"50",	--2594
		x"00",	--2595
		x"3f",	--2596
		x"43",	--2597
		x"43",	--2598
		x"43",	--2599
		x"3f",	--2600
		x"d3",	--2601
		x"d0",	--2602
		x"00",	--2603
		x"f3",	--2604
		x"f0",	--2605
		x"00",	--2606
		x"43",	--2607
		x"3f",	--2608
		x"40",	--2609
		x"ff",	--2610
		x"8b",	--2611
		x"90",	--2612
		x"00",	--2613
		x"34",	--2614
		x"4e",	--2615
		x"4f",	--2616
		x"47",	--2617
		x"f0",	--2618
		x"00",	--2619
		x"24",	--2620
		x"c3",	--2621
		x"10",	--2622
		x"10",	--2623
		x"53",	--2624
		x"23",	--2625
		x"43",	--2626
		x"43",	--2627
		x"f0",	--2628
		x"00",	--2629
		x"24",	--2630
		x"58",	--2631
		x"69",	--2632
		x"53",	--2633
		x"23",	--2634
		x"53",	--2635
		x"63",	--2636
		x"fe",	--2637
		x"ff",	--2638
		x"43",	--2639
		x"43",	--2640
		x"93",	--2641
		x"20",	--2642
		x"93",	--2643
		x"20",	--2644
		x"43",	--2645
		x"43",	--2646
		x"4e",	--2647
		x"4f",	--2648
		x"dc",	--2649
		x"dd",	--2650
		x"48",	--2651
		x"49",	--2652
		x"f0",	--2653
		x"00",	--2654
		x"f3",	--2655
		x"90",	--2656
		x"00",	--2657
		x"24",	--2658
		x"50",	--2659
		x"00",	--2660
		x"63",	--2661
		x"48",	--2662
		x"49",	--2663
		x"c3",	--2664
		x"10",	--2665
		x"10",	--2666
		x"c3",	--2667
		x"10",	--2668
		x"10",	--2669
		x"c3",	--2670
		x"10",	--2671
		x"10",	--2672
		x"c3",	--2673
		x"10",	--2674
		x"10",	--2675
		x"c3",	--2676
		x"10",	--2677
		x"10",	--2678
		x"c3",	--2679
		x"10",	--2680
		x"10",	--2681
		x"c3",	--2682
		x"10",	--2683
		x"10",	--2684
		x"f3",	--2685
		x"f0",	--2686
		x"00",	--2687
		x"43",	--2688
		x"90",	--2689
		x"40",	--2690
		x"2f",	--2691
		x"43",	--2692
		x"3f",	--2693
		x"43",	--2694
		x"43",	--2695
		x"3f",	--2696
		x"93",	--2697
		x"23",	--2698
		x"48",	--2699
		x"49",	--2700
		x"f0",	--2701
		x"00",	--2702
		x"f3",	--2703
		x"93",	--2704
		x"24",	--2705
		x"50",	--2706
		x"00",	--2707
		x"63",	--2708
		x"3f",	--2709
		x"93",	--2710
		x"27",	--2711
		x"3f",	--2712
		x"12",	--2713
		x"12",	--2714
		x"4f",	--2715
		x"4f",	--2716
		x"00",	--2717
		x"f0",	--2718
		x"00",	--2719
		x"4f",	--2720
		x"00",	--2721
		x"c3",	--2722
		x"10",	--2723
		x"c3",	--2724
		x"10",	--2725
		x"c3",	--2726
		x"10",	--2727
		x"c3",	--2728
		x"10",	--2729
		x"c3",	--2730
		x"10",	--2731
		x"c3",	--2732
		x"10",	--2733
		x"c3",	--2734
		x"10",	--2735
		x"4d",	--2736
		x"4f",	--2737
		x"00",	--2738
		x"b0",	--2739
		x"00",	--2740
		x"43",	--2741
		x"6f",	--2742
		x"4f",	--2743
		x"00",	--2744
		x"93",	--2745
		x"20",	--2746
		x"93",	--2747
		x"24",	--2748
		x"40",	--2749
		x"ff",	--2750
		x"00",	--2751
		x"4a",	--2752
		x"4b",	--2753
		x"5c",	--2754
		x"6d",	--2755
		x"5c",	--2756
		x"6d",	--2757
		x"5c",	--2758
		x"6d",	--2759
		x"5c",	--2760
		x"6d",	--2761
		x"5c",	--2762
		x"6d",	--2763
		x"5c",	--2764
		x"6d",	--2765
		x"5c",	--2766
		x"6d",	--2767
		x"40",	--2768
		x"00",	--2769
		x"00",	--2770
		x"90",	--2771
		x"40",	--2772
		x"2c",	--2773
		x"40",	--2774
		x"ff",	--2775
		x"5c",	--2776
		x"6d",	--2777
		x"4f",	--2778
		x"53",	--2779
		x"90",	--2780
		x"40",	--2781
		x"2b",	--2782
		x"4a",	--2783
		x"00",	--2784
		x"4c",	--2785
		x"00",	--2786
		x"4d",	--2787
		x"00",	--2788
		x"41",	--2789
		x"41",	--2790
		x"41",	--2791
		x"90",	--2792
		x"00",	--2793
		x"24",	--2794
		x"50",	--2795
		x"ff",	--2796
		x"4d",	--2797
		x"00",	--2798
		x"40",	--2799
		x"00",	--2800
		x"00",	--2801
		x"4a",	--2802
		x"4b",	--2803
		x"5c",	--2804
		x"6d",	--2805
		x"5c",	--2806
		x"6d",	--2807
		x"5c",	--2808
		x"6d",	--2809
		x"5c",	--2810
		x"6d",	--2811
		x"5c",	--2812
		x"6d",	--2813
		x"5c",	--2814
		x"6d",	--2815
		x"5c",	--2816
		x"6d",	--2817
		x"4c",	--2818
		x"4d",	--2819
		x"d3",	--2820
		x"d0",	--2821
		x"40",	--2822
		x"4a",	--2823
		x"00",	--2824
		x"4b",	--2825
		x"00",	--2826
		x"41",	--2827
		x"41",	--2828
		x"41",	--2829
		x"93",	--2830
		x"23",	--2831
		x"43",	--2832
		x"00",	--2833
		x"41",	--2834
		x"41",	--2835
		x"41",	--2836
		x"93",	--2837
		x"24",	--2838
		x"4a",	--2839
		x"4b",	--2840
		x"f3",	--2841
		x"f0",	--2842
		x"00",	--2843
		x"93",	--2844
		x"20",	--2845
		x"93",	--2846
		x"24",	--2847
		x"43",	--2848
		x"00",	--2849
		x"3f",	--2850
		x"93",	--2851
		x"23",	--2852
		x"42",	--2853
		x"00",	--2854
		x"3f",	--2855
		x"43",	--2856
		x"00",	--2857
		x"3f",	--2858
		x"12",	--2859
		x"4f",	--2860
		x"93",	--2861
		x"28",	--2862
		x"4e",	--2863
		x"93",	--2864
		x"28",	--2865
		x"92",	--2866
		x"24",	--2867
		x"92",	--2868
		x"24",	--2869
		x"93",	--2870
		x"24",	--2871
		x"93",	--2872
		x"24",	--2873
		x"4f",	--2874
		x"00",	--2875
		x"9e",	--2876
		x"00",	--2877
		x"24",	--2878
		x"93",	--2879
		x"20",	--2880
		x"43",	--2881
		x"4e",	--2882
		x"41",	--2883
		x"41",	--2884
		x"93",	--2885
		x"24",	--2886
		x"93",	--2887
		x"00",	--2888
		x"23",	--2889
		x"43",	--2890
		x"4e",	--2891
		x"41",	--2892
		x"41",	--2893
		x"93",	--2894
		x"00",	--2895
		x"27",	--2896
		x"43",	--2897
		x"3f",	--2898
		x"4f",	--2899
		x"00",	--2900
		x"4e",	--2901
		x"00",	--2902
		x"9b",	--2903
		x"3b",	--2904
		x"9c",	--2905
		x"38",	--2906
		x"4f",	--2907
		x"00",	--2908
		x"4f",	--2909
		x"00",	--2910
		x"4e",	--2911
		x"00",	--2912
		x"4e",	--2913
		x"00",	--2914
		x"9f",	--2915
		x"2b",	--2916
		x"9e",	--2917
		x"28",	--2918
		x"9b",	--2919
		x"2b",	--2920
		x"9e",	--2921
		x"28",	--2922
		x"9f",	--2923
		x"28",	--2924
		x"9c",	--2925
		x"28",	--2926
		x"43",	--2927
		x"3f",	--2928
		x"93",	--2929
		x"23",	--2930
		x"43",	--2931
		x"3f",	--2932
		x"92",	--2933
		x"23",	--2934
		x"4e",	--2935
		x"00",	--2936
		x"4f",	--2937
		x"00",	--2938
		x"8f",	--2939
		x"3f",	--2940
		x"43",	--2941
		x"93",	--2942
		x"34",	--2943
		x"40",	--2944
		x"00",	--2945
		x"e3",	--2946
		x"53",	--2947
		x"93",	--2948
		x"34",	--2949
		x"e3",	--2950
		x"e3",	--2951
		x"53",	--2952
		x"12",	--2953
		x"12",	--2954
		x"f7",	--2955
		x"41",	--2956
		x"b3",	--2957
		x"24",	--2958
		x"e3",	--2959
		x"53",	--2960
		x"b3",	--2961
		x"24",	--2962
		x"e3",	--2963
		x"53",	--2964
		x"41",	--2965
		x"12",	--2966
		x"f6",	--2967
		x"4e",	--2968
		x"41",	--2969
		x"12",	--2970
		x"43",	--2971
		x"93",	--2972
		x"34",	--2973
		x"40",	--2974
		x"00",	--2975
		x"e3",	--2976
		x"e3",	--2977
		x"53",	--2978
		x"63",	--2979
		x"93",	--2980
		x"34",	--2981
		x"e3",	--2982
		x"e3",	--2983
		x"e3",	--2984
		x"53",	--2985
		x"63",	--2986
		x"12",	--2987
		x"f7",	--2988
		x"b3",	--2989
		x"24",	--2990
		x"e3",	--2991
		x"e3",	--2992
		x"53",	--2993
		x"63",	--2994
		x"b3",	--2995
		x"24",	--2996
		x"e3",	--2997
		x"e3",	--2998
		x"53",	--2999
		x"63",	--3000
		x"41",	--3001
		x"41",	--3002
		x"12",	--3003
		x"f7",	--3004
		x"4c",	--3005
		x"4d",	--3006
		x"41",	--3007
		x"40",	--3008
		x"00",	--3009
		x"4e",	--3010
		x"43",	--3011
		x"5f",	--3012
		x"6e",	--3013
		x"9d",	--3014
		x"28",	--3015
		x"8d",	--3016
		x"d3",	--3017
		x"83",	--3018
		x"23",	--3019
		x"41",	--3020
		x"12",	--3021
		x"f7",	--3022
		x"4e",	--3023
		x"41",	--3024
		x"12",	--3025
		x"12",	--3026
		x"12",	--3027
		x"40",	--3028
		x"00",	--3029
		x"4c",	--3030
		x"4d",	--3031
		x"43",	--3032
		x"43",	--3033
		x"5e",	--3034
		x"6f",	--3035
		x"6c",	--3036
		x"6d",	--3037
		x"9b",	--3038
		x"28",	--3039
		x"20",	--3040
		x"9a",	--3041
		x"28",	--3042
		x"8a",	--3043
		x"7b",	--3044
		x"d3",	--3045
		x"83",	--3046
		x"23",	--3047
		x"41",	--3048
		x"41",	--3049
		x"41",	--3050
		x"41",	--3051
		x"12",	--3052
		x"f7",	--3053
		x"4c",	--3054
		x"4d",	--3055
		x"41",	--3056
		x"13",	--3057
		x"d0",	--3058
		x"00",	--3059
		x"3f",	--3060
		x"61",	--3061
		x"74",	--3062
		x"6e",	--3063
		x"20",	--3064
		x"6f",	--3065
		x"20",	--3066
		x"20",	--3067
		x"65",	--3068
		x"20",	--3069
		x"62",	--3070
		x"6e",	--3071
		x"66",	--3072
		x"6c",	--3073
		x"0d",	--3074
		x"00",	--3075
		x"65",	--3076
		x"73",	--3077
		x"6f",	--3078
		x"6c",	--3079
		x"20",	--3080
		x"6f",	--3081
		x"20",	--3082
		x"65",	--3083
		x"20",	--3084
		x"68",	--3085
		x"74",	--3086
		x"0a",	--3087
		x"63",	--3088
		x"72",	--3089
		x"65",	--3090
		x"74",	--3091
		x"75",	--3092
		x"61",	--3093
		x"65",	--3094
		x"0d",	--3095
		x"00",	--3096
		x"25",	--3097
		x"20",	--3098
		x"45",	--3099
		x"54",	--3100
		x"52",	--3101
		x"47",	--3102
		x"54",	--3103
		x"0a",	--3104
		x"53",	--3105
		x"6d",	--3106
		x"74",	--3107
		x"69",	--3108
		x"67",	--3109
		x"77",	--3110
		x"6e",	--3111
		x"20",	--3112
		x"65",	--3113
		x"72",	--3114
		x"62",	--3115
		x"79",	--3116
		x"77",	--3117
		x"6f",	--3118
		x"67",	--3119
		x"0a",	--3120
		x"0d",	--3121
		x"3d",	--3122
		x"3d",	--3123
		x"3d",	--3124
		x"20",	--3125
		x"61",	--3126
		x"63",	--3127
		x"6c",	--3128
		x"4d",	--3129
		x"55",	--3130
		x"3d",	--3131
		x"3d",	--3132
		x"3d",	--3133
		x"0d",	--3134
		x"00",	--3135
		x"72",	--3136
		x"74",	--3137
		x"00",	--3138
		x"65",	--3139
		x"64",	--3140
		x"70",	--3141
		x"6d",	--3142
		x"62",	--3143
		x"6f",	--3144
		x"6c",	--3145
		x"61",	--3146
		x"65",	--3147
		x"00",	--3148
		x"20",	--3149
		x"0d",	--3150
		x"00",	--3151
		x"25",	--3152
		x"0d",	--3153
		x"00",	--3154
		x"20",	--3155
		x"00",	--3156
		x"63",	--3157
		x"77",	--3158
		x"69",	--3159
		x"65",	--3160
		x"0d",	--3161
		x"63",	--3162
		x"72",	--3163
		x"65",	--3164
		x"74",	--3165
		x"75",	--3166
		x"61",	--3167
		x"65",	--3168
		x"0d",	--3169
		x"00",	--3170
		x"25",	--3171
		x"20",	--3172
		x"45",	--3173
		x"49",	--3174
		x"54",	--3175
		x"52",	--3176
		x"56",	--3177
		x"4c",	--3178
		x"45",	--3179
		x"0a",	--3180
		x"53",	--3181
		x"6d",	--3182
		x"74",	--3183
		x"69",	--3184
		x"67",	--3185
		x"77",	--3186
		x"6e",	--3187
		x"20",	--3188
		x"65",	--3189
		x"72",	--3190
		x"62",	--3191
		x"79",	--3192
		x"77",	--3193
		x"6f",	--3194
		x"67",	--3195
		x"0a",	--3196
		x"72",	--3197
		x"25",	--3198
		x"20",	--3199
		x"3d",	--3200
		x"64",	--3201
		x"0a",	--3202
		x"72",	--3203
		x"61",	--3204
		x"0a",	--3205
		x"00",	--3206
		x"25",	--3207
		x"20",	--3208
		x"45",	--3209
		x"49",	--3210
		x"54",	--3211
		x"52",	--3212
		x"0a",	--3213
		x"25",	--3214
		x"20",	--3215
		x"73",	--3216
		x"6e",	--3217
		x"74",	--3218
		x"61",	--3219
		x"6e",	--3220
		x"6d",	--3221
		x"65",	--3222
		x"0d",	--3223
		x"00",	--3224
		x"63",	--3225
		x"25",	--3226
		x"0d",	--3227
		x"00",	--3228
		x"63",	--3229
		x"20",	--3230
		x"6f",	--3231
		x"73",	--3232
		x"63",	--3233
		x"20",	--3234
		x"6f",	--3235
		x"6d",	--3236
		x"6e",	--3237
		x"0d",	--3238
		x"00",	--3239
		x"e9",	--3240
		x"e8",	--3241
		x"e8",	--3242
		x"e8",	--3243
		x"e8",	--3244
		x"e8",	--3245
		x"e8",	--3246
		x"e8",	--3247
		x"e8",	--3248
		x"e8",	--3249
		x"e8",	--3250
		x"e8",	--3251
		x"e8",	--3252
		x"e8",	--3253
		x"e8",	--3254
		x"e8",	--3255
		x"e8",	--3256
		x"e8",	--3257
		x"e8",	--3258
		x"e8",	--3259
		x"e8",	--3260
		x"e8",	--3261
		x"e8",	--3262
		x"e8",	--3263
		x"e8",	--3264
		x"e8",	--3265
		x"e8",	--3266
		x"e8",	--3267
		x"e8",	--3268
		x"e9",	--3269
		x"e8",	--3270
		x"e8",	--3271
		x"e8",	--3272
		x"e8",	--3273
		x"e8",	--3274
		x"e8",	--3275
		x"e8",	--3276
		x"e8",	--3277
		x"e8",	--3278
		x"e8",	--3279
		x"e8",	--3280
		x"e8",	--3281
		x"e8",	--3282
		x"e8",	--3283
		x"e8",	--3284
		x"e8",	--3285
		x"e8",	--3286
		x"e8",	--3287
		x"e8",	--3288
		x"e8",	--3289
		x"e8",	--3290
		x"e8",	--3291
		x"e8",	--3292
		x"e8",	--3293
		x"e8",	--3294
		x"e8",	--3295
		x"e8",	--3296
		x"e8",	--3297
		x"e8",	--3298
		x"e8",	--3299
		x"e8",	--3300
		x"e9",	--3301
		x"e9",	--3302
		x"e9",	--3303
		x"e8",	--3304
		x"e8",	--3305
		x"e8",	--3306
		x"e8",	--3307
		x"e8",	--3308
		x"e8",	--3309
		x"e8",	--3310
		x"e9",	--3311
		x"e8",	--3312
		x"e9",	--3313
		x"e8",	--3314
		x"e8",	--3315
		x"e8",	--3316
		x"e8",	--3317
		x"e9",	--3318
		x"e8",	--3319
		x"e8",	--3320
		x"e8",	--3321
		x"e8",	--3322
		x"e8",	--3323
		x"31",	--3324
		x"33",	--3325
		x"35",	--3326
		x"37",	--3327
		x"39",	--3328
		x"62",	--3329
		x"64",	--3330
		x"66",	--3331
		x"00",	--3332
		x"00",	--3333
		x"00",	--3334
		x"00",	--3335
		x"00",	--3336
		x"01",	--3337
		x"02",	--3338
		x"03",	--3339
		x"03",	--3340
		x"04",	--3341
		x"04",	--3342
		x"04",	--3343
		x"04",	--3344
		x"05",	--3345
		x"05",	--3346
		x"05",	--3347
		x"05",	--3348
		x"05",	--3349
		x"05",	--3350
		x"05",	--3351
		x"05",	--3352
		x"06",	--3353
		x"06",	--3354
		x"06",	--3355
		x"06",	--3356
		x"06",	--3357
		x"06",	--3358
		x"06",	--3359
		x"06",	--3360
		x"06",	--3361
		x"06",	--3362
		x"06",	--3363
		x"06",	--3364
		x"06",	--3365
		x"06",	--3366
		x"06",	--3367
		x"06",	--3368
		x"07",	--3369
		x"07",	--3370
		x"07",	--3371
		x"07",	--3372
		x"07",	--3373
		x"07",	--3374
		x"07",	--3375
		x"07",	--3376
		x"07",	--3377
		x"07",	--3378
		x"07",	--3379
		x"07",	--3380
		x"07",	--3381
		x"07",	--3382
		x"07",	--3383
		x"07",	--3384
		x"07",	--3385
		x"07",	--3386
		x"07",	--3387
		x"07",	--3388
		x"07",	--3389
		x"07",	--3390
		x"07",	--3391
		x"07",	--3392
		x"07",	--3393
		x"07",	--3394
		x"07",	--3395
		x"07",	--3396
		x"07",	--3397
		x"07",	--3398
		x"07",	--3399
		x"07",	--3400
		x"08",	--3401
		x"08",	--3402
		x"08",	--3403
		x"08",	--3404
		x"08",	--3405
		x"08",	--3406
		x"08",	--3407
		x"08",	--3408
		x"08",	--3409
		x"08",	--3410
		x"08",	--3411
		x"08",	--3412
		x"08",	--3413
		x"08",	--3414
		x"08",	--3415
		x"08",	--3416
		x"08",	--3417
		x"08",	--3418
		x"08",	--3419
		x"08",	--3420
		x"08",	--3421
		x"08",	--3422
		x"08",	--3423
		x"08",	--3424
		x"08",	--3425
		x"08",	--3426
		x"08",	--3427
		x"08",	--3428
		x"08",	--3429
		x"08",	--3430
		x"08",	--3431
		x"08",	--3432
		x"08",	--3433
		x"08",	--3434
		x"08",	--3435
		x"08",	--3436
		x"08",	--3437
		x"08",	--3438
		x"08",	--3439
		x"08",	--3440
		x"08",	--3441
		x"08",	--3442
		x"08",	--3443
		x"08",	--3444
		x"08",	--3445
		x"08",	--3446
		x"08",	--3447
		x"08",	--3448
		x"08",	--3449
		x"08",	--3450
		x"08",	--3451
		x"08",	--3452
		x"08",	--3453
		x"08",	--3454
		x"08",	--3455
		x"08",	--3456
		x"08",	--3457
		x"08",	--3458
		x"08",	--3459
		x"08",	--3460
		x"08",	--3461
		x"08",	--3462
		x"08",	--3463
		x"08",	--3464
		x"65",	--3465
		x"70",	--3466
		x"00",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"e9",	--4087
		x"e1",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
