library ieee;
use ieee.std_logic_1164.all;

library work;
use work.ram16_pkg.all;

package init_ram16_pkg is
	constant mcu_firmware_l : ram8_t := (
		x"55",	--0
		x"20",	--1
		x"35",	--2
		x"08",	--3
		x"82",	--4
		x"4a",	--5
		x"31",	--6
		x"00",	--7
		x"3f",	--8
		x"00",	--9
		x"0f",	--10
		x"08",	--11
		x"92",	--12
		x"4a",	--13
		x"20",	--14
		x"2f",	--15
		x"9f",	--16
		x"d0",	--17
		x"00",	--18
		x"f8",	--19
		x"3f",	--20
		x"4a",	--21
		x"0f",	--22
		x"07",	--23
		x"92",	--24
		x"4a",	--25
		x"20",	--26
		x"1f",	--27
		x"cf",	--28
		x"00",	--29
		x"f9",	--30
		x"31",	--31
		x"c2",	--32
		x"b2",	--33
		x"80",	--34
		x"20",	--35
		x"f2",	--36
		x"1a",	--37
		x"c2",	--38
		x"22",	--39
		x"3e",	--40
		x"00",	--41
		x"1f",	--42
		x"b0",	--43
		x"0c",	--44
		x"b0",	--45
		x"74",	--46
		x"c2",	--47
		x"19",	--48
		x"3e",	--49
		x"4c",	--50
		x"7f",	--51
		x"77",	--52
		x"b0",	--53
		x"76",	--54
		x"3e",	--55
		x"ec",	--56
		x"7f",	--57
		x"72",	--58
		x"b0",	--59
		x"76",	--60
		x"3e",	--61
		x"9a",	--62
		x"7f",	--63
		x"70",	--64
		x"b0",	--65
		x"76",	--66
		x"2c",	--67
		x"3d",	--68
		x"20",	--69
		x"3e",	--70
		x"80",	--71
		x"0f",	--72
		x"3f",	--73
		x"0a",	--74
		x"b0",	--75
		x"84",	--76
		x"0f",	--77
		x"3f",	--78
		x"0a",	--79
		x"b0",	--80
		x"cc",	--81
		x"2c",	--82
		x"3d",	--83
		x"20",	--84
		x"3e",	--85
		x"88",	--86
		x"0f",	--87
		x"b0",	--88
		x"84",	--89
		x"0f",	--90
		x"b0",	--91
		x"cc",	--92
		x"0e",	--93
		x"0f",	--94
		x"3f",	--95
		x"0a",	--96
		x"b0",	--97
		x"90",	--98
		x"f2",	--99
		x"80",	--100
		x"19",	--101
		x"32",	--102
		x"0b",	--103
		x"30",	--104
		x"60",	--105
		x"b0",	--106
		x"ca",	--107
		x"21",	--108
		x"0a",	--109
		x"32",	--110
		x"10",	--111
		x"1b",	--112
		x"3b",	--113
		x"09",	--114
		x"0a",	--115
		x"1f",	--116
		x"4e",	--117
		x"7e",	--118
		x"0f",	--119
		x"03",	--120
		x"0f",	--121
		x"7e",	--122
		x"fd",	--123
		x"4f",	--124
		x"02",	--125
		x"5f",	--126
		x"0b",	--127
		x"c2",	--128
		x"19",	--129
		x"b0",	--130
		x"1a",	--131
		x"0f",	--132
		x"e8",	--133
		x"b0",	--134
		x"42",	--135
		x"7f",	--136
		x"1c",	--137
		x"7f",	--138
		x"0d",	--139
		x"22",	--140
		x"30",	--141
		x"63",	--142
		x"b0",	--143
		x"ca",	--144
		x"21",	--145
		x"3f",	--146
		x"14",	--147
		x"0f",	--148
		x"0a",	--149
		x"ca",	--150
		x"00",	--151
		x"0f",	--152
		x"30",	--153
		x"66",	--154
		x"b0",	--155
		x"ca",	--156
		x"21",	--157
		x"0e",	--158
		x"3e",	--159
		x"14",	--160
		x"5f",	--161
		x"14",	--162
		x"b0",	--163
		x"a0",	--164
		x"c2",	--165
		x"0a",	--166
		x"c6",	--167
		x"3a",	--168
		x"30",	--169
		x"6c",	--170
		x"b0",	--171
		x"ca",	--172
		x"21",	--173
		x"bf",	--174
		x"3a",	--175
		x"28",	--176
		x"bc",	--177
		x"4e",	--178
		x"8e",	--179
		x"0e",	--180
		x"30",	--181
		x"70",	--182
		x"81",	--183
		x"40",	--184
		x"b0",	--185
		x"ca",	--186
		x"21",	--187
		x"3e",	--188
		x"14",	--189
		x"0e",	--190
		x"0e",	--191
		x"1f",	--192
		x"3c",	--193
		x"ce",	--194
		x"00",	--195
		x"1a",	--196
		x"a8",	--197
		x"30",	--198
		x"16",	--199
		x"82",	--200
		x"08",	--201
		x"82",	--202
		x"06",	--203
		x"30",	--204
		x"31",	--205
		x"ff",	--206
		x"20",	--207
		x"01",	--208
		x"39",	--209
		x"cf",	--210
		x"02",	--211
		x"36",	--212
		x"0d",	--213
		x"0e",	--214
		x"2e",	--215
		x"0f",	--216
		x"2f",	--217
		x"b0",	--218
		x"6a",	--219
		x"81",	--220
		x"00",	--221
		x"40",	--222
		x"0d",	--223
		x"0e",	--224
		x"0f",	--225
		x"2f",	--226
		x"b0",	--227
		x"6a",	--228
		x"81",	--229
		x"00",	--230
		x"37",	--231
		x"1e",	--232
		x"04",	--233
		x"0f",	--234
		x"b0",	--235
		x"34",	--236
		x"0c",	--237
		x"3d",	--238
		x"c8",	--239
		x"b0",	--240
		x"04",	--241
		x"0d",	--242
		x"0e",	--243
		x"1f",	--244
		x"08",	--245
		x"b0",	--246
		x"20",	--247
		x"1e",	--248
		x"02",	--249
		x"0f",	--250
		x"b0",	--251
		x"34",	--252
		x"0c",	--253
		x"3d",	--254
		x"c8",	--255
		x"b0",	--256
		x"04",	--257
		x"0d",	--258
		x"0e",	--259
		x"1f",	--260
		x"06",	--261
		x"b0",	--262
		x"20",	--263
		x"0f",	--264
		x"31",	--265
		x"30",	--266
		x"30",	--267
		x"1e",	--268
		x"81",	--269
		x"08",	--270
		x"b0",	--271
		x"ca",	--272
		x"1f",	--273
		x"08",	--274
		x"6f",	--275
		x"8f",	--276
		x"81",	--277
		x"00",	--278
		x"30",	--279
		x"2f",	--280
		x"b0",	--281
		x"ca",	--282
		x"21",	--283
		x"3f",	--284
		x"31",	--285
		x"30",	--286
		x"30",	--287
		x"40",	--288
		x"b0",	--289
		x"ca",	--290
		x"21",	--291
		x"3f",	--292
		x"e3",	--293
		x"0b",	--294
		x"31",	--295
		x"fa",	--296
		x"0b",	--297
		x"30",	--298
		x"73",	--299
		x"b0",	--300
		x"ca",	--301
		x"21",	--302
		x"fb",	--303
		x"20",	--304
		x"01",	--305
		x"2a",	--306
		x"cb",	--307
		x"02",	--308
		x"27",	--309
		x"0d",	--310
		x"0e",	--311
		x"2e",	--312
		x"0f",	--313
		x"2f",	--314
		x"b0",	--315
		x"6a",	--316
		x"81",	--317
		x"00",	--318
		x"2f",	--319
		x"0d",	--320
		x"0e",	--321
		x"0f",	--322
		x"2f",	--323
		x"b0",	--324
		x"6a",	--325
		x"81",	--326
		x"00",	--327
		x"26",	--328
		x"11",	--329
		x"04",	--330
		x"11",	--331
		x"08",	--332
		x"30",	--333
		x"c1",	--334
		x"b0",	--335
		x"ca",	--336
		x"31",	--337
		x"06",	--338
		x"1f",	--339
		x"04",	--340
		x"9f",	--341
		x"02",	--342
		x"00",	--343
		x"0f",	--344
		x"31",	--345
		x"06",	--346
		x"3b",	--347
		x"30",	--348
		x"30",	--349
		x"7b",	--350
		x"b0",	--351
		x"ca",	--352
		x"6f",	--353
		x"8f",	--354
		x"81",	--355
		x"00",	--356
		x"30",	--357
		x"8c",	--358
		x"b0",	--359
		x"ca",	--360
		x"21",	--361
		x"3f",	--362
		x"31",	--363
		x"06",	--364
		x"3b",	--365
		x"30",	--366
		x"30",	--367
		x"a1",	--368
		x"b0",	--369
		x"ca",	--370
		x"21",	--371
		x"3f",	--372
		x"e3",	--373
		x"0b",	--374
		x"21",	--375
		x"0b",	--376
		x"30",	--377
		x"cd",	--378
		x"b0",	--379
		x"ca",	--380
		x"21",	--381
		x"fb",	--382
		x"20",	--383
		x"01",	--384
		x"1b",	--385
		x"cb",	--386
		x"02",	--387
		x"18",	--388
		x"0d",	--389
		x"0e",	--390
		x"2e",	--391
		x"0f",	--392
		x"2f",	--393
		x"b0",	--394
		x"6a",	--395
		x"81",	--396
		x"00",	--397
		x"1f",	--398
		x"1f",	--399
		x"02",	--400
		x"2f",	--401
		x"0f",	--402
		x"30",	--403
		x"c1",	--404
		x"b0",	--405
		x"ca",	--406
		x"31",	--407
		x"06",	--408
		x"0f",	--409
		x"21",	--410
		x"3b",	--411
		x"30",	--412
		x"30",	--413
		x"7b",	--414
		x"b0",	--415
		x"ca",	--416
		x"6f",	--417
		x"8f",	--418
		x"81",	--419
		x"00",	--420
		x"30",	--421
		x"d4",	--422
		x"b0",	--423
		x"ca",	--424
		x"21",	--425
		x"3f",	--426
		x"21",	--427
		x"3b",	--428
		x"30",	--429
		x"30",	--430
		x"a1",	--431
		x"b0",	--432
		x"ca",	--433
		x"21",	--434
		x"3f",	--435
		x"e5",	--436
		x"0b",	--437
		x"0a",	--438
		x"09",	--439
		x"08",	--440
		x"07",	--441
		x"8f",	--442
		x"00",	--443
		x"8d",	--444
		x"00",	--445
		x"6c",	--446
		x"4c",	--447
		x"5f",	--448
		x"0b",	--449
		x"1b",	--450
		x"08",	--451
		x"0a",	--452
		x"07",	--453
		x"09",	--454
		x"18",	--455
		x"7a",	--456
		x"0a",	--457
		x"35",	--458
		x"2c",	--459
		x"0c",	--460
		x"0c",	--461
		x"0c",	--462
		x"0c",	--463
		x"8f",	--464
		x"00",	--465
		x"3c",	--466
		x"d0",	--467
		x"6a",	--468
		x"8a",	--469
		x"0c",	--470
		x"8f",	--471
		x"00",	--472
		x"17",	--473
		x"19",	--474
		x"0a",	--475
		x"08",	--476
		x"7c",	--477
		x"4c",	--478
		x"40",	--479
		x"7c",	--480
		x"78",	--481
		x"1b",	--482
		x"7c",	--483
		x"20",	--484
		x"43",	--485
		x"4a",	--486
		x"7a",	--487
		x"d0",	--488
		x"07",	--489
		x"dd",	--490
		x"7a",	--491
		x"0a",	--492
		x"46",	--493
		x"2a",	--494
		x"0a",	--495
		x"0c",	--496
		x"0c",	--497
		x"0c",	--498
		x"0c",	--499
		x"8f",	--500
		x"00",	--501
		x"3c",	--502
		x"d0",	--503
		x"68",	--504
		x"88",	--505
		x"0c",	--506
		x"8f",	--507
		x"00",	--508
		x"dc",	--509
		x"17",	--510
		x"da",	--511
		x"4a",	--512
		x"7a",	--513
		x"9f",	--514
		x"7a",	--515
		x"06",	--516
		x"0a",	--517
		x"2c",	--518
		x"0c",	--519
		x"0c",	--520
		x"0c",	--521
		x"0c",	--522
		x"8f",	--523
		x"00",	--524
		x"3c",	--525
		x"a9",	--526
		x"c4",	--527
		x"4a",	--528
		x"7a",	--529
		x"bf",	--530
		x"7a",	--531
		x"06",	--532
		x"1e",	--533
		x"2c",	--534
		x"0c",	--535
		x"0c",	--536
		x"0c",	--537
		x"0c",	--538
		x"8f",	--539
		x"00",	--540
		x"3c",	--541
		x"c9",	--542
		x"b4",	--543
		x"9d",	--544
		x"00",	--545
		x"0f",	--546
		x"37",	--547
		x"38",	--548
		x"39",	--549
		x"3a",	--550
		x"3b",	--551
		x"30",	--552
		x"9d",	--553
		x"00",	--554
		x"0f",	--555
		x"1f",	--556
		x"0f",	--557
		x"37",	--558
		x"38",	--559
		x"39",	--560
		x"3a",	--561
		x"3b",	--562
		x"30",	--563
		x"8c",	--564
		x"0c",	--565
		x"30",	--566
		x"e3",	--567
		x"b0",	--568
		x"ca",	--569
		x"21",	--570
		x"0f",	--571
		x"37",	--572
		x"38",	--573
		x"39",	--574
		x"3a",	--575
		x"3b",	--576
		x"30",	--577
		x"0b",	--578
		x"0a",	--579
		x"0b",	--580
		x"0a",	--581
		x"8f",	--582
		x"00",	--583
		x"8f",	--584
		x"02",	--585
		x"8f",	--586
		x"04",	--587
		x"0c",	--588
		x"0d",	--589
		x"3e",	--590
		x"00",	--591
		x"3f",	--592
		x"6e",	--593
		x"b0",	--594
		x"68",	--595
		x"8b",	--596
		x"02",	--597
		x"02",	--598
		x"32",	--599
		x"03",	--600
		x"82",	--601
		x"32",	--602
		x"b2",	--603
		x"18",	--604
		x"38",	--605
		x"9b",	--606
		x"3a",	--607
		x"06",	--608
		x"32",	--609
		x"0f",	--610
		x"3a",	--611
		x"3b",	--612
		x"30",	--613
		x"0b",	--614
		x"09",	--615
		x"08",	--616
		x"8f",	--617
		x"06",	--618
		x"bf",	--619
		x"00",	--620
		x"08",	--621
		x"2b",	--622
		x"1e",	--623
		x"02",	--624
		x"0f",	--625
		x"b0",	--626
		x"34",	--627
		x"0c",	--628
		x"3d",	--629
		x"00",	--630
		x"b0",	--631
		x"e0",	--632
		x"08",	--633
		x"09",	--634
		x"1e",	--635
		x"06",	--636
		x"0f",	--637
		x"b0",	--638
		x"34",	--639
		x"0c",	--640
		x"0d",	--641
		x"0e",	--642
		x"0f",	--643
		x"b0",	--644
		x"90",	--645
		x"b0",	--646
		x"70",	--647
		x"8b",	--648
		x"04",	--649
		x"9b",	--650
		x"00",	--651
		x"38",	--652
		x"39",	--653
		x"3b",	--654
		x"30",	--655
		x"0b",	--656
		x"0a",	--657
		x"09",	--658
		x"0a",	--659
		x"0b",	--660
		x"8f",	--661
		x"06",	--662
		x"8f",	--663
		x"08",	--664
		x"29",	--665
		x"1e",	--666
		x"02",	--667
		x"0f",	--668
		x"b0",	--669
		x"34",	--670
		x"0c",	--671
		x"0d",	--672
		x"0e",	--673
		x"0f",	--674
		x"b0",	--675
		x"e0",	--676
		x"0a",	--677
		x"0b",	--678
		x"1e",	--679
		x"06",	--680
		x"0f",	--681
		x"b0",	--682
		x"34",	--683
		x"0c",	--684
		x"0d",	--685
		x"0e",	--686
		x"0f",	--687
		x"b0",	--688
		x"90",	--689
		x"b0",	--690
		x"70",	--691
		x"89",	--692
		x"04",	--693
		x"39",	--694
		x"3a",	--695
		x"3b",	--696
		x"30",	--697
		x"30",	--698
		x"1c",	--699
		x"00",	--700
		x"3c",	--701
		x"40",	--702
		x"0e",	--703
		x"0d",	--704
		x"0d",	--705
		x"0d",	--706
		x"3d",	--707
		x"0a",	--708
		x"cd",	--709
		x"00",	--710
		x"8d",	--711
		x"02",	--712
		x"1c",	--713
		x"82",	--714
		x"00",	--715
		x"0f",	--716
		x"30",	--717
		x"3f",	--718
		x"30",	--719
		x"0b",	--720
		x"1b",	--721
		x"00",	--722
		x"1b",	--723
		x"0e",	--724
		x"5f",	--725
		x"0a",	--726
		x"13",	--727
		x"3d",	--728
		x"0e",	--729
		x"0c",	--730
		x"04",	--731
		x"2d",	--732
		x"cd",	--733
		x"fc",	--734
		x"0c",	--735
		x"1c",	--736
		x"0c",	--737
		x"f9",	--738
		x"30",	--739
		x"f8",	--740
		x"b0",	--741
		x"ca",	--742
		x"21",	--743
		x"3f",	--744
		x"3b",	--745
		x"30",	--746
		x"0c",	--747
		x"0c",	--748
		x"0c",	--749
		x"3c",	--750
		x"0a",	--751
		x"0f",	--752
		x"9c",	--753
		x"02",	--754
		x"3b",	--755
		x"30",	--756
		x"5e",	--757
		x"81",	--758
		x"3e",	--759
		x"fc",	--760
		x"c2",	--761
		x"19",	--762
		x"c2",	--763
		x"84",	--764
		x"0f",	--765
		x"30",	--766
		x"3f",	--767
		x"0f",	--768
		x"5f",	--769
		x"b6",	--770
		x"8f",	--771
		x"b0",	--772
		x"ea",	--773
		x"30",	--774
		x"0b",	--775
		x"0b",	--776
		x"0e",	--777
		x"0e",	--778
		x"0e",	--779
		x"0e",	--780
		x"0e",	--781
		x"0f",	--782
		x"b0",	--783
		x"fe",	--784
		x"0f",	--785
		x"b0",	--786
		x"fe",	--787
		x"3b",	--788
		x"30",	--789
		x"0b",	--790
		x"0a",	--791
		x"0a",	--792
		x"3b",	--793
		x"07",	--794
		x"0e",	--795
		x"4d",	--796
		x"7d",	--797
		x"0f",	--798
		x"03",	--799
		x"0e",	--800
		x"7d",	--801
		x"fd",	--802
		x"1e",	--803
		x"0a",	--804
		x"3f",	--805
		x"31",	--806
		x"b0",	--807
		x"ea",	--808
		x"3b",	--809
		x"3b",	--810
		x"ef",	--811
		x"3a",	--812
		x"3b",	--813
		x"30",	--814
		x"3f",	--815
		x"30",	--816
		x"f5",	--817
		x"0b",	--818
		x"0b",	--819
		x"0e",	--820
		x"8e",	--821
		x"8e",	--822
		x"0f",	--823
		x"b0",	--824
		x"0e",	--825
		x"0f",	--826
		x"b0",	--827
		x"0e",	--828
		x"3b",	--829
		x"30",	--830
		x"0b",	--831
		x"0a",	--832
		x"0a",	--833
		x"0b",	--834
		x"0d",	--835
		x"8d",	--836
		x"8d",	--837
		x"0f",	--838
		x"b0",	--839
		x"0e",	--840
		x"0f",	--841
		x"b0",	--842
		x"0e",	--843
		x"0c",	--844
		x"0d",	--845
		x"8d",	--846
		x"8c",	--847
		x"4d",	--848
		x"0d",	--849
		x"0f",	--850
		x"b0",	--851
		x"0e",	--852
		x"0f",	--853
		x"b0",	--854
		x"0e",	--855
		x"3a",	--856
		x"3b",	--857
		x"30",	--858
		x"0b",	--859
		x"0a",	--860
		x"09",	--861
		x"0a",	--862
		x"0e",	--863
		x"19",	--864
		x"09",	--865
		x"39",	--866
		x"0b",	--867
		x"0d",	--868
		x"0d",	--869
		x"6f",	--870
		x"8f",	--871
		x"b0",	--872
		x"0e",	--873
		x"0b",	--874
		x"0e",	--875
		x"1b",	--876
		x"3b",	--877
		x"07",	--878
		x"05",	--879
		x"3f",	--880
		x"20",	--881
		x"b0",	--882
		x"ea",	--883
		x"ef",	--884
		x"3f",	--885
		x"3a",	--886
		x"b0",	--887
		x"ea",	--888
		x"ea",	--889
		x"39",	--890
		x"3a",	--891
		x"3b",	--892
		x"30",	--893
		x"0b",	--894
		x"0a",	--895
		x"09",	--896
		x"0a",	--897
		x"0e",	--898
		x"17",	--899
		x"09",	--900
		x"39",	--901
		x"0b",	--902
		x"6f",	--903
		x"8f",	--904
		x"b0",	--905
		x"fe",	--906
		x"0b",	--907
		x"0e",	--908
		x"1b",	--909
		x"3b",	--910
		x"07",	--911
		x"f6",	--912
		x"3f",	--913
		x"20",	--914
		x"b0",	--915
		x"ea",	--916
		x"6f",	--917
		x"8f",	--918
		x"b0",	--919
		x"fe",	--920
		x"0b",	--921
		x"f2",	--922
		x"39",	--923
		x"3a",	--924
		x"3b",	--925
		x"30",	--926
		x"0b",	--927
		x"0a",	--928
		x"09",	--929
		x"31",	--930
		x"ec",	--931
		x"0b",	--932
		x"0f",	--933
		x"34",	--934
		x"3b",	--935
		x"0a",	--936
		x"38",	--937
		x"09",	--938
		x"0a",	--939
		x"0a",	--940
		x"3e",	--941
		x"0a",	--942
		x"0f",	--943
		x"b0",	--944
		x"60",	--945
		x"7f",	--946
		x"30",	--947
		x"ca",	--948
		x"00",	--949
		x"19",	--950
		x"3e",	--951
		x"0a",	--952
		x"0f",	--953
		x"b0",	--954
		x"2e",	--955
		x"0b",	--956
		x"3f",	--957
		x"0a",	--958
		x"eb",	--959
		x"0a",	--960
		x"1a",	--961
		x"09",	--962
		x"3e",	--963
		x"0a",	--964
		x"0f",	--965
		x"b0",	--966
		x"60",	--967
		x"7f",	--968
		x"30",	--969
		x"c9",	--970
		x"00",	--971
		x"3a",	--972
		x"0f",	--973
		x"0f",	--974
		x"6f",	--975
		x"8f",	--976
		x"b0",	--977
		x"ea",	--978
		x"0a",	--979
		x"f7",	--980
		x"31",	--981
		x"14",	--982
		x"39",	--983
		x"3a",	--984
		x"3b",	--985
		x"30",	--986
		x"3f",	--987
		x"2d",	--988
		x"b0",	--989
		x"ea",	--990
		x"3b",	--991
		x"1b",	--992
		x"c5",	--993
		x"1a",	--994
		x"09",	--995
		x"dd",	--996
		x"0b",	--997
		x"0a",	--998
		x"09",	--999
		x"0b",	--1000
		x"3b",	--1001
		x"39",	--1002
		x"6f",	--1003
		x"4f",	--1004
		x"0b",	--1005
		x"1a",	--1006
		x"8f",	--1007
		x"b0",	--1008
		x"ea",	--1009
		x"0a",	--1010
		x"09",	--1011
		x"19",	--1012
		x"5f",	--1013
		x"01",	--1014
		x"4f",	--1015
		x"10",	--1016
		x"7f",	--1017
		x"25",	--1018
		x"f3",	--1019
		x"0a",	--1020
		x"1a",	--1021
		x"5f",	--1022
		x"01",	--1023
		x"7f",	--1024
		x"db",	--1025
		x"7f",	--1026
		x"54",	--1027
		x"ee",	--1028
		x"4f",	--1029
		x"0f",	--1030
		x"10",	--1031
		x"0e",	--1032
		x"39",	--1033
		x"3a",	--1034
		x"3b",	--1035
		x"30",	--1036
		x"09",	--1037
		x"29",	--1038
		x"1e",	--1039
		x"02",	--1040
		x"2f",	--1041
		x"b0",	--1042
		x"b6",	--1043
		x"0b",	--1044
		x"dd",	--1045
		x"09",	--1046
		x"29",	--1047
		x"2f",	--1048
		x"b0",	--1049
		x"64",	--1050
		x"0b",	--1051
		x"d6",	--1052
		x"0f",	--1053
		x"2b",	--1054
		x"29",	--1055
		x"6f",	--1056
		x"4f",	--1057
		x"d0",	--1058
		x"19",	--1059
		x"8f",	--1060
		x"b0",	--1061
		x"ea",	--1062
		x"7f",	--1063
		x"4f",	--1064
		x"fa",	--1065
		x"c8",	--1066
		x"09",	--1067
		x"29",	--1068
		x"1e",	--1069
		x"02",	--1070
		x"2f",	--1071
		x"b0",	--1072
		x"fc",	--1073
		x"0b",	--1074
		x"bf",	--1075
		x"09",	--1076
		x"29",	--1077
		x"2e",	--1078
		x"0f",	--1079
		x"8f",	--1080
		x"8f",	--1081
		x"8f",	--1082
		x"8f",	--1083
		x"b0",	--1084
		x"7e",	--1085
		x"0b",	--1086
		x"b3",	--1087
		x"09",	--1088
		x"29",	--1089
		x"2f",	--1090
		x"b0",	--1091
		x"3e",	--1092
		x"0b",	--1093
		x"ac",	--1094
		x"09",	--1095
		x"29",	--1096
		x"2f",	--1097
		x"b0",	--1098
		x"ea",	--1099
		x"0b",	--1100
		x"a5",	--1101
		x"09",	--1102
		x"29",	--1103
		x"2f",	--1104
		x"b0",	--1105
		x"0e",	--1106
		x"0b",	--1107
		x"9e",	--1108
		x"09",	--1109
		x"29",	--1110
		x"2f",	--1111
		x"b0",	--1112
		x"2c",	--1113
		x"0b",	--1114
		x"97",	--1115
		x"3f",	--1116
		x"25",	--1117
		x"b0",	--1118
		x"ea",	--1119
		x"92",	--1120
		x"0f",	--1121
		x"0e",	--1122
		x"1f",	--1123
		x"02",	--1124
		x"df",	--1125
		x"85",	--1126
		x"0a",	--1127
		x"1f",	--1128
		x"02",	--1129
		x"3f",	--1130
		x"3f",	--1131
		x"16",	--1132
		x"92",	--1133
		x"02",	--1134
		x"1e",	--1135
		x"02",	--1136
		x"1f",	--1137
		x"04",	--1138
		x"0e",	--1139
		x"02",	--1140
		x"92",	--1141
		x"04",	--1142
		x"f2",	--1143
		x"10",	--1144
		x"81",	--1145
		x"b1",	--1146
		x"10",	--1147
		x"04",	--1148
		x"3e",	--1149
		x"3f",	--1150
		x"b1",	--1151
		x"f0",	--1152
		x"00",	--1153
		x"00",	--1154
		x"82",	--1155
		x"02",	--1156
		x"e9",	--1157
		x"b2",	--1158
		x"cf",	--1159
		x"82",	--1160
		x"f2",	--1161
		x"11",	--1162
		x"80",	--1163
		x"30",	--1164
		x"1e",	--1165
		x"02",	--1166
		x"1f",	--1167
		x"04",	--1168
		x"0e",	--1169
		x"05",	--1170
		x"1f",	--1171
		x"02",	--1172
		x"1f",	--1173
		x"04",	--1174
		x"30",	--1175
		x"1d",	--1176
		x"02",	--1177
		x"1e",	--1178
		x"04",	--1179
		x"3f",	--1180
		x"40",	--1181
		x"0f",	--1182
		x"0f",	--1183
		x"30",	--1184
		x"1f",	--1185
		x"04",	--1186
		x"5f",	--1187
		x"0a",	--1188
		x"1d",	--1189
		x"04",	--1190
		x"1e",	--1191
		x"02",	--1192
		x"0d",	--1193
		x"0b",	--1194
		x"1e",	--1195
		x"04",	--1196
		x"3e",	--1197
		x"3f",	--1198
		x"03",	--1199
		x"82",	--1200
		x"04",	--1201
		x"30",	--1202
		x"92",	--1203
		x"04",	--1204
		x"30",	--1205
		x"4f",	--1206
		x"30",	--1207
		x"0b",	--1208
		x"0a",	--1209
		x"0a",	--1210
		x"0b",	--1211
		x"0c",	--1212
		x"3d",	--1213
		x"00",	--1214
		x"b0",	--1215
		x"54",	--1216
		x"0f",	--1217
		x"07",	--1218
		x"0e",	--1219
		x"0f",	--1220
		x"b0",	--1221
		x"a4",	--1222
		x"3a",	--1223
		x"3b",	--1224
		x"30",	--1225
		x"0c",	--1226
		x"3d",	--1227
		x"00",	--1228
		x"0e",	--1229
		x"0f",	--1230
		x"b0",	--1231
		x"90",	--1232
		x"b0",	--1233
		x"a4",	--1234
		x"0e",	--1235
		x"3f",	--1236
		x"00",	--1237
		x"3a",	--1238
		x"3b",	--1239
		x"30",	--1240
		x"0b",	--1241
		x"0a",	--1242
		x"09",	--1243
		x"08",	--1244
		x"07",	--1245
		x"06",	--1246
		x"05",	--1247
		x"04",	--1248
		x"31",	--1249
		x"fa",	--1250
		x"08",	--1251
		x"6b",	--1252
		x"6b",	--1253
		x"67",	--1254
		x"6c",	--1255
		x"6c",	--1256
		x"e9",	--1257
		x"6b",	--1258
		x"02",	--1259
		x"30",	--1260
		x"32",	--1261
		x"6c",	--1262
		x"e3",	--1263
		x"6c",	--1264
		x"bb",	--1265
		x"6b",	--1266
		x"df",	--1267
		x"91",	--1268
		x"02",	--1269
		x"00",	--1270
		x"1b",	--1271
		x"02",	--1272
		x"14",	--1273
		x"04",	--1274
		x"15",	--1275
		x"06",	--1276
		x"16",	--1277
		x"04",	--1278
		x"17",	--1279
		x"06",	--1280
		x"2c",	--1281
		x"0c",	--1282
		x"09",	--1283
		x"0c",	--1284
		x"bf",	--1285
		x"39",	--1286
		x"20",	--1287
		x"50",	--1288
		x"1c",	--1289
		x"d7",	--1290
		x"81",	--1291
		x"02",	--1292
		x"81",	--1293
		x"04",	--1294
		x"4c",	--1295
		x"7c",	--1296
		x"1f",	--1297
		x"0b",	--1298
		x"0a",	--1299
		x"0b",	--1300
		x"12",	--1301
		x"0b",	--1302
		x"0a",	--1303
		x"7c",	--1304
		x"fb",	--1305
		x"81",	--1306
		x"02",	--1307
		x"81",	--1308
		x"04",	--1309
		x"1c",	--1310
		x"0d",	--1311
		x"79",	--1312
		x"1f",	--1313
		x"04",	--1314
		x"0c",	--1315
		x"0d",	--1316
		x"79",	--1317
		x"fc",	--1318
		x"3c",	--1319
		x"3d",	--1320
		x"0c",	--1321
		x"0d",	--1322
		x"1a",	--1323
		x"0b",	--1324
		x"0c",	--1325
		x"02",	--1326
		x"0d",	--1327
		x"e5",	--1328
		x"16",	--1329
		x"02",	--1330
		x"17",	--1331
		x"04",	--1332
		x"06",	--1333
		x"07",	--1334
		x"5f",	--1335
		x"01",	--1336
		x"5f",	--1337
		x"01",	--1338
		x"28",	--1339
		x"c8",	--1340
		x"01",	--1341
		x"a8",	--1342
		x"02",	--1343
		x"0e",	--1344
		x"0f",	--1345
		x"0e",	--1346
		x"0f",	--1347
		x"88",	--1348
		x"04",	--1349
		x"88",	--1350
		x"06",	--1351
		x"f8",	--1352
		x"03",	--1353
		x"00",	--1354
		x"0f",	--1355
		x"4d",	--1356
		x"0f",	--1357
		x"31",	--1358
		x"06",	--1359
		x"34",	--1360
		x"35",	--1361
		x"36",	--1362
		x"37",	--1363
		x"38",	--1364
		x"39",	--1365
		x"3a",	--1366
		x"3b",	--1367
		x"30",	--1368
		x"2b",	--1369
		x"67",	--1370
		x"81",	--1371
		x"00",	--1372
		x"04",	--1373
		x"05",	--1374
		x"5f",	--1375
		x"01",	--1376
		x"5f",	--1377
		x"01",	--1378
		x"d8",	--1379
		x"4f",	--1380
		x"68",	--1381
		x"0e",	--1382
		x"0f",	--1383
		x"0e",	--1384
		x"0f",	--1385
		x"0f",	--1386
		x"69",	--1387
		x"c8",	--1388
		x"01",	--1389
		x"a8",	--1390
		x"02",	--1391
		x"88",	--1392
		x"04",	--1393
		x"88",	--1394
		x"06",	--1395
		x"0c",	--1396
		x"0d",	--1397
		x"3c",	--1398
		x"3d",	--1399
		x"3d",	--1400
		x"ff",	--1401
		x"05",	--1402
		x"3d",	--1403
		x"00",	--1404
		x"17",	--1405
		x"3c",	--1406
		x"15",	--1407
		x"1b",	--1408
		x"02",	--1409
		x"3b",	--1410
		x"0e",	--1411
		x"0f",	--1412
		x"0a",	--1413
		x"3b",	--1414
		x"0c",	--1415
		x"0d",	--1416
		x"3c",	--1417
		x"3d",	--1418
		x"3d",	--1419
		x"ff",	--1420
		x"f5",	--1421
		x"3c",	--1422
		x"88",	--1423
		x"04",	--1424
		x"88",	--1425
		x"06",	--1426
		x"88",	--1427
		x"02",	--1428
		x"f8",	--1429
		x"03",	--1430
		x"00",	--1431
		x"0f",	--1432
		x"b3",	--1433
		x"0c",	--1434
		x"0d",	--1435
		x"1c",	--1436
		x"0d",	--1437
		x"12",	--1438
		x"0f",	--1439
		x"0e",	--1440
		x"0a",	--1441
		x"0b",	--1442
		x"0a",	--1443
		x"0b",	--1444
		x"88",	--1445
		x"04",	--1446
		x"88",	--1447
		x"06",	--1448
		x"98",	--1449
		x"02",	--1450
		x"0f",	--1451
		x"a1",	--1452
		x"6b",	--1453
		x"9f",	--1454
		x"ad",	--1455
		x"00",	--1456
		x"9d",	--1457
		x"02",	--1458
		x"02",	--1459
		x"9d",	--1460
		x"04",	--1461
		x"04",	--1462
		x"9d",	--1463
		x"06",	--1464
		x"06",	--1465
		x"5e",	--1466
		x"01",	--1467
		x"5e",	--1468
		x"01",	--1469
		x"cd",	--1470
		x"01",	--1471
		x"0f",	--1472
		x"8c",	--1473
		x"06",	--1474
		x"07",	--1475
		x"9a",	--1476
		x"39",	--1477
		x"19",	--1478
		x"39",	--1479
		x"20",	--1480
		x"8f",	--1481
		x"3e",	--1482
		x"3c",	--1483
		x"b6",	--1484
		x"c1",	--1485
		x"0e",	--1486
		x"0f",	--1487
		x"0e",	--1488
		x"0f",	--1489
		x"97",	--1490
		x"0f",	--1491
		x"79",	--1492
		x"d8",	--1493
		x"01",	--1494
		x"a8",	--1495
		x"02",	--1496
		x"3e",	--1497
		x"3f",	--1498
		x"1e",	--1499
		x"0f",	--1500
		x"88",	--1501
		x"04",	--1502
		x"88",	--1503
		x"06",	--1504
		x"92",	--1505
		x"0c",	--1506
		x"7b",	--1507
		x"81",	--1508
		x"00",	--1509
		x"81",	--1510
		x"02",	--1511
		x"81",	--1512
		x"04",	--1513
		x"4d",	--1514
		x"7d",	--1515
		x"1f",	--1516
		x"0c",	--1517
		x"4b",	--1518
		x"0c",	--1519
		x"0d",	--1520
		x"12",	--1521
		x"0d",	--1522
		x"0c",	--1523
		x"7b",	--1524
		x"fb",	--1525
		x"81",	--1526
		x"02",	--1527
		x"81",	--1528
		x"04",	--1529
		x"1c",	--1530
		x"0d",	--1531
		x"79",	--1532
		x"1f",	--1533
		x"04",	--1534
		x"0c",	--1535
		x"0d",	--1536
		x"79",	--1537
		x"fc",	--1538
		x"3c",	--1539
		x"3d",	--1540
		x"0c",	--1541
		x"0d",	--1542
		x"1a",	--1543
		x"0b",	--1544
		x"0c",	--1545
		x"04",	--1546
		x"0d",	--1547
		x"02",	--1548
		x"0a",	--1549
		x"0b",	--1550
		x"14",	--1551
		x"02",	--1552
		x"15",	--1553
		x"04",	--1554
		x"04",	--1555
		x"05",	--1556
		x"49",	--1557
		x"0a",	--1558
		x"0b",	--1559
		x"18",	--1560
		x"6c",	--1561
		x"33",	--1562
		x"df",	--1563
		x"01",	--1564
		x"01",	--1565
		x"2f",	--1566
		x"3f",	--1567
		x"c8",	--1568
		x"2c",	--1569
		x"31",	--1570
		x"e0",	--1571
		x"81",	--1572
		x"04",	--1573
		x"81",	--1574
		x"06",	--1575
		x"81",	--1576
		x"00",	--1577
		x"81",	--1578
		x"02",	--1579
		x"0e",	--1580
		x"3e",	--1581
		x"18",	--1582
		x"0f",	--1583
		x"2f",	--1584
		x"b0",	--1585
		x"66",	--1586
		x"0e",	--1587
		x"3e",	--1588
		x"10",	--1589
		x"0f",	--1590
		x"b0",	--1591
		x"66",	--1592
		x"0d",	--1593
		x"3d",	--1594
		x"0e",	--1595
		x"3e",	--1596
		x"10",	--1597
		x"0f",	--1598
		x"3f",	--1599
		x"18",	--1600
		x"b0",	--1601
		x"b2",	--1602
		x"b0",	--1603
		x"88",	--1604
		x"31",	--1605
		x"20",	--1606
		x"30",	--1607
		x"31",	--1608
		x"e0",	--1609
		x"81",	--1610
		x"04",	--1611
		x"81",	--1612
		x"06",	--1613
		x"81",	--1614
		x"00",	--1615
		x"81",	--1616
		x"02",	--1617
		x"0e",	--1618
		x"3e",	--1619
		x"18",	--1620
		x"0f",	--1621
		x"2f",	--1622
		x"b0",	--1623
		x"66",	--1624
		x"0e",	--1625
		x"3e",	--1626
		x"10",	--1627
		x"0f",	--1628
		x"b0",	--1629
		x"66",	--1630
		x"d1",	--1631
		x"11",	--1632
		x"0d",	--1633
		x"3d",	--1634
		x"0e",	--1635
		x"3e",	--1636
		x"10",	--1637
		x"0f",	--1638
		x"3f",	--1639
		x"18",	--1640
		x"b0",	--1641
		x"b2",	--1642
		x"b0",	--1643
		x"88",	--1644
		x"31",	--1645
		x"20",	--1646
		x"30",	--1647
		x"0b",	--1648
		x"0a",	--1649
		x"09",	--1650
		x"08",	--1651
		x"07",	--1652
		x"06",	--1653
		x"05",	--1654
		x"04",	--1655
		x"31",	--1656
		x"dc",	--1657
		x"81",	--1658
		x"04",	--1659
		x"81",	--1660
		x"06",	--1661
		x"81",	--1662
		x"00",	--1663
		x"81",	--1664
		x"02",	--1665
		x"0e",	--1666
		x"3e",	--1667
		x"18",	--1668
		x"0f",	--1669
		x"2f",	--1670
		x"b0",	--1671
		x"66",	--1672
		x"0e",	--1673
		x"3e",	--1674
		x"10",	--1675
		x"0f",	--1676
		x"b0",	--1677
		x"66",	--1678
		x"5f",	--1679
		x"18",	--1680
		x"6f",	--1681
		x"b6",	--1682
		x"5e",	--1683
		x"10",	--1684
		x"6e",	--1685
		x"d9",	--1686
		x"6f",	--1687
		x"ae",	--1688
		x"6e",	--1689
		x"e2",	--1690
		x"6f",	--1691
		x"ac",	--1692
		x"6e",	--1693
		x"d1",	--1694
		x"14",	--1695
		x"1c",	--1696
		x"15",	--1697
		x"1e",	--1698
		x"18",	--1699
		x"14",	--1700
		x"19",	--1701
		x"16",	--1702
		x"3c",	--1703
		x"20",	--1704
		x"0e",	--1705
		x"0f",	--1706
		x"06",	--1707
		x"07",	--1708
		x"81",	--1709
		x"20",	--1710
		x"81",	--1711
		x"22",	--1712
		x"0a",	--1713
		x"0b",	--1714
		x"81",	--1715
		x"20",	--1716
		x"08",	--1717
		x"08",	--1718
		x"09",	--1719
		x"12",	--1720
		x"05",	--1721
		x"04",	--1722
		x"b1",	--1723
		x"20",	--1724
		x"19",	--1725
		x"14",	--1726
		x"0d",	--1727
		x"0a",	--1728
		x"0b",	--1729
		x"0e",	--1730
		x"0f",	--1731
		x"1c",	--1732
		x"0d",	--1733
		x"0b",	--1734
		x"03",	--1735
		x"0b",	--1736
		x"0c",	--1737
		x"0d",	--1738
		x"0e",	--1739
		x"0f",	--1740
		x"06",	--1741
		x"07",	--1742
		x"09",	--1743
		x"e5",	--1744
		x"16",	--1745
		x"07",	--1746
		x"e2",	--1747
		x"0a",	--1748
		x"f5",	--1749
		x"f2",	--1750
		x"81",	--1751
		x"20",	--1752
		x"81",	--1753
		x"22",	--1754
		x"0c",	--1755
		x"1a",	--1756
		x"1a",	--1757
		x"1a",	--1758
		x"12",	--1759
		x"06",	--1760
		x"26",	--1761
		x"81",	--1762
		x"0a",	--1763
		x"5d",	--1764
		x"d1",	--1765
		x"11",	--1766
		x"19",	--1767
		x"83",	--1768
		x"c1",	--1769
		x"09",	--1770
		x"0c",	--1771
		x"3c",	--1772
		x"3f",	--1773
		x"00",	--1774
		x"18",	--1775
		x"1d",	--1776
		x"0a",	--1777
		x"3d",	--1778
		x"1a",	--1779
		x"20",	--1780
		x"1b",	--1781
		x"22",	--1782
		x"0c",	--1783
		x"0e",	--1784
		x"0f",	--1785
		x"0b",	--1786
		x"2a",	--1787
		x"0a",	--1788
		x"0b",	--1789
		x"3d",	--1790
		x"3f",	--1791
		x"00",	--1792
		x"f5",	--1793
		x"81",	--1794
		x"20",	--1795
		x"81",	--1796
		x"22",	--1797
		x"81",	--1798
		x"0a",	--1799
		x"0c",	--1800
		x"0d",	--1801
		x"3c",	--1802
		x"7f",	--1803
		x"0d",	--1804
		x"3c",	--1805
		x"40",	--1806
		x"44",	--1807
		x"81",	--1808
		x"0c",	--1809
		x"81",	--1810
		x"0e",	--1811
		x"f1",	--1812
		x"03",	--1813
		x"08",	--1814
		x"0f",	--1815
		x"3f",	--1816
		x"b0",	--1817
		x"88",	--1818
		x"31",	--1819
		x"24",	--1820
		x"34",	--1821
		x"35",	--1822
		x"36",	--1823
		x"37",	--1824
		x"38",	--1825
		x"39",	--1826
		x"3a",	--1827
		x"3b",	--1828
		x"30",	--1829
		x"1e",	--1830
		x"0f",	--1831
		x"d3",	--1832
		x"3a",	--1833
		x"03",	--1834
		x"08",	--1835
		x"1e",	--1836
		x"10",	--1837
		x"1c",	--1838
		x"20",	--1839
		x"1d",	--1840
		x"22",	--1841
		x"12",	--1842
		x"0d",	--1843
		x"0c",	--1844
		x"06",	--1845
		x"07",	--1846
		x"06",	--1847
		x"37",	--1848
		x"00",	--1849
		x"81",	--1850
		x"20",	--1851
		x"81",	--1852
		x"22",	--1853
		x"12",	--1854
		x"0f",	--1855
		x"0e",	--1856
		x"1a",	--1857
		x"0f",	--1858
		x"e7",	--1859
		x"81",	--1860
		x"0a",	--1861
		x"a6",	--1862
		x"6e",	--1863
		x"36",	--1864
		x"5f",	--1865
		x"d1",	--1866
		x"11",	--1867
		x"19",	--1868
		x"20",	--1869
		x"c1",	--1870
		x"19",	--1871
		x"0f",	--1872
		x"3f",	--1873
		x"18",	--1874
		x"c5",	--1875
		x"0d",	--1876
		x"ba",	--1877
		x"0c",	--1878
		x"0d",	--1879
		x"3c",	--1880
		x"80",	--1881
		x"0d",	--1882
		x"0c",	--1883
		x"b3",	--1884
		x"0d",	--1885
		x"b1",	--1886
		x"81",	--1887
		x"20",	--1888
		x"03",	--1889
		x"81",	--1890
		x"22",	--1891
		x"ab",	--1892
		x"3e",	--1893
		x"40",	--1894
		x"0f",	--1895
		x"3e",	--1896
		x"80",	--1897
		x"3f",	--1898
		x"a4",	--1899
		x"4d",	--1900
		x"7b",	--1901
		x"4f",	--1902
		x"de",	--1903
		x"5f",	--1904
		x"d1",	--1905
		x"11",	--1906
		x"19",	--1907
		x"06",	--1908
		x"c1",	--1909
		x"11",	--1910
		x"0f",	--1911
		x"3f",	--1912
		x"10",	--1913
		x"9e",	--1914
		x"4f",	--1915
		x"f8",	--1916
		x"6f",	--1917
		x"f1",	--1918
		x"3f",	--1919
		x"c8",	--1920
		x"97",	--1921
		x"0b",	--1922
		x"0a",	--1923
		x"09",	--1924
		x"08",	--1925
		x"07",	--1926
		x"31",	--1927
		x"e8",	--1928
		x"81",	--1929
		x"04",	--1930
		x"81",	--1931
		x"06",	--1932
		x"81",	--1933
		x"00",	--1934
		x"81",	--1935
		x"02",	--1936
		x"0e",	--1937
		x"3e",	--1938
		x"10",	--1939
		x"0f",	--1940
		x"2f",	--1941
		x"b0",	--1942
		x"66",	--1943
		x"0e",	--1944
		x"3e",	--1945
		x"0f",	--1946
		x"b0",	--1947
		x"66",	--1948
		x"5f",	--1949
		x"10",	--1950
		x"6f",	--1951
		x"5d",	--1952
		x"5e",	--1953
		x"08",	--1954
		x"6e",	--1955
		x"82",	--1956
		x"d1",	--1957
		x"09",	--1958
		x"11",	--1959
		x"6f",	--1960
		x"58",	--1961
		x"6f",	--1962
		x"56",	--1963
		x"6e",	--1964
		x"6f",	--1965
		x"6e",	--1966
		x"4c",	--1967
		x"1d",	--1968
		x"12",	--1969
		x"1d",	--1970
		x"0a",	--1971
		x"81",	--1972
		x"12",	--1973
		x"1e",	--1974
		x"14",	--1975
		x"1f",	--1976
		x"16",	--1977
		x"18",	--1978
		x"0c",	--1979
		x"19",	--1980
		x"0e",	--1981
		x"0f",	--1982
		x"1e",	--1983
		x"0e",	--1984
		x"0f",	--1985
		x"3d",	--1986
		x"81",	--1987
		x"12",	--1988
		x"37",	--1989
		x"1f",	--1990
		x"0c",	--1991
		x"3d",	--1992
		x"00",	--1993
		x"0a",	--1994
		x"0b",	--1995
		x"0b",	--1996
		x"0a",	--1997
		x"0b",	--1998
		x"0e",	--1999
		x"0f",	--2000
		x"12",	--2001
		x"0d",	--2002
		x"0c",	--2003
		x"0e",	--2004
		x"0f",	--2005
		x"37",	--2006
		x"0b",	--2007
		x"0f",	--2008
		x"f7",	--2009
		x"f2",	--2010
		x"0e",	--2011
		x"f4",	--2012
		x"ef",	--2013
		x"09",	--2014
		x"e5",	--2015
		x"0e",	--2016
		x"e3",	--2017
		x"dd",	--2018
		x"0c",	--2019
		x"0d",	--2020
		x"3c",	--2021
		x"7f",	--2022
		x"0d",	--2023
		x"3c",	--2024
		x"40",	--2025
		x"1c",	--2026
		x"81",	--2027
		x"14",	--2028
		x"81",	--2029
		x"16",	--2030
		x"0f",	--2031
		x"3f",	--2032
		x"10",	--2033
		x"b0",	--2034
		x"88",	--2035
		x"31",	--2036
		x"18",	--2037
		x"37",	--2038
		x"38",	--2039
		x"39",	--2040
		x"3a",	--2041
		x"3b",	--2042
		x"30",	--2043
		x"e1",	--2044
		x"10",	--2045
		x"0f",	--2046
		x"3f",	--2047
		x"10",	--2048
		x"f0",	--2049
		x"4f",	--2050
		x"fa",	--2051
		x"3f",	--2052
		x"c8",	--2053
		x"eb",	--2054
		x"0d",	--2055
		x"e2",	--2056
		x"0c",	--2057
		x"0d",	--2058
		x"3c",	--2059
		x"80",	--2060
		x"0d",	--2061
		x"0c",	--2062
		x"db",	--2063
		x"0d",	--2064
		x"d9",	--2065
		x"0e",	--2066
		x"02",	--2067
		x"0f",	--2068
		x"d5",	--2069
		x"3a",	--2070
		x"40",	--2071
		x"0b",	--2072
		x"3a",	--2073
		x"80",	--2074
		x"3b",	--2075
		x"ce",	--2076
		x"81",	--2077
		x"14",	--2078
		x"81",	--2079
		x"16",	--2080
		x"81",	--2081
		x"12",	--2082
		x"0f",	--2083
		x"3f",	--2084
		x"10",	--2085
		x"cb",	--2086
		x"0f",	--2087
		x"3f",	--2088
		x"c8",	--2089
		x"31",	--2090
		x"e8",	--2091
		x"81",	--2092
		x"04",	--2093
		x"81",	--2094
		x"06",	--2095
		x"81",	--2096
		x"00",	--2097
		x"81",	--2098
		x"02",	--2099
		x"0e",	--2100
		x"3e",	--2101
		x"10",	--2102
		x"0f",	--2103
		x"2f",	--2104
		x"b0",	--2105
		x"66",	--2106
		x"0e",	--2107
		x"3e",	--2108
		x"0f",	--2109
		x"b0",	--2110
		x"66",	--2111
		x"e1",	--2112
		x"10",	--2113
		x"0d",	--2114
		x"e1",	--2115
		x"08",	--2116
		x"0a",	--2117
		x"0e",	--2118
		x"3e",	--2119
		x"0f",	--2120
		x"3f",	--2121
		x"10",	--2122
		x"b0",	--2123
		x"8a",	--2124
		x"31",	--2125
		x"18",	--2126
		x"30",	--2127
		x"3f",	--2128
		x"fb",	--2129
		x"31",	--2130
		x"f4",	--2131
		x"81",	--2132
		x"00",	--2133
		x"81",	--2134
		x"02",	--2135
		x"0e",	--2136
		x"2e",	--2137
		x"0f",	--2138
		x"b0",	--2139
		x"66",	--2140
		x"5f",	--2141
		x"04",	--2142
		x"6f",	--2143
		x"28",	--2144
		x"27",	--2145
		x"6f",	--2146
		x"07",	--2147
		x"1d",	--2148
		x"06",	--2149
		x"0d",	--2150
		x"21",	--2151
		x"3d",	--2152
		x"1f",	--2153
		x"09",	--2154
		x"c1",	--2155
		x"05",	--2156
		x"26",	--2157
		x"3e",	--2158
		x"3f",	--2159
		x"ff",	--2160
		x"31",	--2161
		x"0c",	--2162
		x"30",	--2163
		x"1e",	--2164
		x"08",	--2165
		x"1f",	--2166
		x"0a",	--2167
		x"3c",	--2168
		x"1e",	--2169
		x"4c",	--2170
		x"4d",	--2171
		x"7d",	--2172
		x"1f",	--2173
		x"0f",	--2174
		x"c1",	--2175
		x"05",	--2176
		x"ef",	--2177
		x"3e",	--2178
		x"3f",	--2179
		x"1e",	--2180
		x"0f",	--2181
		x"31",	--2182
		x"0c",	--2183
		x"30",	--2184
		x"0e",	--2185
		x"0f",	--2186
		x"31",	--2187
		x"0c",	--2188
		x"30",	--2189
		x"12",	--2190
		x"0f",	--2191
		x"0e",	--2192
		x"7d",	--2193
		x"fb",	--2194
		x"eb",	--2195
		x"0e",	--2196
		x"3f",	--2197
		x"00",	--2198
		x"31",	--2199
		x"0c",	--2200
		x"30",	--2201
		x"0b",	--2202
		x"0a",	--2203
		x"09",	--2204
		x"08",	--2205
		x"31",	--2206
		x"0a",	--2207
		x"0b",	--2208
		x"c1",	--2209
		x"01",	--2210
		x"0e",	--2211
		x"0d",	--2212
		x"0b",	--2213
		x"0b",	--2214
		x"e1",	--2215
		x"00",	--2216
		x"0f",	--2217
		x"b0",	--2218
		x"88",	--2219
		x"31",	--2220
		x"38",	--2221
		x"39",	--2222
		x"3a",	--2223
		x"3b",	--2224
		x"30",	--2225
		x"f1",	--2226
		x"03",	--2227
		x"00",	--2228
		x"b1",	--2229
		x"1e",	--2230
		x"02",	--2231
		x"81",	--2232
		x"04",	--2233
		x"81",	--2234
		x"06",	--2235
		x"0e",	--2236
		x"0f",	--2237
		x"b0",	--2238
		x"16",	--2239
		x"3f",	--2240
		x"0f",	--2241
		x"18",	--2242
		x"e5",	--2243
		x"81",	--2244
		x"04",	--2245
		x"81",	--2246
		x"06",	--2247
		x"4e",	--2248
		x"7e",	--2249
		x"1f",	--2250
		x"06",	--2251
		x"3e",	--2252
		x"1e",	--2253
		x"0e",	--2254
		x"81",	--2255
		x"02",	--2256
		x"d7",	--2257
		x"91",	--2258
		x"04",	--2259
		x"04",	--2260
		x"91",	--2261
		x"06",	--2262
		x"06",	--2263
		x"7e",	--2264
		x"f8",	--2265
		x"f1",	--2266
		x"0e",	--2267
		x"3e",	--2268
		x"1e",	--2269
		x"1c",	--2270
		x"0d",	--2271
		x"48",	--2272
		x"78",	--2273
		x"1f",	--2274
		x"04",	--2275
		x"0c",	--2276
		x"0d",	--2277
		x"78",	--2278
		x"fc",	--2279
		x"3c",	--2280
		x"3d",	--2281
		x"0c",	--2282
		x"0d",	--2283
		x"18",	--2284
		x"09",	--2285
		x"0c",	--2286
		x"04",	--2287
		x"0d",	--2288
		x"02",	--2289
		x"08",	--2290
		x"09",	--2291
		x"7e",	--2292
		x"1f",	--2293
		x"0e",	--2294
		x"0d",	--2295
		x"0e",	--2296
		x"0d",	--2297
		x"0e",	--2298
		x"81",	--2299
		x"04",	--2300
		x"81",	--2301
		x"06",	--2302
		x"3e",	--2303
		x"1e",	--2304
		x"0e",	--2305
		x"81",	--2306
		x"02",	--2307
		x"a4",	--2308
		x"12",	--2309
		x"0b",	--2310
		x"0a",	--2311
		x"7e",	--2312
		x"fb",	--2313
		x"ec",	--2314
		x"0b",	--2315
		x"0a",	--2316
		x"09",	--2317
		x"1f",	--2318
		x"17",	--2319
		x"3e",	--2320
		x"00",	--2321
		x"2c",	--2322
		x"3a",	--2323
		x"18",	--2324
		x"0b",	--2325
		x"39",	--2326
		x"0c",	--2327
		x"0d",	--2328
		x"4f",	--2329
		x"4f",	--2330
		x"17",	--2331
		x"3c",	--2332
		x"d0",	--2333
		x"6e",	--2334
		x"0f",	--2335
		x"0a",	--2336
		x"0b",	--2337
		x"0f",	--2338
		x"39",	--2339
		x"3a",	--2340
		x"3b",	--2341
		x"30",	--2342
		x"3f",	--2343
		x"00",	--2344
		x"0f",	--2345
		x"3a",	--2346
		x"0b",	--2347
		x"39",	--2348
		x"18",	--2349
		x"0c",	--2350
		x"0d",	--2351
		x"4f",	--2352
		x"4f",	--2353
		x"e9",	--2354
		x"12",	--2355
		x"0d",	--2356
		x"0c",	--2357
		x"7f",	--2358
		x"fb",	--2359
		x"e3",	--2360
		x"3a",	--2361
		x"10",	--2362
		x"0b",	--2363
		x"39",	--2364
		x"10",	--2365
		x"ef",	--2366
		x"3a",	--2367
		x"20",	--2368
		x"0b",	--2369
		x"09",	--2370
		x"ea",	--2371
		x"0b",	--2372
		x"0a",	--2373
		x"09",	--2374
		x"08",	--2375
		x"07",	--2376
		x"0d",	--2377
		x"1e",	--2378
		x"04",	--2379
		x"1f",	--2380
		x"06",	--2381
		x"5a",	--2382
		x"01",	--2383
		x"6c",	--2384
		x"6c",	--2385
		x"70",	--2386
		x"6c",	--2387
		x"6a",	--2388
		x"6c",	--2389
		x"36",	--2390
		x"0e",	--2391
		x"32",	--2392
		x"1b",	--2393
		x"02",	--2394
		x"3b",	--2395
		x"82",	--2396
		x"6d",	--2397
		x"3b",	--2398
		x"80",	--2399
		x"5e",	--2400
		x"0c",	--2401
		x"0d",	--2402
		x"3c",	--2403
		x"7f",	--2404
		x"0d",	--2405
		x"3c",	--2406
		x"40",	--2407
		x"40",	--2408
		x"3e",	--2409
		x"3f",	--2410
		x"0f",	--2411
		x"0f",	--2412
		x"4a",	--2413
		x"0d",	--2414
		x"3d",	--2415
		x"7f",	--2416
		x"12",	--2417
		x"0f",	--2418
		x"0e",	--2419
		x"12",	--2420
		x"0f",	--2421
		x"0e",	--2422
		x"12",	--2423
		x"0f",	--2424
		x"0e",	--2425
		x"12",	--2426
		x"0f",	--2427
		x"0e",	--2428
		x"12",	--2429
		x"0f",	--2430
		x"0e",	--2431
		x"12",	--2432
		x"0f",	--2433
		x"0e",	--2434
		x"12",	--2435
		x"0f",	--2436
		x"0e",	--2437
		x"3e",	--2438
		x"3f",	--2439
		x"7f",	--2440
		x"4d",	--2441
		x"05",	--2442
		x"0f",	--2443
		x"cc",	--2444
		x"4d",	--2445
		x"0e",	--2446
		x"0f",	--2447
		x"4d",	--2448
		x"0d",	--2449
		x"0d",	--2450
		x"0d",	--2451
		x"0d",	--2452
		x"0d",	--2453
		x"0d",	--2454
		x"0d",	--2455
		x"0c",	--2456
		x"3c",	--2457
		x"7f",	--2458
		x"0c",	--2459
		x"4f",	--2460
		x"0f",	--2461
		x"0f",	--2462
		x"0f",	--2463
		x"0d",	--2464
		x"0d",	--2465
		x"0f",	--2466
		x"37",	--2467
		x"38",	--2468
		x"39",	--2469
		x"3a",	--2470
		x"3b",	--2471
		x"30",	--2472
		x"0d",	--2473
		x"be",	--2474
		x"0c",	--2475
		x"0d",	--2476
		x"3c",	--2477
		x"80",	--2478
		x"0d",	--2479
		x"0c",	--2480
		x"02",	--2481
		x"0d",	--2482
		x"b8",	--2483
		x"3e",	--2484
		x"40",	--2485
		x"0f",	--2486
		x"b4",	--2487
		x"12",	--2488
		x"0f",	--2489
		x"0e",	--2490
		x"0d",	--2491
		x"3d",	--2492
		x"80",	--2493
		x"b2",	--2494
		x"7d",	--2495
		x"0e",	--2496
		x"0f",	--2497
		x"cd",	--2498
		x"0e",	--2499
		x"3f",	--2500
		x"10",	--2501
		x"3e",	--2502
		x"3f",	--2503
		x"7f",	--2504
		x"7d",	--2505
		x"c5",	--2506
		x"37",	--2507
		x"82",	--2508
		x"07",	--2509
		x"37",	--2510
		x"1a",	--2511
		x"4f",	--2512
		x"0c",	--2513
		x"0d",	--2514
		x"4b",	--2515
		x"7b",	--2516
		x"1f",	--2517
		x"05",	--2518
		x"12",	--2519
		x"0d",	--2520
		x"0c",	--2521
		x"7b",	--2522
		x"fb",	--2523
		x"18",	--2524
		x"09",	--2525
		x"77",	--2526
		x"1f",	--2527
		x"04",	--2528
		x"08",	--2529
		x"09",	--2530
		x"77",	--2531
		x"fc",	--2532
		x"38",	--2533
		x"39",	--2534
		x"08",	--2535
		x"09",	--2536
		x"1e",	--2537
		x"0f",	--2538
		x"08",	--2539
		x"04",	--2540
		x"09",	--2541
		x"02",	--2542
		x"0e",	--2543
		x"0f",	--2544
		x"08",	--2545
		x"09",	--2546
		x"08",	--2547
		x"09",	--2548
		x"0e",	--2549
		x"0f",	--2550
		x"3e",	--2551
		x"7f",	--2552
		x"0f",	--2553
		x"3e",	--2554
		x"40",	--2555
		x"26",	--2556
		x"38",	--2557
		x"3f",	--2558
		x"09",	--2559
		x"0e",	--2560
		x"0f",	--2561
		x"12",	--2562
		x"0f",	--2563
		x"0e",	--2564
		x"12",	--2565
		x"0f",	--2566
		x"0e",	--2567
		x"12",	--2568
		x"0f",	--2569
		x"0e",	--2570
		x"12",	--2571
		x"0f",	--2572
		x"0e",	--2573
		x"12",	--2574
		x"0f",	--2575
		x"0e",	--2576
		x"12",	--2577
		x"0f",	--2578
		x"0e",	--2579
		x"12",	--2580
		x"0f",	--2581
		x"0e",	--2582
		x"3e",	--2583
		x"3f",	--2584
		x"7f",	--2585
		x"5d",	--2586
		x"39",	--2587
		x"00",	--2588
		x"72",	--2589
		x"4d",	--2590
		x"70",	--2591
		x"08",	--2592
		x"09",	--2593
		x"da",	--2594
		x"0f",	--2595
		x"d8",	--2596
		x"0e",	--2597
		x"0f",	--2598
		x"3e",	--2599
		x"80",	--2600
		x"0f",	--2601
		x"0e",	--2602
		x"04",	--2603
		x"38",	--2604
		x"40",	--2605
		x"09",	--2606
		x"d0",	--2607
		x"0f",	--2608
		x"ce",	--2609
		x"f9",	--2610
		x"0b",	--2611
		x"0a",	--2612
		x"2a",	--2613
		x"5b",	--2614
		x"02",	--2615
		x"3b",	--2616
		x"7f",	--2617
		x"1d",	--2618
		x"02",	--2619
		x"12",	--2620
		x"0d",	--2621
		x"12",	--2622
		x"0d",	--2623
		x"12",	--2624
		x"0d",	--2625
		x"12",	--2626
		x"0d",	--2627
		x"12",	--2628
		x"0d",	--2629
		x"12",	--2630
		x"0d",	--2631
		x"12",	--2632
		x"0d",	--2633
		x"4d",	--2634
		x"5f",	--2635
		x"03",	--2636
		x"3f",	--2637
		x"80",	--2638
		x"0f",	--2639
		x"0f",	--2640
		x"ce",	--2641
		x"01",	--2642
		x"0d",	--2643
		x"2d",	--2644
		x"0a",	--2645
		x"51",	--2646
		x"be",	--2647
		x"82",	--2648
		x"02",	--2649
		x"0c",	--2650
		x"0d",	--2651
		x"0c",	--2652
		x"0d",	--2653
		x"0c",	--2654
		x"0d",	--2655
		x"0c",	--2656
		x"0d",	--2657
		x"0c",	--2658
		x"0d",	--2659
		x"0c",	--2660
		x"0d",	--2661
		x"0c",	--2662
		x"0d",	--2663
		x"0c",	--2664
		x"0d",	--2665
		x"fe",	--2666
		x"03",	--2667
		x"00",	--2668
		x"3d",	--2669
		x"00",	--2670
		x"0b",	--2671
		x"3f",	--2672
		x"81",	--2673
		x"0c",	--2674
		x"0d",	--2675
		x"0a",	--2676
		x"3f",	--2677
		x"3d",	--2678
		x"00",	--2679
		x"f9",	--2680
		x"8e",	--2681
		x"02",	--2682
		x"8e",	--2683
		x"04",	--2684
		x"8e",	--2685
		x"06",	--2686
		x"3a",	--2687
		x"3b",	--2688
		x"30",	--2689
		x"3d",	--2690
		x"ff",	--2691
		x"2a",	--2692
		x"3d",	--2693
		x"81",	--2694
		x"8e",	--2695
		x"02",	--2696
		x"fe",	--2697
		x"03",	--2698
		x"00",	--2699
		x"0c",	--2700
		x"0d",	--2701
		x"0c",	--2702
		x"0d",	--2703
		x"0c",	--2704
		x"0d",	--2705
		x"0c",	--2706
		x"0d",	--2707
		x"0c",	--2708
		x"0d",	--2709
		x"0c",	--2710
		x"0d",	--2711
		x"0c",	--2712
		x"0d",	--2713
		x"0c",	--2714
		x"0d",	--2715
		x"0a",	--2716
		x"0b",	--2717
		x"0a",	--2718
		x"3b",	--2719
		x"00",	--2720
		x"8e",	--2721
		x"04",	--2722
		x"8e",	--2723
		x"06",	--2724
		x"3a",	--2725
		x"3b",	--2726
		x"30",	--2727
		x"0b",	--2728
		x"ad",	--2729
		x"ee",	--2730
		x"00",	--2731
		x"3a",	--2732
		x"3b",	--2733
		x"30",	--2734
		x"0a",	--2735
		x"0c",	--2736
		x"0c",	--2737
		x"0d",	--2738
		x"0c",	--2739
		x"3d",	--2740
		x"10",	--2741
		x"0c",	--2742
		x"02",	--2743
		x"0d",	--2744
		x"08",	--2745
		x"de",	--2746
		x"00",	--2747
		x"e4",	--2748
		x"0b",	--2749
		x"f2",	--2750
		x"ee",	--2751
		x"00",	--2752
		x"e3",	--2753
		x"ce",	--2754
		x"00",	--2755
		x"dc",	--2756
		x"0b",	--2757
		x"6d",	--2758
		x"6d",	--2759
		x"12",	--2760
		x"6c",	--2761
		x"6c",	--2762
		x"0f",	--2763
		x"6d",	--2764
		x"41",	--2765
		x"6c",	--2766
		x"11",	--2767
		x"6d",	--2768
		x"0d",	--2769
		x"6c",	--2770
		x"14",	--2771
		x"5d",	--2772
		x"01",	--2773
		x"5d",	--2774
		x"01",	--2775
		x"14",	--2776
		x"4d",	--2777
		x"09",	--2778
		x"1e",	--2779
		x"0f",	--2780
		x"3b",	--2781
		x"30",	--2782
		x"6c",	--2783
		x"28",	--2784
		x"ce",	--2785
		x"01",	--2786
		x"f7",	--2787
		x"3e",	--2788
		x"0f",	--2789
		x"3b",	--2790
		x"30",	--2791
		x"cf",	--2792
		x"01",	--2793
		x"f0",	--2794
		x"3e",	--2795
		x"f8",	--2796
		x"1b",	--2797
		x"02",	--2798
		x"1c",	--2799
		x"02",	--2800
		x"0c",	--2801
		x"e6",	--2802
		x"0b",	--2803
		x"16",	--2804
		x"1b",	--2805
		x"04",	--2806
		x"1f",	--2807
		x"06",	--2808
		x"1c",	--2809
		x"04",	--2810
		x"1e",	--2811
		x"06",	--2812
		x"0e",	--2813
		x"da",	--2814
		x"0f",	--2815
		x"02",	--2816
		x"0c",	--2817
		x"d6",	--2818
		x"0f",	--2819
		x"06",	--2820
		x"0e",	--2821
		x"02",	--2822
		x"0b",	--2823
		x"02",	--2824
		x"0e",	--2825
		x"d1",	--2826
		x"4d",	--2827
		x"ce",	--2828
		x"3e",	--2829
		x"d6",	--2830
		x"6c",	--2831
		x"d7",	--2832
		x"5e",	--2833
		x"01",	--2834
		x"5f",	--2835
		x"01",	--2836
		x"0e",	--2837
		x"c5",	--2838
		x"0d",	--2839
		x"0f",	--2840
		x"04",	--2841
		x"3d",	--2842
		x"03",	--2843
		x"3f",	--2844
		x"1f",	--2845
		x"0e",	--2846
		x"03",	--2847
		x"5d",	--2848
		x"3e",	--2849
		x"1e",	--2850
		x"0d",	--2851
		x"b0",	--2852
		x"b4",	--2853
		x"3d",	--2854
		x"6d",	--2855
		x"02",	--2856
		x"3e",	--2857
		x"1e",	--2858
		x"5d",	--2859
		x"02",	--2860
		x"3f",	--2861
		x"1f",	--2862
		x"30",	--2863
		x"b0",	--2864
		x"2e",	--2865
		x"0f",	--2866
		x"30",	--2867
		x"0b",	--2868
		x"0b",	--2869
		x"0f",	--2870
		x"06",	--2871
		x"3b",	--2872
		x"03",	--2873
		x"3e",	--2874
		x"3f",	--2875
		x"1e",	--2876
		x"0f",	--2877
		x"0d",	--2878
		x"05",	--2879
		x"5b",	--2880
		x"3c",	--2881
		x"3d",	--2882
		x"1c",	--2883
		x"0d",	--2884
		x"b0",	--2885
		x"d6",	--2886
		x"6b",	--2887
		x"04",	--2888
		x"3c",	--2889
		x"3d",	--2890
		x"1c",	--2891
		x"0d",	--2892
		x"5b",	--2893
		x"04",	--2894
		x"3e",	--2895
		x"3f",	--2896
		x"1e",	--2897
		x"0f",	--2898
		x"3b",	--2899
		x"30",	--2900
		x"b0",	--2901
		x"68",	--2902
		x"0e",	--2903
		x"0f",	--2904
		x"30",	--2905
		x"7c",	--2906
		x"10",	--2907
		x"0d",	--2908
		x"0e",	--2909
		x"0f",	--2910
		x"0e",	--2911
		x"0e",	--2912
		x"02",	--2913
		x"0e",	--2914
		x"1f",	--2915
		x"1c",	--2916
		x"f8",	--2917
		x"30",	--2918
		x"b0",	--2919
		x"b4",	--2920
		x"0f",	--2921
		x"30",	--2922
		x"0b",	--2923
		x"0a",	--2924
		x"09",	--2925
		x"79",	--2926
		x"20",	--2927
		x"0a",	--2928
		x"0b",	--2929
		x"0c",	--2930
		x"0d",	--2931
		x"0e",	--2932
		x"0f",	--2933
		x"0c",	--2934
		x"0d",	--2935
		x"0d",	--2936
		x"06",	--2937
		x"02",	--2938
		x"0c",	--2939
		x"03",	--2940
		x"0c",	--2941
		x"0d",	--2942
		x"1e",	--2943
		x"19",	--2944
		x"f2",	--2945
		x"39",	--2946
		x"3a",	--2947
		x"3b",	--2948
		x"30",	--2949
		x"b0",	--2950
		x"d6",	--2951
		x"0e",	--2952
		x"0f",	--2953
		x"30",	--2954
		x"00",	--2955
		x"32",	--2956
		x"f0",	--2957
		x"fd",	--2958
		x"63",	--2959
		x"72",	--2960
		x"65",	--2961
		x"74",	--2962
		x"75",	--2963
		x"61",	--2964
		x"65",	--2965
		x"0d",	--2966
		x"00",	--2967
		x"25",	--2968
		x"20",	--2969
		x"45",	--2970
		x"54",	--2971
		x"52",	--2972
		x"47",	--2973
		x"54",	--2974
		x"0a",	--2975
		x"53",	--2976
		x"6d",	--2977
		x"74",	--2978
		x"69",	--2979
		x"67",	--2980
		x"77",	--2981
		x"6e",	--2982
		x"20",	--2983
		x"65",	--2984
		x"72",	--2985
		x"62",	--2986
		x"79",	--2987
		x"77",	--2988
		x"6f",	--2989
		x"67",	--2990
		x"0a",	--2991
		x"3e",	--2992
		x"00",	--2993
		x"0a",	--2994
		x"3a",	--2995
		x"73",	--2996
		x"0a",	--2997
		x"08",	--2998
		x"08",	--2999
		x"25",	--3000
		x"00",	--3001
		x"72",	--3002
		x"74",	--3003
		x"0a",	--3004
		x"00",	--3005
		x"6f",	--3006
		x"72",	--3007
		x"63",	--3008
		x"20",	--3009
		x"73",	--3010
		x"67",	--3011
		x"3a",	--3012
		x"0a",	--3013
		x"09",	--3014
		x"63",	--3015
		x"52",	--3016
		x"47",	--3017
		x"53",	--3018
		x"45",	--3019
		x"20",	--3020
		x"41",	--3021
		x"55",	--3022
		x"0d",	--3023
		x"00",	--3024
		x"6f",	--3025
		x"65",	--3026
		x"68",	--3027
		x"6e",	--3028
		x"20",	--3029
		x"65",	--3030
		x"74",	--3031
		x"74",	--3032
		x"72",	--3033
		x"69",	--3034
		x"6c",	--3035
		x"20",	--3036
		x"72",	--3037
		x"6e",	--3038
		x"0d",	--3039
		x"00",	--3040
		x"3d",	--3041
		x"64",	--3042
		x"76",	--3043
		x"25",	--3044
		x"0d",	--3045
		x"00",	--3046
		x"65",	--3047
		x"64",	--3048
		x"0d",	--3049
		x"09",	--3050
		x"63",	--3051
		x"52",	--3052
		x"47",	--3053
		x"53",	--3054
		x"45",	--3055
		x"0d",	--3056
		x"00",	--3057
		x"63",	--3058
		x"69",	--3059
		x"20",	--3060
		x"6f",	--3061
		x"20",	--3062
		x"20",	--3063
		x"75",	--3064
		x"62",	--3065
		x"72",	--3066
		x"0a",	--3067
		x"25",	--3068
		x"3a",	--3069
		x"6e",	--3070
		x"20",	--3071
		x"75",	--3072
		x"68",	--3073
		x"63",	--3074
		x"6d",	--3075
		x"61",	--3076
		x"64",	--3077
		x"0a",	--3078
		x"b8",	--3079
		x"e6",	--3080
		x"e6",	--3081
		x"e6",	--3082
		x"e6",	--3083
		x"e6",	--3084
		x"e6",	--3085
		x"e6",	--3086
		x"e6",	--3087
		x"e6",	--3088
		x"e6",	--3089
		x"e6",	--3090
		x"e6",	--3091
		x"e6",	--3092
		x"e6",	--3093
		x"e6",	--3094
		x"e6",	--3095
		x"e6",	--3096
		x"e6",	--3097
		x"e6",	--3098
		x"e6",	--3099
		x"e6",	--3100
		x"e6",	--3101
		x"e6",	--3102
		x"e6",	--3103
		x"e6",	--3104
		x"e6",	--3105
		x"e6",	--3106
		x"e6",	--3107
		x"aa",	--3108
		x"e6",	--3109
		x"e6",	--3110
		x"e6",	--3111
		x"e6",	--3112
		x"e6",	--3113
		x"e6",	--3114
		x"e6",	--3115
		x"e6",	--3116
		x"e6",	--3117
		x"e6",	--3118
		x"e6",	--3119
		x"e6",	--3120
		x"e6",	--3121
		x"e6",	--3122
		x"e6",	--3123
		x"e6",	--3124
		x"e6",	--3125
		x"e6",	--3126
		x"e6",	--3127
		x"e6",	--3128
		x"e6",	--3129
		x"e6",	--3130
		x"e6",	--3131
		x"e6",	--3132
		x"e6",	--3133
		x"e6",	--3134
		x"e6",	--3135
		x"e6",	--3136
		x"e6",	--3137
		x"e6",	--3138
		x"e6",	--3139
		x"9c",	--3140
		x"8e",	--3141
		x"80",	--3142
		x"e6",	--3143
		x"e6",	--3144
		x"e6",	--3145
		x"e6",	--3146
		x"e6",	--3147
		x"e6",	--3148
		x"e6",	--3149
		x"68",	--3150
		x"e6",	--3151
		x"56",	--3152
		x"e6",	--3153
		x"e6",	--3154
		x"e6",	--3155
		x"e6",	--3156
		x"3a",	--3157
		x"e6",	--3158
		x"e6",	--3159
		x"e6",	--3160
		x"2c",	--3161
		x"1a",	--3162
		x"30",	--3163
		x"32",	--3164
		x"34",	--3165
		x"36",	--3166
		x"38",	--3167
		x"61",	--3168
		x"63",	--3169
		x"65",	--3170
		x"00",	--3171
		x"00",	--3172
		x"00",	--3173
		x"00",	--3174
		x"00",	--3175
		x"00",	--3176
		x"02",	--3177
		x"03",	--3178
		x"03",	--3179
		x"04",	--3180
		x"04",	--3181
		x"04",	--3182
		x"04",	--3183
		x"05",	--3184
		x"05",	--3185
		x"05",	--3186
		x"05",	--3187
		x"05",	--3188
		x"05",	--3189
		x"05",	--3190
		x"05",	--3191
		x"06",	--3192
		x"06",	--3193
		x"06",	--3194
		x"06",	--3195
		x"06",	--3196
		x"06",	--3197
		x"06",	--3198
		x"06",	--3199
		x"06",	--3200
		x"06",	--3201
		x"06",	--3202
		x"06",	--3203
		x"06",	--3204
		x"06",	--3205
		x"06",	--3206
		x"06",	--3207
		x"07",	--3208
		x"07",	--3209
		x"07",	--3210
		x"07",	--3211
		x"07",	--3212
		x"07",	--3213
		x"07",	--3214
		x"07",	--3215
		x"07",	--3216
		x"07",	--3217
		x"07",	--3218
		x"07",	--3219
		x"07",	--3220
		x"07",	--3221
		x"07",	--3222
		x"07",	--3223
		x"07",	--3224
		x"07",	--3225
		x"07",	--3226
		x"07",	--3227
		x"07",	--3228
		x"07",	--3229
		x"07",	--3230
		x"07",	--3231
		x"07",	--3232
		x"07",	--3233
		x"07",	--3234
		x"07",	--3235
		x"07",	--3236
		x"07",	--3237
		x"07",	--3238
		x"07",	--3239
		x"08",	--3240
		x"08",	--3241
		x"08",	--3242
		x"08",	--3243
		x"08",	--3244
		x"08",	--3245
		x"08",	--3246
		x"08",	--3247
		x"08",	--3248
		x"08",	--3249
		x"08",	--3250
		x"08",	--3251
		x"08",	--3252
		x"08",	--3253
		x"08",	--3254
		x"08",	--3255
		x"08",	--3256
		x"08",	--3257
		x"08",	--3258
		x"08",	--3259
		x"08",	--3260
		x"08",	--3261
		x"08",	--3262
		x"08",	--3263
		x"08",	--3264
		x"08",	--3265
		x"08",	--3266
		x"08",	--3267
		x"08",	--3268
		x"08",	--3269
		x"08",	--3270
		x"08",	--3271
		x"08",	--3272
		x"08",	--3273
		x"08",	--3274
		x"08",	--3275
		x"08",	--3276
		x"08",	--3277
		x"08",	--3278
		x"08",	--3279
		x"08",	--3280
		x"08",	--3281
		x"08",	--3282
		x"08",	--3283
		x"08",	--3284
		x"08",	--3285
		x"08",	--3286
		x"08",	--3287
		x"08",	--3288
		x"08",	--3289
		x"08",	--3290
		x"08",	--3291
		x"08",	--3292
		x"08",	--3293
		x"08",	--3294
		x"08",	--3295
		x"08",	--3296
		x"08",	--3297
		x"08",	--3298
		x"08",	--3299
		x"08",	--3300
		x"08",	--3301
		x"08",	--3302
		x"08",	--3303
		x"ff",	--3304
		x"ff",	--3305
		x"ff",	--3306
		x"ff",	--3307
		x"ff",	--3308
		x"ff",	--3309
		x"ff",	--3310
		x"ff",	--3311
		x"ff",	--3312
		x"ff",	--3313
		x"ff",	--3314
		x"ff",	--3315
		x"ff",	--3316
		x"ff",	--3317
		x"ff",	--3318
		x"ff",	--3319
		x"ff",	--3320
		x"ff",	--3321
		x"ff",	--3322
		x"ff",	--3323
		x"ff",	--3324
		x"ff",	--3325
		x"ff",	--3326
		x"ff",	--3327
		x"ff",	--3328
		x"ff",	--3329
		x"ff",	--3330
		x"ff",	--3331
		x"ff",	--3332
		x"ff",	--3333
		x"ff",	--3334
		x"ff",	--3335
		x"ff",	--3336
		x"ff",	--3337
		x"ff",	--3338
		x"ff",	--3339
		x"ff",	--3340
		x"ff",	--3341
		x"ff",	--3342
		x"ff",	--3343
		x"ff",	--3344
		x"ff",	--3345
		x"ff",	--3346
		x"ff",	--3347
		x"ff",	--3348
		x"ff",	--3349
		x"ff",	--3350
		x"ff",	--3351
		x"ff",	--3352
		x"ff",	--3353
		x"ff",	--3354
		x"ff",	--3355
		x"ff",	--3356
		x"ff",	--3357
		x"ff",	--3358
		x"ff",	--3359
		x"ff",	--3360
		x"ff",	--3361
		x"ff",	--3362
		x"ff",	--3363
		x"ff",	--3364
		x"ff",	--3365
		x"ff",	--3366
		x"ff",	--3367
		x"ff",	--3368
		x"ff",	--3369
		x"ff",	--3370
		x"ff",	--3371
		x"ff",	--3372
		x"ff",	--3373
		x"ff",	--3374
		x"ff",	--3375
		x"ff",	--3376
		x"ff",	--3377
		x"ff",	--3378
		x"ff",	--3379
		x"ff",	--3380
		x"ff",	--3381
		x"ff",	--3382
		x"ff",	--3383
		x"ff",	--3384
		x"ff",	--3385
		x"ff",	--3386
		x"ff",	--3387
		x"ff",	--3388
		x"ff",	--3389
		x"ff",	--3390
		x"ff",	--3391
		x"ff",	--3392
		x"ff",	--3393
		x"ff",	--3394
		x"ff",	--3395
		x"ff",	--3396
		x"ff",	--3397
		x"ff",	--3398
		x"ff",	--3399
		x"ff",	--3400
		x"ff",	--3401
		x"ff",	--3402
		x"ff",	--3403
		x"ff",	--3404
		x"ff",	--3405
		x"ff",	--3406
		x"ff",	--3407
		x"ff",	--3408
		x"ff",	--3409
		x"ff",	--3410
		x"ff",	--3411
		x"ff",	--3412
		x"ff",	--3413
		x"ff",	--3414
		x"ff",	--3415
		x"ff",	--3416
		x"ff",	--3417
		x"ff",	--3418
		x"ff",	--3419
		x"ff",	--3420
		x"ff",	--3421
		x"ff",	--3422
		x"ff",	--3423
		x"ff",	--3424
		x"ff",	--3425
		x"ff",	--3426
		x"ff",	--3427
		x"ff",	--3428
		x"ff",	--3429
		x"ff",	--3430
		x"ff",	--3431
		x"ff",	--3432
		x"ff",	--3433
		x"ff",	--3434
		x"ff",	--3435
		x"ff",	--3436
		x"ff",	--3437
		x"ff",	--3438
		x"ff",	--3439
		x"ff",	--3440
		x"ff",	--3441
		x"ff",	--3442
		x"ff",	--3443
		x"ff",	--3444
		x"ff",	--3445
		x"ff",	--3446
		x"ff",	--3447
		x"ff",	--3448
		x"ff",	--3449
		x"ff",	--3450
		x"ff",	--3451
		x"ff",	--3452
		x"ff",	--3453
		x"ff",	--3454
		x"ff",	--3455
		x"ff",	--3456
		x"ff",	--3457
		x"ff",	--3458
		x"ff",	--3459
		x"ff",	--3460
		x"ff",	--3461
		x"ff",	--3462
		x"ff",	--3463
		x"ff",	--3464
		x"ff",	--3465
		x"ff",	--3466
		x"ff",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"8c",	--4080
		x"8c",	--4081
		x"8c",	--4082
		x"8c",	--4083
		x"8c",	--4084
		x"8c",	--4085
		x"8c",	--4086
		x"c2",	--4087
		x"8c",	--4088
		x"8c",	--4089
		x"8c",	--4090
		x"8c",	--4091
		x"8c",	--4092
		x"8c",	--4093
		x"8c",	--4094
		x"00");	--4095
	constant mcu_firmware_h : ram8_t := (
		x"42",	--0
		x"01",	--1
		x"d0",	--2
		x"5a",	--3
		x"45",	--4
		x"03",	--5
		x"40",	--6
		x"06",	--7
		x"40",	--8
		x"00",	--9
		x"93",	--10
		x"24",	--11
		x"42",	--12
		x"03",	--13
		x"01",	--14
		x"83",	--15
		x"4f",	--16
		x"f9",	--17
		x"02",	--18
		x"23",	--19
		x"40",	--20
		x"01",	--21
		x"93",	--22
		x"24",	--23
		x"42",	--24
		x"03",	--25
		x"01",	--26
		x"83",	--27
		x"43",	--28
		x"02",	--29
		x"23",	--30
		x"50",	--31
		x"ff",	--32
		x"40",	--33
		x"5a",	--34
		x"01",	--35
		x"43",	--36
		x"00",	--37
		x"43",	--38
		x"00",	--39
		x"40",	--40
		x"c2",	--41
		x"43",	--42
		x"12",	--43
		x"e9",	--44
		x"12",	--45
		x"e5",	--46
		x"43",	--47
		x"00",	--48
		x"40",	--49
		x"e2",	--50
		x"40",	--51
		x"00",	--52
		x"12",	--53
		x"e5",	--54
		x"40",	--55
		x"e2",	--56
		x"40",	--57
		x"00",	--58
		x"12",	--59
		x"e5",	--60
		x"40",	--61
		x"e1",	--62
		x"40",	--63
		x"00",	--64
		x"12",	--65
		x"e5",	--66
		x"43",	--67
		x"40",	--68
		x"4e",	--69
		x"40",	--70
		x"01",	--71
		x"41",	--72
		x"50",	--73
		x"00",	--74
		x"12",	--75
		x"e4",	--76
		x"41",	--77
		x"50",	--78
		x"00",	--79
		x"12",	--80
		x"e4",	--81
		x"43",	--82
		x"40",	--83
		x"4e",	--84
		x"40",	--85
		x"01",	--86
		x"41",	--87
		x"12",	--88
		x"e4",	--89
		x"41",	--90
		x"12",	--91
		x"e4",	--92
		x"41",	--93
		x"41",	--94
		x"50",	--95
		x"00",	--96
		x"12",	--97
		x"e1",	--98
		x"40",	--99
		x"ff",	--100
		x"00",	--101
		x"d2",	--102
		x"43",	--103
		x"12",	--104
		x"f7",	--105
		x"12",	--106
		x"e7",	--107
		x"53",	--108
		x"43",	--109
		x"d0",	--110
		x"00",	--111
		x"53",	--112
		x"90",	--113
		x"00",	--114
		x"24",	--115
		x"43",	--116
		x"4b",	--117
		x"f0",	--118
		x"00",	--119
		x"24",	--120
		x"5f",	--121
		x"53",	--122
		x"23",	--123
		x"4f",	--124
		x"3c",	--125
		x"43",	--126
		x"43",	--127
		x"4f",	--128
		x"00",	--129
		x"12",	--130
		x"e9",	--131
		x"93",	--132
		x"27",	--133
		x"12",	--134
		x"e9",	--135
		x"92",	--136
		x"24",	--137
		x"90",	--138
		x"00",	--139
		x"20",	--140
		x"12",	--141
		x"f7",	--142
		x"12",	--143
		x"e7",	--144
		x"53",	--145
		x"40",	--146
		x"00",	--147
		x"51",	--148
		x"5f",	--149
		x"43",	--150
		x"00",	--151
		x"12",	--152
		x"12",	--153
		x"f7",	--154
		x"12",	--155
		x"e7",	--156
		x"52",	--157
		x"41",	--158
		x"50",	--159
		x"00",	--160
		x"41",	--161
		x"00",	--162
		x"12",	--163
		x"e5",	--164
		x"3f",	--165
		x"93",	--166
		x"27",	--167
		x"53",	--168
		x"12",	--169
		x"f7",	--170
		x"12",	--171
		x"e7",	--172
		x"53",	--173
		x"3f",	--174
		x"90",	--175
		x"00",	--176
		x"2f",	--177
		x"4f",	--178
		x"11",	--179
		x"12",	--180
		x"12",	--181
		x"f7",	--182
		x"4f",	--183
		x"00",	--184
		x"12",	--185
		x"e7",	--186
		x"52",	--187
		x"40",	--188
		x"00",	--189
		x"51",	--190
		x"5a",	--191
		x"41",	--192
		x"00",	--193
		x"4f",	--194
		x"00",	--195
		x"53",	--196
		x"3f",	--197
		x"40",	--198
		x"f7",	--199
		x"4f",	--200
		x"02",	--201
		x"4e",	--202
		x"02",	--203
		x"41",	--204
		x"82",	--205
		x"90",	--206
		x"00",	--207
		x"00",	--208
		x"20",	--209
		x"93",	--210
		x"00",	--211
		x"24",	--212
		x"41",	--213
		x"4f",	--214
		x"53",	--215
		x"41",	--216
		x"52",	--217
		x"12",	--218
		x"e3",	--219
		x"93",	--220
		x"00",	--221
		x"24",	--222
		x"41",	--223
		x"4f",	--224
		x"41",	--225
		x"53",	--226
		x"12",	--227
		x"e3",	--228
		x"93",	--229
		x"00",	--230
		x"24",	--231
		x"41",	--232
		x"00",	--233
		x"43",	--234
		x"12",	--235
		x"f1",	--236
		x"43",	--237
		x"40",	--238
		x"42",	--239
		x"12",	--240
		x"ef",	--241
		x"4e",	--242
		x"4f",	--243
		x"42",	--244
		x"02",	--245
		x"12",	--246
		x"e5",	--247
		x"41",	--248
		x"00",	--249
		x"43",	--250
		x"12",	--251
		x"f1",	--252
		x"43",	--253
		x"40",	--254
		x"42",	--255
		x"12",	--256
		x"ef",	--257
		x"4e",	--258
		x"4f",	--259
		x"42",	--260
		x"02",	--261
		x"12",	--262
		x"e5",	--263
		x"43",	--264
		x"52",	--265
		x"41",	--266
		x"12",	--267
		x"f7",	--268
		x"4f",	--269
		x"00",	--270
		x"12",	--271
		x"e7",	--272
		x"41",	--273
		x"00",	--274
		x"4f",	--275
		x"11",	--276
		x"4f",	--277
		x"00",	--278
		x"12",	--279
		x"f7",	--280
		x"12",	--281
		x"e7",	--282
		x"52",	--283
		x"43",	--284
		x"52",	--285
		x"41",	--286
		x"12",	--287
		x"f7",	--288
		x"12",	--289
		x"e7",	--290
		x"53",	--291
		x"43",	--292
		x"3f",	--293
		x"12",	--294
		x"50",	--295
		x"ff",	--296
		x"4f",	--297
		x"12",	--298
		x"f7",	--299
		x"12",	--300
		x"e7",	--301
		x"53",	--302
		x"90",	--303
		x"00",	--304
		x"00",	--305
		x"20",	--306
		x"93",	--307
		x"00",	--308
		x"24",	--309
		x"41",	--310
		x"4b",	--311
		x"53",	--312
		x"41",	--313
		x"52",	--314
		x"12",	--315
		x"e3",	--316
		x"93",	--317
		x"00",	--318
		x"24",	--319
		x"41",	--320
		x"4f",	--321
		x"41",	--322
		x"53",	--323
		x"12",	--324
		x"e3",	--325
		x"93",	--326
		x"00",	--327
		x"24",	--328
		x"12",	--329
		x"00",	--330
		x"12",	--331
		x"00",	--332
		x"12",	--333
		x"f7",	--334
		x"12",	--335
		x"e7",	--336
		x"50",	--337
		x"00",	--338
		x"41",	--339
		x"00",	--340
		x"41",	--341
		x"00",	--342
		x"00",	--343
		x"43",	--344
		x"50",	--345
		x"00",	--346
		x"41",	--347
		x"41",	--348
		x"12",	--349
		x"f7",	--350
		x"12",	--351
		x"e7",	--352
		x"4b",	--353
		x"11",	--354
		x"4f",	--355
		x"00",	--356
		x"12",	--357
		x"f7",	--358
		x"12",	--359
		x"e7",	--360
		x"52",	--361
		x"43",	--362
		x"50",	--363
		x"00",	--364
		x"41",	--365
		x"41",	--366
		x"12",	--367
		x"f7",	--368
		x"12",	--369
		x"e7",	--370
		x"53",	--371
		x"43",	--372
		x"3f",	--373
		x"12",	--374
		x"82",	--375
		x"4f",	--376
		x"12",	--377
		x"f7",	--378
		x"12",	--379
		x"e7",	--380
		x"53",	--381
		x"90",	--382
		x"00",	--383
		x"00",	--384
		x"20",	--385
		x"93",	--386
		x"00",	--387
		x"24",	--388
		x"41",	--389
		x"4b",	--390
		x"53",	--391
		x"41",	--392
		x"53",	--393
		x"12",	--394
		x"e3",	--395
		x"93",	--396
		x"00",	--397
		x"24",	--398
		x"41",	--399
		x"00",	--400
		x"12",	--401
		x"12",	--402
		x"12",	--403
		x"f7",	--404
		x"12",	--405
		x"e7",	--406
		x"50",	--407
		x"00",	--408
		x"43",	--409
		x"52",	--410
		x"41",	--411
		x"41",	--412
		x"12",	--413
		x"f7",	--414
		x"12",	--415
		x"e7",	--416
		x"4b",	--417
		x"11",	--418
		x"4f",	--419
		x"00",	--420
		x"12",	--421
		x"f7",	--422
		x"12",	--423
		x"e7",	--424
		x"52",	--425
		x"43",	--426
		x"52",	--427
		x"41",	--428
		x"41",	--429
		x"12",	--430
		x"f7",	--431
		x"12",	--432
		x"e7",	--433
		x"53",	--434
		x"43",	--435
		x"3f",	--436
		x"12",	--437
		x"12",	--438
		x"12",	--439
		x"12",	--440
		x"12",	--441
		x"43",	--442
		x"00",	--443
		x"43",	--444
		x"00",	--445
		x"4e",	--446
		x"93",	--447
		x"24",	--448
		x"4e",	--449
		x"53",	--450
		x"4e",	--451
		x"43",	--452
		x"43",	--453
		x"43",	--454
		x"3c",	--455
		x"90",	--456
		x"00",	--457
		x"2c",	--458
		x"4f",	--459
		x"5c",	--460
		x"5c",	--461
		x"5c",	--462
		x"5c",	--463
		x"4c",	--464
		x"00",	--465
		x"50",	--466
		x"ff",	--467
		x"48",	--468
		x"11",	--469
		x"5a",	--470
		x"4c",	--471
		x"00",	--472
		x"43",	--473
		x"53",	--474
		x"49",	--475
		x"4b",	--476
		x"4b",	--477
		x"93",	--478
		x"24",	--479
		x"90",	--480
		x"00",	--481
		x"24",	--482
		x"90",	--483
		x"00",	--484
		x"24",	--485
		x"4c",	--486
		x"50",	--487
		x"ff",	--488
		x"93",	--489
		x"23",	--490
		x"90",	--491
		x"00",	--492
		x"2c",	--493
		x"4f",	--494
		x"5a",	--495
		x"4a",	--496
		x"5c",	--497
		x"5c",	--498
		x"5a",	--499
		x"4c",	--500
		x"00",	--501
		x"50",	--502
		x"ff",	--503
		x"48",	--504
		x"11",	--505
		x"58",	--506
		x"4c",	--507
		x"00",	--508
		x"3f",	--509
		x"43",	--510
		x"3f",	--511
		x"4c",	--512
		x"50",	--513
		x"ff",	--514
		x"90",	--515
		x"00",	--516
		x"2c",	--517
		x"4f",	--518
		x"5c",	--519
		x"5c",	--520
		x"5c",	--521
		x"5c",	--522
		x"4c",	--523
		x"00",	--524
		x"50",	--525
		x"ff",	--526
		x"3f",	--527
		x"4c",	--528
		x"50",	--529
		x"ff",	--530
		x"90",	--531
		x"00",	--532
		x"2c",	--533
		x"4f",	--534
		x"5c",	--535
		x"5c",	--536
		x"5c",	--537
		x"5c",	--538
		x"4c",	--539
		x"00",	--540
		x"50",	--541
		x"ff",	--542
		x"3f",	--543
		x"43",	--544
		x"00",	--545
		x"43",	--546
		x"41",	--547
		x"41",	--548
		x"41",	--549
		x"41",	--550
		x"41",	--551
		x"41",	--552
		x"43",	--553
		x"00",	--554
		x"4a",	--555
		x"53",	--556
		x"5e",	--557
		x"41",	--558
		x"41",	--559
		x"41",	--560
		x"41",	--561
		x"41",	--562
		x"41",	--563
		x"11",	--564
		x"12",	--565
		x"12",	--566
		x"f7",	--567
		x"12",	--568
		x"e7",	--569
		x"52",	--570
		x"43",	--571
		x"41",	--572
		x"41",	--573
		x"41",	--574
		x"41",	--575
		x"41",	--576
		x"41",	--577
		x"12",	--578
		x"12",	--579
		x"4e",	--580
		x"4c",	--581
		x"4e",	--582
		x"00",	--583
		x"4d",	--584
		x"00",	--585
		x"4c",	--586
		x"00",	--587
		x"4d",	--588
		x"43",	--589
		x"40",	--590
		x"36",	--591
		x"40",	--592
		x"01",	--593
		x"12",	--594
		x"f6",	--595
		x"4e",	--596
		x"00",	--597
		x"12",	--598
		x"c2",	--599
		x"43",	--600
		x"4a",	--601
		x"01",	--602
		x"40",	--603
		x"00",	--604
		x"01",	--605
		x"42",	--606
		x"01",	--607
		x"00",	--608
		x"41",	--609
		x"43",	--610
		x"41",	--611
		x"41",	--612
		x"41",	--613
		x"12",	--614
		x"12",	--615
		x"12",	--616
		x"43",	--617
		x"00",	--618
		x"40",	--619
		x"3f",	--620
		x"00",	--621
		x"4f",	--622
		x"4b",	--623
		x"00",	--624
		x"43",	--625
		x"12",	--626
		x"f1",	--627
		x"43",	--628
		x"40",	--629
		x"3f",	--630
		x"12",	--631
		x"ec",	--632
		x"4e",	--633
		x"4f",	--634
		x"4b",	--635
		x"00",	--636
		x"43",	--637
		x"12",	--638
		x"f1",	--639
		x"4e",	--640
		x"4f",	--641
		x"48",	--642
		x"49",	--643
		x"12",	--644
		x"ec",	--645
		x"12",	--646
		x"e9",	--647
		x"4e",	--648
		x"00",	--649
		x"43",	--650
		x"00",	--651
		x"41",	--652
		x"41",	--653
		x"41",	--654
		x"41",	--655
		x"12",	--656
		x"12",	--657
		x"12",	--658
		x"4d",	--659
		x"4e",	--660
		x"4d",	--661
		x"00",	--662
		x"4e",	--663
		x"00",	--664
		x"4f",	--665
		x"49",	--666
		x"00",	--667
		x"43",	--668
		x"12",	--669
		x"f1",	--670
		x"4e",	--671
		x"4f",	--672
		x"4a",	--673
		x"4b",	--674
		x"12",	--675
		x"ec",	--676
		x"4e",	--677
		x"4f",	--678
		x"49",	--679
		x"00",	--680
		x"43",	--681
		x"12",	--682
		x"f1",	--683
		x"4e",	--684
		x"4f",	--685
		x"4a",	--686
		x"4b",	--687
		x"12",	--688
		x"ec",	--689
		x"12",	--690
		x"e9",	--691
		x"4e",	--692
		x"00",	--693
		x"41",	--694
		x"41",	--695
		x"41",	--696
		x"41",	--697
		x"41",	--698
		x"42",	--699
		x"02",	--700
		x"90",	--701
		x"00",	--702
		x"34",	--703
		x"4c",	--704
		x"5d",	--705
		x"5d",	--706
		x"50",	--707
		x"02",	--708
		x"4f",	--709
		x"00",	--710
		x"4e",	--711
		x"00",	--712
		x"53",	--713
		x"4c",	--714
		x"02",	--715
		x"43",	--716
		x"41",	--717
		x"43",	--718
		x"41",	--719
		x"12",	--720
		x"42",	--721
		x"02",	--722
		x"93",	--723
		x"38",	--724
		x"92",	--725
		x"02",	--726
		x"24",	--727
		x"40",	--728
		x"02",	--729
		x"43",	--730
		x"3c",	--731
		x"52",	--732
		x"9f",	--733
		x"ff",	--734
		x"24",	--735
		x"53",	--736
		x"9b",	--737
		x"23",	--738
		x"12",	--739
		x"f7",	--740
		x"12",	--741
		x"e7",	--742
		x"53",	--743
		x"43",	--744
		x"41",	--745
		x"41",	--746
		x"43",	--747
		x"5c",	--748
		x"5c",	--749
		x"50",	--750
		x"02",	--751
		x"4e",	--752
		x"12",	--753
		x"00",	--754
		x"41",	--755
		x"41",	--756
		x"42",	--757
		x"00",	--758
		x"f2",	--759
		x"23",	--760
		x"4f",	--761
		x"00",	--762
		x"4f",	--763
		x"00",	--764
		x"43",	--765
		x"41",	--766
		x"f0",	--767
		x"00",	--768
		x"4f",	--769
		x"f8",	--770
		x"11",	--771
		x"12",	--772
		x"e5",	--773
		x"41",	--774
		x"12",	--775
		x"4f",	--776
		x"4f",	--777
		x"11",	--778
		x"11",	--779
		x"11",	--780
		x"11",	--781
		x"4e",	--782
		x"12",	--783
		x"e5",	--784
		x"4b",	--785
		x"12",	--786
		x"e5",	--787
		x"41",	--788
		x"41",	--789
		x"12",	--790
		x"12",	--791
		x"4f",	--792
		x"40",	--793
		x"00",	--794
		x"4a",	--795
		x"4b",	--796
		x"f0",	--797
		x"00",	--798
		x"24",	--799
		x"11",	--800
		x"53",	--801
		x"23",	--802
		x"f3",	--803
		x"24",	--804
		x"40",	--805
		x"00",	--806
		x"12",	--807
		x"e5",	--808
		x"53",	--809
		x"93",	--810
		x"23",	--811
		x"41",	--812
		x"41",	--813
		x"41",	--814
		x"40",	--815
		x"00",	--816
		x"3f",	--817
		x"12",	--818
		x"4f",	--819
		x"4f",	--820
		x"10",	--821
		x"11",	--822
		x"4e",	--823
		x"12",	--824
		x"e6",	--825
		x"4b",	--826
		x"12",	--827
		x"e6",	--828
		x"41",	--829
		x"41",	--830
		x"12",	--831
		x"12",	--832
		x"4e",	--833
		x"4f",	--834
		x"4f",	--835
		x"10",	--836
		x"11",	--837
		x"4d",	--838
		x"12",	--839
		x"e6",	--840
		x"4b",	--841
		x"12",	--842
		x"e6",	--843
		x"4b",	--844
		x"4a",	--845
		x"10",	--846
		x"10",	--847
		x"ec",	--848
		x"ec",	--849
		x"4d",	--850
		x"12",	--851
		x"e6",	--852
		x"4a",	--853
		x"12",	--854
		x"e6",	--855
		x"41",	--856
		x"41",	--857
		x"41",	--858
		x"12",	--859
		x"12",	--860
		x"12",	--861
		x"4f",	--862
		x"93",	--863
		x"24",	--864
		x"4e",	--865
		x"53",	--866
		x"43",	--867
		x"4a",	--868
		x"5b",	--869
		x"4d",	--870
		x"11",	--871
		x"12",	--872
		x"e6",	--873
		x"99",	--874
		x"24",	--875
		x"53",	--876
		x"b0",	--877
		x"00",	--878
		x"20",	--879
		x"40",	--880
		x"00",	--881
		x"12",	--882
		x"e5",	--883
		x"3f",	--884
		x"40",	--885
		x"00",	--886
		x"12",	--887
		x"e5",	--888
		x"3f",	--889
		x"41",	--890
		x"41",	--891
		x"41",	--892
		x"41",	--893
		x"12",	--894
		x"12",	--895
		x"12",	--896
		x"4f",	--897
		x"93",	--898
		x"24",	--899
		x"4e",	--900
		x"53",	--901
		x"43",	--902
		x"4a",	--903
		x"11",	--904
		x"12",	--905
		x"e5",	--906
		x"99",	--907
		x"24",	--908
		x"53",	--909
		x"b0",	--910
		x"00",	--911
		x"23",	--912
		x"40",	--913
		x"00",	--914
		x"12",	--915
		x"e5",	--916
		x"4a",	--917
		x"11",	--918
		x"12",	--919
		x"e5",	--920
		x"99",	--921
		x"23",	--922
		x"41",	--923
		x"41",	--924
		x"41",	--925
		x"41",	--926
		x"12",	--927
		x"12",	--928
		x"12",	--929
		x"50",	--930
		x"ff",	--931
		x"4f",	--932
		x"93",	--933
		x"38",	--934
		x"90",	--935
		x"00",	--936
		x"38",	--937
		x"43",	--938
		x"41",	--939
		x"59",	--940
		x"40",	--941
		x"00",	--942
		x"4b",	--943
		x"12",	--944
		x"f6",	--945
		x"50",	--946
		x"00",	--947
		x"4f",	--948
		x"00",	--949
		x"53",	--950
		x"40",	--951
		x"00",	--952
		x"4b",	--953
		x"12",	--954
		x"f6",	--955
		x"4f",	--956
		x"90",	--957
		x"00",	--958
		x"37",	--959
		x"49",	--960
		x"53",	--961
		x"51",	--962
		x"40",	--963
		x"00",	--964
		x"4b",	--965
		x"12",	--966
		x"f6",	--967
		x"50",	--968
		x"00",	--969
		x"4f",	--970
		x"00",	--971
		x"53",	--972
		x"41",	--973
		x"5a",	--974
		x"4f",	--975
		x"11",	--976
		x"12",	--977
		x"e5",	--978
		x"93",	--979
		x"23",	--980
		x"50",	--981
		x"00",	--982
		x"41",	--983
		x"41",	--984
		x"41",	--985
		x"41",	--986
		x"40",	--987
		x"00",	--988
		x"12",	--989
		x"e5",	--990
		x"e3",	--991
		x"53",	--992
		x"3f",	--993
		x"43",	--994
		x"43",	--995
		x"3f",	--996
		x"12",	--997
		x"12",	--998
		x"12",	--999
		x"41",	--1000
		x"52",	--1001
		x"4b",	--1002
		x"49",	--1003
		x"93",	--1004
		x"20",	--1005
		x"3c",	--1006
		x"11",	--1007
		x"12",	--1008
		x"e5",	--1009
		x"49",	--1010
		x"4a",	--1011
		x"53",	--1012
		x"4a",	--1013
		x"00",	--1014
		x"93",	--1015
		x"24",	--1016
		x"90",	--1017
		x"00",	--1018
		x"23",	--1019
		x"49",	--1020
		x"53",	--1021
		x"49",	--1022
		x"00",	--1023
		x"50",	--1024
		x"ff",	--1025
		x"90",	--1026
		x"00",	--1027
		x"2f",	--1028
		x"4f",	--1029
		x"5f",	--1030
		x"4f",	--1031
		x"f8",	--1032
		x"41",	--1033
		x"41",	--1034
		x"41",	--1035
		x"41",	--1036
		x"4b",	--1037
		x"52",	--1038
		x"4b",	--1039
		x"00",	--1040
		x"4b",	--1041
		x"12",	--1042
		x"e6",	--1043
		x"49",	--1044
		x"3f",	--1045
		x"4b",	--1046
		x"53",	--1047
		x"4b",	--1048
		x"12",	--1049
		x"e6",	--1050
		x"49",	--1051
		x"3f",	--1052
		x"4b",	--1053
		x"53",	--1054
		x"4f",	--1055
		x"49",	--1056
		x"93",	--1057
		x"27",	--1058
		x"53",	--1059
		x"11",	--1060
		x"12",	--1061
		x"e5",	--1062
		x"49",	--1063
		x"93",	--1064
		x"23",	--1065
		x"3f",	--1066
		x"4b",	--1067
		x"52",	--1068
		x"4b",	--1069
		x"00",	--1070
		x"4b",	--1071
		x"12",	--1072
		x"e6",	--1073
		x"49",	--1074
		x"3f",	--1075
		x"4b",	--1076
		x"53",	--1077
		x"4b",	--1078
		x"4e",	--1079
		x"10",	--1080
		x"11",	--1081
		x"10",	--1082
		x"11",	--1083
		x"12",	--1084
		x"e6",	--1085
		x"49",	--1086
		x"3f",	--1087
		x"4b",	--1088
		x"53",	--1089
		x"4b",	--1090
		x"12",	--1091
		x"e7",	--1092
		x"49",	--1093
		x"3f",	--1094
		x"4b",	--1095
		x"53",	--1096
		x"4b",	--1097
		x"12",	--1098
		x"e5",	--1099
		x"49",	--1100
		x"3f",	--1101
		x"4b",	--1102
		x"53",	--1103
		x"4b",	--1104
		x"12",	--1105
		x"e6",	--1106
		x"49",	--1107
		x"3f",	--1108
		x"4b",	--1109
		x"53",	--1110
		x"4b",	--1111
		x"12",	--1112
		x"e6",	--1113
		x"49",	--1114
		x"3f",	--1115
		x"40",	--1116
		x"00",	--1117
		x"12",	--1118
		x"e5",	--1119
		x"3f",	--1120
		x"12",	--1121
		x"12",	--1122
		x"42",	--1123
		x"02",	--1124
		x"42",	--1125
		x"00",	--1126
		x"03",	--1127
		x"42",	--1128
		x"02",	--1129
		x"90",	--1130
		x"00",	--1131
		x"34",	--1132
		x"53",	--1133
		x"02",	--1134
		x"42",	--1135
		x"02",	--1136
		x"42",	--1137
		x"02",	--1138
		x"9f",	--1139
		x"20",	--1140
		x"53",	--1141
		x"02",	--1142
		x"40",	--1143
		x"00",	--1144
		x"00",	--1145
		x"c0",	--1146
		x"00",	--1147
		x"00",	--1148
		x"41",	--1149
		x"41",	--1150
		x"c0",	--1151
		x"00",	--1152
		x"00",	--1153
		x"13",	--1154
		x"43",	--1155
		x"02",	--1156
		x"3f",	--1157
		x"40",	--1158
		x"00",	--1159
		x"00",	--1160
		x"40",	--1161
		x"00",	--1162
		x"00",	--1163
		x"41",	--1164
		x"42",	--1165
		x"02",	--1166
		x"42",	--1167
		x"02",	--1168
		x"9f",	--1169
		x"38",	--1170
		x"42",	--1171
		x"02",	--1172
		x"82",	--1173
		x"02",	--1174
		x"41",	--1175
		x"42",	--1176
		x"02",	--1177
		x"42",	--1178
		x"02",	--1179
		x"40",	--1180
		x"00",	--1181
		x"8d",	--1182
		x"8e",	--1183
		x"41",	--1184
		x"42",	--1185
		x"02",	--1186
		x"4f",	--1187
		x"03",	--1188
		x"42",	--1189
		x"02",	--1190
		x"42",	--1191
		x"02",	--1192
		x"9e",	--1193
		x"24",	--1194
		x"42",	--1195
		x"02",	--1196
		x"90",	--1197
		x"00",	--1198
		x"38",	--1199
		x"43",	--1200
		x"02",	--1201
		x"41",	--1202
		x"53",	--1203
		x"02",	--1204
		x"41",	--1205
		x"43",	--1206
		x"41",	--1207
		x"12",	--1208
		x"12",	--1209
		x"4e",	--1210
		x"4f",	--1211
		x"43",	--1212
		x"40",	--1213
		x"4f",	--1214
		x"12",	--1215
		x"f0",	--1216
		x"93",	--1217
		x"34",	--1218
		x"4a",	--1219
		x"4b",	--1220
		x"12",	--1221
		x"f0",	--1222
		x"41",	--1223
		x"41",	--1224
		x"41",	--1225
		x"43",	--1226
		x"40",	--1227
		x"4f",	--1228
		x"4a",	--1229
		x"4b",	--1230
		x"12",	--1231
		x"ec",	--1232
		x"12",	--1233
		x"f0",	--1234
		x"53",	--1235
		x"60",	--1236
		x"80",	--1237
		x"41",	--1238
		x"41",	--1239
		x"41",	--1240
		x"12",	--1241
		x"12",	--1242
		x"12",	--1243
		x"12",	--1244
		x"12",	--1245
		x"12",	--1246
		x"12",	--1247
		x"12",	--1248
		x"50",	--1249
		x"ff",	--1250
		x"4d",	--1251
		x"4f",	--1252
		x"93",	--1253
		x"28",	--1254
		x"4e",	--1255
		x"93",	--1256
		x"28",	--1257
		x"92",	--1258
		x"20",	--1259
		x"40",	--1260
		x"ec",	--1261
		x"92",	--1262
		x"24",	--1263
		x"93",	--1264
		x"24",	--1265
		x"93",	--1266
		x"24",	--1267
		x"4f",	--1268
		x"00",	--1269
		x"00",	--1270
		x"4e",	--1271
		x"00",	--1272
		x"4f",	--1273
		x"00",	--1274
		x"4f",	--1275
		x"00",	--1276
		x"4e",	--1277
		x"00",	--1278
		x"4e",	--1279
		x"00",	--1280
		x"41",	--1281
		x"8b",	--1282
		x"4c",	--1283
		x"93",	--1284
		x"38",	--1285
		x"90",	--1286
		x"00",	--1287
		x"34",	--1288
		x"93",	--1289
		x"38",	--1290
		x"46",	--1291
		x"00",	--1292
		x"47",	--1293
		x"00",	--1294
		x"49",	--1295
		x"f0",	--1296
		x"00",	--1297
		x"24",	--1298
		x"46",	--1299
		x"47",	--1300
		x"c3",	--1301
		x"10",	--1302
		x"10",	--1303
		x"53",	--1304
		x"23",	--1305
		x"4a",	--1306
		x"00",	--1307
		x"4b",	--1308
		x"00",	--1309
		x"43",	--1310
		x"43",	--1311
		x"f0",	--1312
		x"00",	--1313
		x"24",	--1314
		x"5c",	--1315
		x"6d",	--1316
		x"53",	--1317
		x"23",	--1318
		x"53",	--1319
		x"63",	--1320
		x"f6",	--1321
		x"f7",	--1322
		x"43",	--1323
		x"43",	--1324
		x"93",	--1325
		x"20",	--1326
		x"93",	--1327
		x"24",	--1328
		x"41",	--1329
		x"00",	--1330
		x"41",	--1331
		x"00",	--1332
		x"da",	--1333
		x"db",	--1334
		x"4f",	--1335
		x"00",	--1336
		x"9e",	--1337
		x"00",	--1338
		x"20",	--1339
		x"4f",	--1340
		x"00",	--1341
		x"41",	--1342
		x"00",	--1343
		x"46",	--1344
		x"47",	--1345
		x"54",	--1346
		x"65",	--1347
		x"4e",	--1348
		x"00",	--1349
		x"4f",	--1350
		x"00",	--1351
		x"40",	--1352
		x"00",	--1353
		x"00",	--1354
		x"93",	--1355
		x"38",	--1356
		x"48",	--1357
		x"50",	--1358
		x"00",	--1359
		x"41",	--1360
		x"41",	--1361
		x"41",	--1362
		x"41",	--1363
		x"41",	--1364
		x"41",	--1365
		x"41",	--1366
		x"41",	--1367
		x"41",	--1368
		x"91",	--1369
		x"38",	--1370
		x"4b",	--1371
		x"00",	--1372
		x"43",	--1373
		x"43",	--1374
		x"4f",	--1375
		x"00",	--1376
		x"9e",	--1377
		x"00",	--1378
		x"27",	--1379
		x"93",	--1380
		x"24",	--1381
		x"46",	--1382
		x"47",	--1383
		x"84",	--1384
		x"75",	--1385
		x"93",	--1386
		x"38",	--1387
		x"43",	--1388
		x"00",	--1389
		x"41",	--1390
		x"00",	--1391
		x"4e",	--1392
		x"00",	--1393
		x"4f",	--1394
		x"00",	--1395
		x"4e",	--1396
		x"4f",	--1397
		x"53",	--1398
		x"63",	--1399
		x"90",	--1400
		x"3f",	--1401
		x"28",	--1402
		x"90",	--1403
		x"40",	--1404
		x"2c",	--1405
		x"93",	--1406
		x"2c",	--1407
		x"48",	--1408
		x"00",	--1409
		x"53",	--1410
		x"5e",	--1411
		x"6f",	--1412
		x"4b",	--1413
		x"53",	--1414
		x"4e",	--1415
		x"4f",	--1416
		x"53",	--1417
		x"63",	--1418
		x"90",	--1419
		x"3f",	--1420
		x"2b",	--1421
		x"24",	--1422
		x"4e",	--1423
		x"00",	--1424
		x"4f",	--1425
		x"00",	--1426
		x"4a",	--1427
		x"00",	--1428
		x"40",	--1429
		x"00",	--1430
		x"00",	--1431
		x"93",	--1432
		x"37",	--1433
		x"4e",	--1434
		x"4f",	--1435
		x"f3",	--1436
		x"f3",	--1437
		x"c3",	--1438
		x"10",	--1439
		x"10",	--1440
		x"4c",	--1441
		x"4d",	--1442
		x"de",	--1443
		x"df",	--1444
		x"4a",	--1445
		x"00",	--1446
		x"4b",	--1447
		x"00",	--1448
		x"53",	--1449
		x"00",	--1450
		x"48",	--1451
		x"3f",	--1452
		x"93",	--1453
		x"23",	--1454
		x"4f",	--1455
		x"00",	--1456
		x"4f",	--1457
		x"00",	--1458
		x"00",	--1459
		x"4f",	--1460
		x"00",	--1461
		x"00",	--1462
		x"4f",	--1463
		x"00",	--1464
		x"00",	--1465
		x"4e",	--1466
		x"00",	--1467
		x"ff",	--1468
		x"00",	--1469
		x"4e",	--1470
		x"00",	--1471
		x"4d",	--1472
		x"3f",	--1473
		x"43",	--1474
		x"43",	--1475
		x"3f",	--1476
		x"e3",	--1477
		x"53",	--1478
		x"90",	--1479
		x"00",	--1480
		x"37",	--1481
		x"3f",	--1482
		x"93",	--1483
		x"2b",	--1484
		x"3f",	--1485
		x"44",	--1486
		x"45",	--1487
		x"86",	--1488
		x"77",	--1489
		x"3f",	--1490
		x"4e",	--1491
		x"3f",	--1492
		x"43",	--1493
		x"00",	--1494
		x"41",	--1495
		x"00",	--1496
		x"e3",	--1497
		x"e3",	--1498
		x"53",	--1499
		x"63",	--1500
		x"4e",	--1501
		x"00",	--1502
		x"4f",	--1503
		x"00",	--1504
		x"3f",	--1505
		x"93",	--1506
		x"27",	--1507
		x"59",	--1508
		x"00",	--1509
		x"44",	--1510
		x"00",	--1511
		x"45",	--1512
		x"00",	--1513
		x"49",	--1514
		x"f0",	--1515
		x"00",	--1516
		x"24",	--1517
		x"4d",	--1518
		x"44",	--1519
		x"45",	--1520
		x"c3",	--1521
		x"10",	--1522
		x"10",	--1523
		x"53",	--1524
		x"23",	--1525
		x"4c",	--1526
		x"00",	--1527
		x"4d",	--1528
		x"00",	--1529
		x"43",	--1530
		x"43",	--1531
		x"f0",	--1532
		x"00",	--1533
		x"24",	--1534
		x"5c",	--1535
		x"6d",	--1536
		x"53",	--1537
		x"23",	--1538
		x"53",	--1539
		x"63",	--1540
		x"f4",	--1541
		x"f5",	--1542
		x"43",	--1543
		x"43",	--1544
		x"93",	--1545
		x"20",	--1546
		x"93",	--1547
		x"20",	--1548
		x"43",	--1549
		x"43",	--1550
		x"41",	--1551
		x"00",	--1552
		x"41",	--1553
		x"00",	--1554
		x"da",	--1555
		x"db",	--1556
		x"3f",	--1557
		x"43",	--1558
		x"43",	--1559
		x"3f",	--1560
		x"92",	--1561
		x"23",	--1562
		x"9e",	--1563
		x"00",	--1564
		x"00",	--1565
		x"27",	--1566
		x"40",	--1567
		x"f8",	--1568
		x"3f",	--1569
		x"50",	--1570
		x"ff",	--1571
		x"4e",	--1572
		x"00",	--1573
		x"4f",	--1574
		x"00",	--1575
		x"4c",	--1576
		x"00",	--1577
		x"4d",	--1578
		x"00",	--1579
		x"41",	--1580
		x"50",	--1581
		x"00",	--1582
		x"41",	--1583
		x"52",	--1584
		x"12",	--1585
		x"f4",	--1586
		x"41",	--1587
		x"50",	--1588
		x"00",	--1589
		x"41",	--1590
		x"12",	--1591
		x"f4",	--1592
		x"41",	--1593
		x"52",	--1594
		x"41",	--1595
		x"50",	--1596
		x"00",	--1597
		x"41",	--1598
		x"50",	--1599
		x"00",	--1600
		x"12",	--1601
		x"e9",	--1602
		x"12",	--1603
		x"f2",	--1604
		x"50",	--1605
		x"00",	--1606
		x"41",	--1607
		x"50",	--1608
		x"ff",	--1609
		x"4e",	--1610
		x"00",	--1611
		x"4f",	--1612
		x"00",	--1613
		x"4c",	--1614
		x"00",	--1615
		x"4d",	--1616
		x"00",	--1617
		x"41",	--1618
		x"50",	--1619
		x"00",	--1620
		x"41",	--1621
		x"52",	--1622
		x"12",	--1623
		x"f4",	--1624
		x"41",	--1625
		x"50",	--1626
		x"00",	--1627
		x"41",	--1628
		x"12",	--1629
		x"f4",	--1630
		x"e3",	--1631
		x"00",	--1632
		x"41",	--1633
		x"52",	--1634
		x"41",	--1635
		x"50",	--1636
		x"00",	--1637
		x"41",	--1638
		x"50",	--1639
		x"00",	--1640
		x"12",	--1641
		x"e9",	--1642
		x"12",	--1643
		x"f2",	--1644
		x"50",	--1645
		x"00",	--1646
		x"41",	--1647
		x"12",	--1648
		x"12",	--1649
		x"12",	--1650
		x"12",	--1651
		x"12",	--1652
		x"12",	--1653
		x"12",	--1654
		x"12",	--1655
		x"50",	--1656
		x"ff",	--1657
		x"4e",	--1658
		x"00",	--1659
		x"4f",	--1660
		x"00",	--1661
		x"4c",	--1662
		x"00",	--1663
		x"4d",	--1664
		x"00",	--1665
		x"41",	--1666
		x"50",	--1667
		x"00",	--1668
		x"41",	--1669
		x"52",	--1670
		x"12",	--1671
		x"f4",	--1672
		x"41",	--1673
		x"50",	--1674
		x"00",	--1675
		x"41",	--1676
		x"12",	--1677
		x"f4",	--1678
		x"41",	--1679
		x"00",	--1680
		x"93",	--1681
		x"28",	--1682
		x"41",	--1683
		x"00",	--1684
		x"93",	--1685
		x"28",	--1686
		x"92",	--1687
		x"24",	--1688
		x"92",	--1689
		x"24",	--1690
		x"93",	--1691
		x"24",	--1692
		x"93",	--1693
		x"24",	--1694
		x"41",	--1695
		x"00",	--1696
		x"41",	--1697
		x"00",	--1698
		x"41",	--1699
		x"00",	--1700
		x"41",	--1701
		x"00",	--1702
		x"40",	--1703
		x"00",	--1704
		x"43",	--1705
		x"43",	--1706
		x"43",	--1707
		x"43",	--1708
		x"43",	--1709
		x"00",	--1710
		x"43",	--1711
		x"00",	--1712
		x"43",	--1713
		x"43",	--1714
		x"4c",	--1715
		x"00",	--1716
		x"3c",	--1717
		x"58",	--1718
		x"69",	--1719
		x"c3",	--1720
		x"10",	--1721
		x"10",	--1722
		x"53",	--1723
		x"00",	--1724
		x"24",	--1725
		x"b3",	--1726
		x"24",	--1727
		x"58",	--1728
		x"69",	--1729
		x"56",	--1730
		x"67",	--1731
		x"43",	--1732
		x"43",	--1733
		x"99",	--1734
		x"28",	--1735
		x"24",	--1736
		x"43",	--1737
		x"43",	--1738
		x"5c",	--1739
		x"6d",	--1740
		x"56",	--1741
		x"67",	--1742
		x"93",	--1743
		x"37",	--1744
		x"d3",	--1745
		x"d3",	--1746
		x"3f",	--1747
		x"98",	--1748
		x"2b",	--1749
		x"3f",	--1750
		x"4a",	--1751
		x"00",	--1752
		x"4b",	--1753
		x"00",	--1754
		x"4f",	--1755
		x"41",	--1756
		x"00",	--1757
		x"51",	--1758
		x"00",	--1759
		x"4a",	--1760
		x"53",	--1761
		x"46",	--1762
		x"00",	--1763
		x"43",	--1764
		x"91",	--1765
		x"00",	--1766
		x"00",	--1767
		x"24",	--1768
		x"4d",	--1769
		x"00",	--1770
		x"93",	--1771
		x"38",	--1772
		x"90",	--1773
		x"40",	--1774
		x"2c",	--1775
		x"41",	--1776
		x"00",	--1777
		x"53",	--1778
		x"41",	--1779
		x"00",	--1780
		x"41",	--1781
		x"00",	--1782
		x"4d",	--1783
		x"5e",	--1784
		x"6f",	--1785
		x"93",	--1786
		x"38",	--1787
		x"5a",	--1788
		x"6b",	--1789
		x"53",	--1790
		x"90",	--1791
		x"40",	--1792
		x"2b",	--1793
		x"4a",	--1794
		x"00",	--1795
		x"4b",	--1796
		x"00",	--1797
		x"4c",	--1798
		x"00",	--1799
		x"4e",	--1800
		x"4f",	--1801
		x"f0",	--1802
		x"00",	--1803
		x"f3",	--1804
		x"90",	--1805
		x"00",	--1806
		x"24",	--1807
		x"4e",	--1808
		x"00",	--1809
		x"4f",	--1810
		x"00",	--1811
		x"40",	--1812
		x"00",	--1813
		x"00",	--1814
		x"41",	--1815
		x"52",	--1816
		x"12",	--1817
		x"f2",	--1818
		x"50",	--1819
		x"00",	--1820
		x"41",	--1821
		x"41",	--1822
		x"41",	--1823
		x"41",	--1824
		x"41",	--1825
		x"41",	--1826
		x"41",	--1827
		x"41",	--1828
		x"41",	--1829
		x"d3",	--1830
		x"d3",	--1831
		x"3f",	--1832
		x"50",	--1833
		x"00",	--1834
		x"4a",	--1835
		x"b3",	--1836
		x"24",	--1837
		x"41",	--1838
		x"00",	--1839
		x"41",	--1840
		x"00",	--1841
		x"c3",	--1842
		x"10",	--1843
		x"10",	--1844
		x"4c",	--1845
		x"4d",	--1846
		x"d3",	--1847
		x"d0",	--1848
		x"80",	--1849
		x"46",	--1850
		x"00",	--1851
		x"47",	--1852
		x"00",	--1853
		x"c3",	--1854
		x"10",	--1855
		x"10",	--1856
		x"53",	--1857
		x"93",	--1858
		x"3b",	--1859
		x"48",	--1860
		x"00",	--1861
		x"3f",	--1862
		x"93",	--1863
		x"24",	--1864
		x"43",	--1865
		x"91",	--1866
		x"00",	--1867
		x"00",	--1868
		x"24",	--1869
		x"4f",	--1870
		x"00",	--1871
		x"41",	--1872
		x"50",	--1873
		x"00",	--1874
		x"3f",	--1875
		x"93",	--1876
		x"23",	--1877
		x"4e",	--1878
		x"4f",	--1879
		x"f0",	--1880
		x"00",	--1881
		x"f3",	--1882
		x"93",	--1883
		x"23",	--1884
		x"93",	--1885
		x"23",	--1886
		x"93",	--1887
		x"00",	--1888
		x"20",	--1889
		x"93",	--1890
		x"00",	--1891
		x"27",	--1892
		x"50",	--1893
		x"00",	--1894
		x"63",	--1895
		x"f0",	--1896
		x"ff",	--1897
		x"f3",	--1898
		x"3f",	--1899
		x"43",	--1900
		x"3f",	--1901
		x"43",	--1902
		x"3f",	--1903
		x"43",	--1904
		x"91",	--1905
		x"00",	--1906
		x"00",	--1907
		x"24",	--1908
		x"4f",	--1909
		x"00",	--1910
		x"41",	--1911
		x"50",	--1912
		x"00",	--1913
		x"3f",	--1914
		x"43",	--1915
		x"3f",	--1916
		x"93",	--1917
		x"23",	--1918
		x"40",	--1919
		x"f8",	--1920
		x"3f",	--1921
		x"12",	--1922
		x"12",	--1923
		x"12",	--1924
		x"12",	--1925
		x"12",	--1926
		x"50",	--1927
		x"ff",	--1928
		x"4e",	--1929
		x"00",	--1930
		x"4f",	--1931
		x"00",	--1932
		x"4c",	--1933
		x"00",	--1934
		x"4d",	--1935
		x"00",	--1936
		x"41",	--1937
		x"50",	--1938
		x"00",	--1939
		x"41",	--1940
		x"52",	--1941
		x"12",	--1942
		x"f4",	--1943
		x"41",	--1944
		x"52",	--1945
		x"41",	--1946
		x"12",	--1947
		x"f4",	--1948
		x"41",	--1949
		x"00",	--1950
		x"93",	--1951
		x"28",	--1952
		x"41",	--1953
		x"00",	--1954
		x"93",	--1955
		x"28",	--1956
		x"e1",	--1957
		x"00",	--1958
		x"00",	--1959
		x"92",	--1960
		x"24",	--1961
		x"93",	--1962
		x"24",	--1963
		x"92",	--1964
		x"24",	--1965
		x"93",	--1966
		x"24",	--1967
		x"41",	--1968
		x"00",	--1969
		x"81",	--1970
		x"00",	--1971
		x"4d",	--1972
		x"00",	--1973
		x"41",	--1974
		x"00",	--1975
		x"41",	--1976
		x"00",	--1977
		x"41",	--1978
		x"00",	--1979
		x"41",	--1980
		x"00",	--1981
		x"99",	--1982
		x"2c",	--1983
		x"5e",	--1984
		x"6f",	--1985
		x"53",	--1986
		x"4d",	--1987
		x"00",	--1988
		x"40",	--1989
		x"00",	--1990
		x"43",	--1991
		x"40",	--1992
		x"40",	--1993
		x"43",	--1994
		x"43",	--1995
		x"3c",	--1996
		x"dc",	--1997
		x"dd",	--1998
		x"88",	--1999
		x"79",	--2000
		x"c3",	--2001
		x"10",	--2002
		x"10",	--2003
		x"5e",	--2004
		x"6f",	--2005
		x"53",	--2006
		x"24",	--2007
		x"99",	--2008
		x"2b",	--2009
		x"23",	--2010
		x"98",	--2011
		x"2b",	--2012
		x"3f",	--2013
		x"9f",	--2014
		x"2b",	--2015
		x"98",	--2016
		x"2f",	--2017
		x"3f",	--2018
		x"4a",	--2019
		x"4b",	--2020
		x"f0",	--2021
		x"00",	--2022
		x"f3",	--2023
		x"90",	--2024
		x"00",	--2025
		x"24",	--2026
		x"4a",	--2027
		x"00",	--2028
		x"4b",	--2029
		x"00",	--2030
		x"41",	--2031
		x"50",	--2032
		x"00",	--2033
		x"12",	--2034
		x"f2",	--2035
		x"50",	--2036
		x"00",	--2037
		x"41",	--2038
		x"41",	--2039
		x"41",	--2040
		x"41",	--2041
		x"41",	--2042
		x"41",	--2043
		x"42",	--2044
		x"00",	--2045
		x"41",	--2046
		x"50",	--2047
		x"00",	--2048
		x"3f",	--2049
		x"9e",	--2050
		x"23",	--2051
		x"40",	--2052
		x"f8",	--2053
		x"3f",	--2054
		x"93",	--2055
		x"23",	--2056
		x"4a",	--2057
		x"4b",	--2058
		x"f0",	--2059
		x"00",	--2060
		x"f3",	--2061
		x"93",	--2062
		x"23",	--2063
		x"93",	--2064
		x"23",	--2065
		x"93",	--2066
		x"20",	--2067
		x"93",	--2068
		x"27",	--2069
		x"50",	--2070
		x"00",	--2071
		x"63",	--2072
		x"f0",	--2073
		x"ff",	--2074
		x"f3",	--2075
		x"3f",	--2076
		x"43",	--2077
		x"00",	--2078
		x"43",	--2079
		x"00",	--2080
		x"43",	--2081
		x"00",	--2082
		x"41",	--2083
		x"50",	--2084
		x"00",	--2085
		x"3f",	--2086
		x"41",	--2087
		x"52",	--2088
		x"3f",	--2089
		x"50",	--2090
		x"ff",	--2091
		x"4e",	--2092
		x"00",	--2093
		x"4f",	--2094
		x"00",	--2095
		x"4c",	--2096
		x"00",	--2097
		x"4d",	--2098
		x"00",	--2099
		x"41",	--2100
		x"50",	--2101
		x"00",	--2102
		x"41",	--2103
		x"52",	--2104
		x"12",	--2105
		x"f4",	--2106
		x"41",	--2107
		x"52",	--2108
		x"41",	--2109
		x"12",	--2110
		x"f4",	--2111
		x"93",	--2112
		x"00",	--2113
		x"28",	--2114
		x"93",	--2115
		x"00",	--2116
		x"28",	--2117
		x"41",	--2118
		x"52",	--2119
		x"41",	--2120
		x"50",	--2121
		x"00",	--2122
		x"12",	--2123
		x"f5",	--2124
		x"50",	--2125
		x"00",	--2126
		x"41",	--2127
		x"43",	--2128
		x"3f",	--2129
		x"50",	--2130
		x"ff",	--2131
		x"4e",	--2132
		x"00",	--2133
		x"4f",	--2134
		x"00",	--2135
		x"41",	--2136
		x"52",	--2137
		x"41",	--2138
		x"12",	--2139
		x"f4",	--2140
		x"41",	--2141
		x"00",	--2142
		x"93",	--2143
		x"24",	--2144
		x"28",	--2145
		x"92",	--2146
		x"24",	--2147
		x"41",	--2148
		x"00",	--2149
		x"93",	--2150
		x"38",	--2151
		x"90",	--2152
		x"00",	--2153
		x"38",	--2154
		x"93",	--2155
		x"00",	--2156
		x"20",	--2157
		x"43",	--2158
		x"40",	--2159
		x"7f",	--2160
		x"50",	--2161
		x"00",	--2162
		x"41",	--2163
		x"41",	--2164
		x"00",	--2165
		x"41",	--2166
		x"00",	--2167
		x"40",	--2168
		x"00",	--2169
		x"8d",	--2170
		x"4c",	--2171
		x"f0",	--2172
		x"00",	--2173
		x"20",	--2174
		x"93",	--2175
		x"00",	--2176
		x"27",	--2177
		x"e3",	--2178
		x"e3",	--2179
		x"53",	--2180
		x"63",	--2181
		x"50",	--2182
		x"00",	--2183
		x"41",	--2184
		x"43",	--2185
		x"43",	--2186
		x"50",	--2187
		x"00",	--2188
		x"41",	--2189
		x"c3",	--2190
		x"10",	--2191
		x"10",	--2192
		x"53",	--2193
		x"23",	--2194
		x"3f",	--2195
		x"43",	--2196
		x"40",	--2197
		x"80",	--2198
		x"50",	--2199
		x"00",	--2200
		x"41",	--2201
		x"12",	--2202
		x"12",	--2203
		x"12",	--2204
		x"12",	--2205
		x"82",	--2206
		x"4e",	--2207
		x"4f",	--2208
		x"43",	--2209
		x"00",	--2210
		x"93",	--2211
		x"20",	--2212
		x"93",	--2213
		x"20",	--2214
		x"43",	--2215
		x"00",	--2216
		x"41",	--2217
		x"12",	--2218
		x"f2",	--2219
		x"52",	--2220
		x"41",	--2221
		x"41",	--2222
		x"41",	--2223
		x"41",	--2224
		x"41",	--2225
		x"40",	--2226
		x"00",	--2227
		x"00",	--2228
		x"40",	--2229
		x"00",	--2230
		x"00",	--2231
		x"4a",	--2232
		x"00",	--2233
		x"4b",	--2234
		x"00",	--2235
		x"4a",	--2236
		x"4b",	--2237
		x"12",	--2238
		x"f2",	--2239
		x"53",	--2240
		x"93",	--2241
		x"38",	--2242
		x"27",	--2243
		x"4a",	--2244
		x"00",	--2245
		x"4b",	--2246
		x"00",	--2247
		x"4f",	--2248
		x"f0",	--2249
		x"00",	--2250
		x"20",	--2251
		x"40",	--2252
		x"00",	--2253
		x"8f",	--2254
		x"4e",	--2255
		x"00",	--2256
		x"3f",	--2257
		x"51",	--2258
		x"00",	--2259
		x"00",	--2260
		x"61",	--2261
		x"00",	--2262
		x"00",	--2263
		x"53",	--2264
		x"23",	--2265
		x"3f",	--2266
		x"4f",	--2267
		x"e3",	--2268
		x"53",	--2269
		x"43",	--2270
		x"43",	--2271
		x"4e",	--2272
		x"f0",	--2273
		x"00",	--2274
		x"24",	--2275
		x"5c",	--2276
		x"6d",	--2277
		x"53",	--2278
		x"23",	--2279
		x"53",	--2280
		x"63",	--2281
		x"fa",	--2282
		x"fb",	--2283
		x"43",	--2284
		x"43",	--2285
		x"93",	--2286
		x"20",	--2287
		x"93",	--2288
		x"20",	--2289
		x"43",	--2290
		x"43",	--2291
		x"f0",	--2292
		x"00",	--2293
		x"20",	--2294
		x"48",	--2295
		x"49",	--2296
		x"da",	--2297
		x"db",	--2298
		x"4d",	--2299
		x"00",	--2300
		x"4e",	--2301
		x"00",	--2302
		x"40",	--2303
		x"00",	--2304
		x"8f",	--2305
		x"4e",	--2306
		x"00",	--2307
		x"3f",	--2308
		x"c3",	--2309
		x"10",	--2310
		x"10",	--2311
		x"53",	--2312
		x"23",	--2313
		x"3f",	--2314
		x"12",	--2315
		x"12",	--2316
		x"12",	--2317
		x"93",	--2318
		x"2c",	--2319
		x"90",	--2320
		x"01",	--2321
		x"28",	--2322
		x"40",	--2323
		x"00",	--2324
		x"43",	--2325
		x"42",	--2326
		x"4e",	--2327
		x"4f",	--2328
		x"49",	--2329
		x"93",	--2330
		x"20",	--2331
		x"50",	--2332
		x"f8",	--2333
		x"4c",	--2334
		x"43",	--2335
		x"8e",	--2336
		x"7f",	--2337
		x"4a",	--2338
		x"41",	--2339
		x"41",	--2340
		x"41",	--2341
		x"41",	--2342
		x"90",	--2343
		x"01",	--2344
		x"28",	--2345
		x"42",	--2346
		x"43",	--2347
		x"40",	--2348
		x"00",	--2349
		x"4e",	--2350
		x"4f",	--2351
		x"49",	--2352
		x"93",	--2353
		x"27",	--2354
		x"c3",	--2355
		x"10",	--2356
		x"10",	--2357
		x"53",	--2358
		x"23",	--2359
		x"3f",	--2360
		x"40",	--2361
		x"00",	--2362
		x"43",	--2363
		x"40",	--2364
		x"00",	--2365
		x"3f",	--2366
		x"40",	--2367
		x"00",	--2368
		x"43",	--2369
		x"43",	--2370
		x"3f",	--2371
		x"12",	--2372
		x"12",	--2373
		x"12",	--2374
		x"12",	--2375
		x"12",	--2376
		x"4f",	--2377
		x"4f",	--2378
		x"00",	--2379
		x"4f",	--2380
		x"00",	--2381
		x"4d",	--2382
		x"00",	--2383
		x"4d",	--2384
		x"93",	--2385
		x"28",	--2386
		x"92",	--2387
		x"24",	--2388
		x"93",	--2389
		x"24",	--2390
		x"93",	--2391
		x"24",	--2392
		x"4d",	--2393
		x"00",	--2394
		x"90",	--2395
		x"ff",	--2396
		x"38",	--2397
		x"90",	--2398
		x"00",	--2399
		x"34",	--2400
		x"4e",	--2401
		x"4f",	--2402
		x"f0",	--2403
		x"00",	--2404
		x"f3",	--2405
		x"90",	--2406
		x"00",	--2407
		x"24",	--2408
		x"50",	--2409
		x"00",	--2410
		x"63",	--2411
		x"93",	--2412
		x"38",	--2413
		x"4b",	--2414
		x"50",	--2415
		x"00",	--2416
		x"c3",	--2417
		x"10",	--2418
		x"10",	--2419
		x"c3",	--2420
		x"10",	--2421
		x"10",	--2422
		x"c3",	--2423
		x"10",	--2424
		x"10",	--2425
		x"c3",	--2426
		x"10",	--2427
		x"10",	--2428
		x"c3",	--2429
		x"10",	--2430
		x"10",	--2431
		x"c3",	--2432
		x"10",	--2433
		x"10",	--2434
		x"c3",	--2435
		x"10",	--2436
		x"10",	--2437
		x"f3",	--2438
		x"f0",	--2439
		x"00",	--2440
		x"4d",	--2441
		x"3c",	--2442
		x"93",	--2443
		x"23",	--2444
		x"43",	--2445
		x"43",	--2446
		x"43",	--2447
		x"4d",	--2448
		x"5d",	--2449
		x"5d",	--2450
		x"5d",	--2451
		x"5d",	--2452
		x"5d",	--2453
		x"5d",	--2454
		x"5d",	--2455
		x"4f",	--2456
		x"f0",	--2457
		x"00",	--2458
		x"dd",	--2459
		x"4a",	--2460
		x"11",	--2461
		x"43",	--2462
		x"10",	--2463
		x"4c",	--2464
		x"df",	--2465
		x"4d",	--2466
		x"41",	--2467
		x"41",	--2468
		x"41",	--2469
		x"41",	--2470
		x"41",	--2471
		x"41",	--2472
		x"93",	--2473
		x"23",	--2474
		x"4e",	--2475
		x"4f",	--2476
		x"f0",	--2477
		x"00",	--2478
		x"f3",	--2479
		x"93",	--2480
		x"20",	--2481
		x"93",	--2482
		x"27",	--2483
		x"50",	--2484
		x"00",	--2485
		x"63",	--2486
		x"3f",	--2487
		x"c3",	--2488
		x"10",	--2489
		x"10",	--2490
		x"4b",	--2491
		x"50",	--2492
		x"00",	--2493
		x"3f",	--2494
		x"43",	--2495
		x"43",	--2496
		x"43",	--2497
		x"3f",	--2498
		x"d3",	--2499
		x"d0",	--2500
		x"00",	--2501
		x"f3",	--2502
		x"f0",	--2503
		x"00",	--2504
		x"43",	--2505
		x"3f",	--2506
		x"40",	--2507
		x"ff",	--2508
		x"8b",	--2509
		x"90",	--2510
		x"00",	--2511
		x"34",	--2512
		x"4e",	--2513
		x"4f",	--2514
		x"47",	--2515
		x"f0",	--2516
		x"00",	--2517
		x"24",	--2518
		x"c3",	--2519
		x"10",	--2520
		x"10",	--2521
		x"53",	--2522
		x"23",	--2523
		x"43",	--2524
		x"43",	--2525
		x"f0",	--2526
		x"00",	--2527
		x"24",	--2528
		x"58",	--2529
		x"69",	--2530
		x"53",	--2531
		x"23",	--2532
		x"53",	--2533
		x"63",	--2534
		x"fe",	--2535
		x"ff",	--2536
		x"43",	--2537
		x"43",	--2538
		x"93",	--2539
		x"20",	--2540
		x"93",	--2541
		x"20",	--2542
		x"43",	--2543
		x"43",	--2544
		x"4e",	--2545
		x"4f",	--2546
		x"dc",	--2547
		x"dd",	--2548
		x"48",	--2549
		x"49",	--2550
		x"f0",	--2551
		x"00",	--2552
		x"f3",	--2553
		x"90",	--2554
		x"00",	--2555
		x"24",	--2556
		x"50",	--2557
		x"00",	--2558
		x"63",	--2559
		x"48",	--2560
		x"49",	--2561
		x"c3",	--2562
		x"10",	--2563
		x"10",	--2564
		x"c3",	--2565
		x"10",	--2566
		x"10",	--2567
		x"c3",	--2568
		x"10",	--2569
		x"10",	--2570
		x"c3",	--2571
		x"10",	--2572
		x"10",	--2573
		x"c3",	--2574
		x"10",	--2575
		x"10",	--2576
		x"c3",	--2577
		x"10",	--2578
		x"10",	--2579
		x"c3",	--2580
		x"10",	--2581
		x"10",	--2582
		x"f3",	--2583
		x"f0",	--2584
		x"00",	--2585
		x"43",	--2586
		x"90",	--2587
		x"40",	--2588
		x"2f",	--2589
		x"43",	--2590
		x"3f",	--2591
		x"43",	--2592
		x"43",	--2593
		x"3f",	--2594
		x"93",	--2595
		x"23",	--2596
		x"48",	--2597
		x"49",	--2598
		x"f0",	--2599
		x"00",	--2600
		x"f3",	--2601
		x"93",	--2602
		x"24",	--2603
		x"50",	--2604
		x"00",	--2605
		x"63",	--2606
		x"3f",	--2607
		x"93",	--2608
		x"27",	--2609
		x"3f",	--2610
		x"12",	--2611
		x"12",	--2612
		x"4f",	--2613
		x"4f",	--2614
		x"00",	--2615
		x"f0",	--2616
		x"00",	--2617
		x"4f",	--2618
		x"00",	--2619
		x"c3",	--2620
		x"10",	--2621
		x"c3",	--2622
		x"10",	--2623
		x"c3",	--2624
		x"10",	--2625
		x"c3",	--2626
		x"10",	--2627
		x"c3",	--2628
		x"10",	--2629
		x"c3",	--2630
		x"10",	--2631
		x"c3",	--2632
		x"10",	--2633
		x"4d",	--2634
		x"4f",	--2635
		x"00",	--2636
		x"b0",	--2637
		x"00",	--2638
		x"43",	--2639
		x"6f",	--2640
		x"4f",	--2641
		x"00",	--2642
		x"93",	--2643
		x"20",	--2644
		x"93",	--2645
		x"24",	--2646
		x"40",	--2647
		x"ff",	--2648
		x"00",	--2649
		x"4a",	--2650
		x"4b",	--2651
		x"5c",	--2652
		x"6d",	--2653
		x"5c",	--2654
		x"6d",	--2655
		x"5c",	--2656
		x"6d",	--2657
		x"5c",	--2658
		x"6d",	--2659
		x"5c",	--2660
		x"6d",	--2661
		x"5c",	--2662
		x"6d",	--2663
		x"5c",	--2664
		x"6d",	--2665
		x"40",	--2666
		x"00",	--2667
		x"00",	--2668
		x"90",	--2669
		x"40",	--2670
		x"2c",	--2671
		x"40",	--2672
		x"ff",	--2673
		x"5c",	--2674
		x"6d",	--2675
		x"4f",	--2676
		x"53",	--2677
		x"90",	--2678
		x"40",	--2679
		x"2b",	--2680
		x"4a",	--2681
		x"00",	--2682
		x"4c",	--2683
		x"00",	--2684
		x"4d",	--2685
		x"00",	--2686
		x"41",	--2687
		x"41",	--2688
		x"41",	--2689
		x"90",	--2690
		x"00",	--2691
		x"24",	--2692
		x"50",	--2693
		x"ff",	--2694
		x"4d",	--2695
		x"00",	--2696
		x"40",	--2697
		x"00",	--2698
		x"00",	--2699
		x"4a",	--2700
		x"4b",	--2701
		x"5c",	--2702
		x"6d",	--2703
		x"5c",	--2704
		x"6d",	--2705
		x"5c",	--2706
		x"6d",	--2707
		x"5c",	--2708
		x"6d",	--2709
		x"5c",	--2710
		x"6d",	--2711
		x"5c",	--2712
		x"6d",	--2713
		x"5c",	--2714
		x"6d",	--2715
		x"4c",	--2716
		x"4d",	--2717
		x"d3",	--2718
		x"d0",	--2719
		x"40",	--2720
		x"4a",	--2721
		x"00",	--2722
		x"4b",	--2723
		x"00",	--2724
		x"41",	--2725
		x"41",	--2726
		x"41",	--2727
		x"93",	--2728
		x"23",	--2729
		x"43",	--2730
		x"00",	--2731
		x"41",	--2732
		x"41",	--2733
		x"41",	--2734
		x"93",	--2735
		x"24",	--2736
		x"4a",	--2737
		x"4b",	--2738
		x"f3",	--2739
		x"f0",	--2740
		x"00",	--2741
		x"93",	--2742
		x"20",	--2743
		x"93",	--2744
		x"24",	--2745
		x"43",	--2746
		x"00",	--2747
		x"3f",	--2748
		x"93",	--2749
		x"23",	--2750
		x"42",	--2751
		x"00",	--2752
		x"3f",	--2753
		x"43",	--2754
		x"00",	--2755
		x"3f",	--2756
		x"12",	--2757
		x"4f",	--2758
		x"93",	--2759
		x"28",	--2760
		x"4e",	--2761
		x"93",	--2762
		x"28",	--2763
		x"92",	--2764
		x"24",	--2765
		x"92",	--2766
		x"24",	--2767
		x"93",	--2768
		x"24",	--2769
		x"93",	--2770
		x"24",	--2771
		x"4f",	--2772
		x"00",	--2773
		x"9e",	--2774
		x"00",	--2775
		x"24",	--2776
		x"93",	--2777
		x"20",	--2778
		x"43",	--2779
		x"4e",	--2780
		x"41",	--2781
		x"41",	--2782
		x"93",	--2783
		x"24",	--2784
		x"93",	--2785
		x"00",	--2786
		x"23",	--2787
		x"43",	--2788
		x"4e",	--2789
		x"41",	--2790
		x"41",	--2791
		x"93",	--2792
		x"00",	--2793
		x"27",	--2794
		x"43",	--2795
		x"3f",	--2796
		x"4f",	--2797
		x"00",	--2798
		x"4e",	--2799
		x"00",	--2800
		x"9b",	--2801
		x"3b",	--2802
		x"9c",	--2803
		x"38",	--2804
		x"4f",	--2805
		x"00",	--2806
		x"4f",	--2807
		x"00",	--2808
		x"4e",	--2809
		x"00",	--2810
		x"4e",	--2811
		x"00",	--2812
		x"9f",	--2813
		x"2b",	--2814
		x"9e",	--2815
		x"28",	--2816
		x"9b",	--2817
		x"2b",	--2818
		x"9e",	--2819
		x"28",	--2820
		x"9f",	--2821
		x"28",	--2822
		x"9c",	--2823
		x"28",	--2824
		x"43",	--2825
		x"3f",	--2826
		x"93",	--2827
		x"23",	--2828
		x"43",	--2829
		x"3f",	--2830
		x"92",	--2831
		x"23",	--2832
		x"4e",	--2833
		x"00",	--2834
		x"4f",	--2835
		x"00",	--2836
		x"8f",	--2837
		x"3f",	--2838
		x"43",	--2839
		x"93",	--2840
		x"34",	--2841
		x"40",	--2842
		x"00",	--2843
		x"e3",	--2844
		x"53",	--2845
		x"93",	--2846
		x"34",	--2847
		x"e3",	--2848
		x"e3",	--2849
		x"53",	--2850
		x"12",	--2851
		x"12",	--2852
		x"f6",	--2853
		x"41",	--2854
		x"b3",	--2855
		x"24",	--2856
		x"e3",	--2857
		x"53",	--2858
		x"b3",	--2859
		x"24",	--2860
		x"e3",	--2861
		x"53",	--2862
		x"41",	--2863
		x"12",	--2864
		x"f6",	--2865
		x"4e",	--2866
		x"41",	--2867
		x"12",	--2868
		x"43",	--2869
		x"93",	--2870
		x"34",	--2871
		x"40",	--2872
		x"00",	--2873
		x"e3",	--2874
		x"e3",	--2875
		x"53",	--2876
		x"63",	--2877
		x"93",	--2878
		x"34",	--2879
		x"e3",	--2880
		x"e3",	--2881
		x"e3",	--2882
		x"53",	--2883
		x"63",	--2884
		x"12",	--2885
		x"f6",	--2886
		x"b3",	--2887
		x"24",	--2888
		x"e3",	--2889
		x"e3",	--2890
		x"53",	--2891
		x"63",	--2892
		x"b3",	--2893
		x"24",	--2894
		x"e3",	--2895
		x"e3",	--2896
		x"53",	--2897
		x"63",	--2898
		x"41",	--2899
		x"41",	--2900
		x"12",	--2901
		x"f6",	--2902
		x"4c",	--2903
		x"4d",	--2904
		x"41",	--2905
		x"40",	--2906
		x"00",	--2907
		x"4e",	--2908
		x"43",	--2909
		x"5f",	--2910
		x"6e",	--2911
		x"9d",	--2912
		x"28",	--2913
		x"8d",	--2914
		x"d3",	--2915
		x"83",	--2916
		x"23",	--2917
		x"41",	--2918
		x"12",	--2919
		x"f6",	--2920
		x"4e",	--2921
		x"41",	--2922
		x"12",	--2923
		x"12",	--2924
		x"12",	--2925
		x"40",	--2926
		x"00",	--2927
		x"4c",	--2928
		x"4d",	--2929
		x"43",	--2930
		x"43",	--2931
		x"5e",	--2932
		x"6f",	--2933
		x"6c",	--2934
		x"6d",	--2935
		x"9b",	--2936
		x"28",	--2937
		x"20",	--2938
		x"9a",	--2939
		x"28",	--2940
		x"8a",	--2941
		x"7b",	--2942
		x"d3",	--2943
		x"83",	--2944
		x"23",	--2945
		x"41",	--2946
		x"41",	--2947
		x"41",	--2948
		x"41",	--2949
		x"12",	--2950
		x"f6",	--2951
		x"4c",	--2952
		x"4d",	--2953
		x"41",	--2954
		x"13",	--2955
		x"d0",	--2956
		x"00",	--2957
		x"3f",	--2958
		x"6f",	--2959
		x"72",	--2960
		x"63",	--2961
		x"20",	--2962
		x"73",	--2963
		x"67",	--2964
		x"3a",	--2965
		x"0a",	--2966
		x"09",	--2967
		x"63",	--2968
		x"4c",	--2969
		x"46",	--2970
		x"20",	--2971
		x"49",	--2972
		x"48",	--2973
		x"0d",	--2974
		x"00",	--2975
		x"6f",	--2976
		x"65",	--2977
		x"68",	--2978
		x"6e",	--2979
		x"20",	--2980
		x"65",	--2981
		x"74",	--2982
		x"74",	--2983
		x"72",	--2984
		x"69",	--2985
		x"6c",	--2986
		x"20",	--2987
		x"72",	--2988
		x"6e",	--2989
		x"0d",	--2990
		x"00",	--2991
		x"20",	--2992
		x"0d",	--2993
		x"00",	--2994
		x"25",	--2995
		x"0d",	--2996
		x"00",	--2997
		x"20",	--2998
		x"00",	--2999
		x"63",	--3000
		x"77",	--3001
		x"69",	--3002
		x"65",	--3003
		x"0d",	--3004
		x"63",	--3005
		x"72",	--3006
		x"65",	--3007
		x"74",	--3008
		x"75",	--3009
		x"61",	--3010
		x"65",	--3011
		x"0d",	--3012
		x"00",	--3013
		x"25",	--3014
		x"20",	--3015
		x"45",	--3016
		x"49",	--3017
		x"54",	--3018
		x"52",	--3019
		x"56",	--3020
		x"4c",	--3021
		x"45",	--3022
		x"0a",	--3023
		x"53",	--3024
		x"6d",	--3025
		x"74",	--3026
		x"69",	--3027
		x"67",	--3028
		x"77",	--3029
		x"6e",	--3030
		x"20",	--3031
		x"65",	--3032
		x"72",	--3033
		x"62",	--3034
		x"79",	--3035
		x"77",	--3036
		x"6f",	--3037
		x"67",	--3038
		x"0a",	--3039
		x"72",	--3040
		x"25",	--3041
		x"20",	--3042
		x"3d",	--3043
		x"64",	--3044
		x"0a",	--3045
		x"72",	--3046
		x"61",	--3047
		x"0a",	--3048
		x"00",	--3049
		x"25",	--3050
		x"20",	--3051
		x"45",	--3052
		x"49",	--3053
		x"54",	--3054
		x"52",	--3055
		x"0a",	--3056
		x"25",	--3057
		x"20",	--3058
		x"73",	--3059
		x"6e",	--3060
		x"74",	--3061
		x"61",	--3062
		x"6e",	--3063
		x"6d",	--3064
		x"65",	--3065
		x"0d",	--3066
		x"00",	--3067
		x"63",	--3068
		x"20",	--3069
		x"6f",	--3070
		x"73",	--3071
		x"63",	--3072
		x"20",	--3073
		x"6f",	--3074
		x"6d",	--3075
		x"6e",	--3076
		x"0d",	--3077
		x"00",	--3078
		x"e8",	--3079
		x"e7",	--3080
		x"e7",	--3081
		x"e7",	--3082
		x"e7",	--3083
		x"e7",	--3084
		x"e7",	--3085
		x"e7",	--3086
		x"e7",	--3087
		x"e7",	--3088
		x"e7",	--3089
		x"e7",	--3090
		x"e7",	--3091
		x"e7",	--3092
		x"e7",	--3093
		x"e7",	--3094
		x"e7",	--3095
		x"e7",	--3096
		x"e7",	--3097
		x"e7",	--3098
		x"e7",	--3099
		x"e7",	--3100
		x"e7",	--3101
		x"e7",	--3102
		x"e7",	--3103
		x"e7",	--3104
		x"e7",	--3105
		x"e7",	--3106
		x"e7",	--3107
		x"e8",	--3108
		x"e7",	--3109
		x"e7",	--3110
		x"e7",	--3111
		x"e7",	--3112
		x"e7",	--3113
		x"e7",	--3114
		x"e7",	--3115
		x"e7",	--3116
		x"e7",	--3117
		x"e7",	--3118
		x"e7",	--3119
		x"e7",	--3120
		x"e7",	--3121
		x"e7",	--3122
		x"e7",	--3123
		x"e7",	--3124
		x"e7",	--3125
		x"e7",	--3126
		x"e7",	--3127
		x"e7",	--3128
		x"e7",	--3129
		x"e7",	--3130
		x"e7",	--3131
		x"e7",	--3132
		x"e7",	--3133
		x"e7",	--3134
		x"e7",	--3135
		x"e7",	--3136
		x"e7",	--3137
		x"e7",	--3138
		x"e7",	--3139
		x"e8",	--3140
		x"e8",	--3141
		x"e8",	--3142
		x"e7",	--3143
		x"e7",	--3144
		x"e7",	--3145
		x"e7",	--3146
		x"e7",	--3147
		x"e7",	--3148
		x"e7",	--3149
		x"e8",	--3150
		x"e7",	--3151
		x"e8",	--3152
		x"e7",	--3153
		x"e7",	--3154
		x"e7",	--3155
		x"e7",	--3156
		x"e8",	--3157
		x"e7",	--3158
		x"e7",	--3159
		x"e7",	--3160
		x"e8",	--3161
		x"e8",	--3162
		x"31",	--3163
		x"33",	--3164
		x"35",	--3165
		x"37",	--3166
		x"39",	--3167
		x"62",	--3168
		x"64",	--3169
		x"66",	--3170
		x"00",	--3171
		x"00",	--3172
		x"00",	--3173
		x"00",	--3174
		x"00",	--3175
		x"01",	--3176
		x"02",	--3177
		x"03",	--3178
		x"03",	--3179
		x"04",	--3180
		x"04",	--3181
		x"04",	--3182
		x"04",	--3183
		x"05",	--3184
		x"05",	--3185
		x"05",	--3186
		x"05",	--3187
		x"05",	--3188
		x"05",	--3189
		x"05",	--3190
		x"05",	--3191
		x"06",	--3192
		x"06",	--3193
		x"06",	--3194
		x"06",	--3195
		x"06",	--3196
		x"06",	--3197
		x"06",	--3198
		x"06",	--3199
		x"06",	--3200
		x"06",	--3201
		x"06",	--3202
		x"06",	--3203
		x"06",	--3204
		x"06",	--3205
		x"06",	--3206
		x"06",	--3207
		x"07",	--3208
		x"07",	--3209
		x"07",	--3210
		x"07",	--3211
		x"07",	--3212
		x"07",	--3213
		x"07",	--3214
		x"07",	--3215
		x"07",	--3216
		x"07",	--3217
		x"07",	--3218
		x"07",	--3219
		x"07",	--3220
		x"07",	--3221
		x"07",	--3222
		x"07",	--3223
		x"07",	--3224
		x"07",	--3225
		x"07",	--3226
		x"07",	--3227
		x"07",	--3228
		x"07",	--3229
		x"07",	--3230
		x"07",	--3231
		x"07",	--3232
		x"07",	--3233
		x"07",	--3234
		x"07",	--3235
		x"07",	--3236
		x"07",	--3237
		x"07",	--3238
		x"07",	--3239
		x"08",	--3240
		x"08",	--3241
		x"08",	--3242
		x"08",	--3243
		x"08",	--3244
		x"08",	--3245
		x"08",	--3246
		x"08",	--3247
		x"08",	--3248
		x"08",	--3249
		x"08",	--3250
		x"08",	--3251
		x"08",	--3252
		x"08",	--3253
		x"08",	--3254
		x"08",	--3255
		x"08",	--3256
		x"08",	--3257
		x"08",	--3258
		x"08",	--3259
		x"08",	--3260
		x"08",	--3261
		x"08",	--3262
		x"08",	--3263
		x"08",	--3264
		x"08",	--3265
		x"08",	--3266
		x"08",	--3267
		x"08",	--3268
		x"08",	--3269
		x"08",	--3270
		x"08",	--3271
		x"08",	--3272
		x"08",	--3273
		x"08",	--3274
		x"08",	--3275
		x"08",	--3276
		x"08",	--3277
		x"08",	--3278
		x"08",	--3279
		x"08",	--3280
		x"08",	--3281
		x"08",	--3282
		x"08",	--3283
		x"08",	--3284
		x"08",	--3285
		x"08",	--3286
		x"08",	--3287
		x"08",	--3288
		x"08",	--3289
		x"08",	--3290
		x"08",	--3291
		x"08",	--3292
		x"08",	--3293
		x"08",	--3294
		x"08",	--3295
		x"08",	--3296
		x"08",	--3297
		x"08",	--3298
		x"08",	--3299
		x"08",	--3300
		x"08",	--3301
		x"08",	--3302
		x"08",	--3303
		x"ff",	--3304
		x"ff",	--3305
		x"ff",	--3306
		x"ff",	--3307
		x"ff",	--3308
		x"ff",	--3309
		x"ff",	--3310
		x"ff",	--3311
		x"ff",	--3312
		x"ff",	--3313
		x"ff",	--3314
		x"ff",	--3315
		x"ff",	--3316
		x"ff",	--3317
		x"ff",	--3318
		x"ff",	--3319
		x"ff",	--3320
		x"ff",	--3321
		x"ff",	--3322
		x"ff",	--3323
		x"ff",	--3324
		x"ff",	--3325
		x"ff",	--3326
		x"ff",	--3327
		x"ff",	--3328
		x"ff",	--3329
		x"ff",	--3330
		x"ff",	--3331
		x"ff",	--3332
		x"ff",	--3333
		x"ff",	--3334
		x"ff",	--3335
		x"ff",	--3336
		x"ff",	--3337
		x"ff",	--3338
		x"ff",	--3339
		x"ff",	--3340
		x"ff",	--3341
		x"ff",	--3342
		x"ff",	--3343
		x"ff",	--3344
		x"ff",	--3345
		x"ff",	--3346
		x"ff",	--3347
		x"ff",	--3348
		x"ff",	--3349
		x"ff",	--3350
		x"ff",	--3351
		x"ff",	--3352
		x"ff",	--3353
		x"ff",	--3354
		x"ff",	--3355
		x"ff",	--3356
		x"ff",	--3357
		x"ff",	--3358
		x"ff",	--3359
		x"ff",	--3360
		x"ff",	--3361
		x"ff",	--3362
		x"ff",	--3363
		x"ff",	--3364
		x"ff",	--3365
		x"ff",	--3366
		x"ff",	--3367
		x"ff",	--3368
		x"ff",	--3369
		x"ff",	--3370
		x"ff",	--3371
		x"ff",	--3372
		x"ff",	--3373
		x"ff",	--3374
		x"ff",	--3375
		x"ff",	--3376
		x"ff",	--3377
		x"ff",	--3378
		x"ff",	--3379
		x"ff",	--3380
		x"ff",	--3381
		x"ff",	--3382
		x"ff",	--3383
		x"ff",	--3384
		x"ff",	--3385
		x"ff",	--3386
		x"ff",	--3387
		x"ff",	--3388
		x"ff",	--3389
		x"ff",	--3390
		x"ff",	--3391
		x"ff",	--3392
		x"ff",	--3393
		x"ff",	--3394
		x"ff",	--3395
		x"ff",	--3396
		x"ff",	--3397
		x"ff",	--3398
		x"ff",	--3399
		x"ff",	--3400
		x"ff",	--3401
		x"ff",	--3402
		x"ff",	--3403
		x"ff",	--3404
		x"ff",	--3405
		x"ff",	--3406
		x"ff",	--3407
		x"ff",	--3408
		x"ff",	--3409
		x"ff",	--3410
		x"ff",	--3411
		x"ff",	--3412
		x"ff",	--3413
		x"ff",	--3414
		x"ff",	--3415
		x"ff",	--3416
		x"ff",	--3417
		x"ff",	--3418
		x"ff",	--3419
		x"ff",	--3420
		x"ff",	--3421
		x"ff",	--3422
		x"ff",	--3423
		x"ff",	--3424
		x"ff",	--3425
		x"ff",	--3426
		x"ff",	--3427
		x"ff",	--3428
		x"ff",	--3429
		x"ff",	--3430
		x"ff",	--3431
		x"ff",	--3432
		x"ff",	--3433
		x"ff",	--3434
		x"ff",	--3435
		x"ff",	--3436
		x"ff",	--3437
		x"ff",	--3438
		x"ff",	--3439
		x"ff",	--3440
		x"ff",	--3441
		x"ff",	--3442
		x"ff",	--3443
		x"ff",	--3444
		x"ff",	--3445
		x"ff",	--3446
		x"ff",	--3447
		x"ff",	--3448
		x"ff",	--3449
		x"ff",	--3450
		x"ff",	--3451
		x"ff",	--3452
		x"ff",	--3453
		x"ff",	--3454
		x"ff",	--3455
		x"ff",	--3456
		x"ff",	--3457
		x"ff",	--3458
		x"ff",	--3459
		x"ff",	--3460
		x"ff",	--3461
		x"ff",	--3462
		x"ff",	--3463
		x"ff",	--3464
		x"ff",	--3465
		x"ff",	--3466
		x"ff",	--3467
		x"ff",	--3468
		x"ff",	--3469
		x"ff",	--3470
		x"ff",	--3471
		x"ff",	--3472
		x"ff",	--3473
		x"ff",	--3474
		x"ff",	--3475
		x"ff",	--3476
		x"ff",	--3477
		x"ff",	--3478
		x"ff",	--3479
		x"ff",	--3480
		x"ff",	--3481
		x"ff",	--3482
		x"ff",	--3483
		x"ff",	--3484
		x"ff",	--3485
		x"ff",	--3486
		x"ff",	--3487
		x"ff",	--3488
		x"ff",	--3489
		x"ff",	--3490
		x"ff",	--3491
		x"ff",	--3492
		x"ff",	--3493
		x"ff",	--3494
		x"ff",	--3495
		x"ff",	--3496
		x"ff",	--3497
		x"ff",	--3498
		x"ff",	--3499
		x"ff",	--3500
		x"ff",	--3501
		x"ff",	--3502
		x"ff",	--3503
		x"ff",	--3504
		x"ff",	--3505
		x"ff",	--3506
		x"ff",	--3507
		x"ff",	--3508
		x"ff",	--3509
		x"ff",	--3510
		x"ff",	--3511
		x"ff",	--3512
		x"ff",	--3513
		x"ff",	--3514
		x"ff",	--3515
		x"ff",	--3516
		x"ff",	--3517
		x"ff",	--3518
		x"ff",	--3519
		x"ff",	--3520
		x"ff",	--3521
		x"ff",	--3522
		x"ff",	--3523
		x"ff",	--3524
		x"ff",	--3525
		x"ff",	--3526
		x"ff",	--3527
		x"ff",	--3528
		x"ff",	--3529
		x"ff",	--3530
		x"ff",	--3531
		x"ff",	--3532
		x"ff",	--3533
		x"ff",	--3534
		x"ff",	--3535
		x"ff",	--3536
		x"ff",	--3537
		x"ff",	--3538
		x"ff",	--3539
		x"ff",	--3540
		x"ff",	--3541
		x"ff",	--3542
		x"ff",	--3543
		x"ff",	--3544
		x"ff",	--3545
		x"ff",	--3546
		x"ff",	--3547
		x"ff",	--3548
		x"ff",	--3549
		x"ff",	--3550
		x"ff",	--3551
		x"ff",	--3552
		x"ff",	--3553
		x"ff",	--3554
		x"ff",	--3555
		x"ff",	--3556
		x"ff",	--3557
		x"ff",	--3558
		x"ff",	--3559
		x"ff",	--3560
		x"ff",	--3561
		x"ff",	--3562
		x"ff",	--3563
		x"ff",	--3564
		x"ff",	--3565
		x"ff",	--3566
		x"ff",	--3567
		x"ff",	--3568
		x"ff",	--3569
		x"ff",	--3570
		x"ff",	--3571
		x"ff",	--3572
		x"ff",	--3573
		x"ff",	--3574
		x"ff",	--3575
		x"ff",	--3576
		x"ff",	--3577
		x"ff",	--3578
		x"ff",	--3579
		x"ff",	--3580
		x"ff",	--3581
		x"ff",	--3582
		x"ff",	--3583
		x"ff",	--3584
		x"ff",	--3585
		x"ff",	--3586
		x"ff",	--3587
		x"ff",	--3588
		x"ff",	--3589
		x"ff",	--3590
		x"ff",	--3591
		x"ff",	--3592
		x"ff",	--3593
		x"ff",	--3594
		x"ff",	--3595
		x"ff",	--3596
		x"ff",	--3597
		x"ff",	--3598
		x"ff",	--3599
		x"ff",	--3600
		x"ff",	--3601
		x"ff",	--3602
		x"ff",	--3603
		x"ff",	--3604
		x"ff",	--3605
		x"ff",	--3606
		x"ff",	--3607
		x"ff",	--3608
		x"ff",	--3609
		x"ff",	--3610
		x"ff",	--3611
		x"ff",	--3612
		x"ff",	--3613
		x"ff",	--3614
		x"ff",	--3615
		x"ff",	--3616
		x"ff",	--3617
		x"ff",	--3618
		x"ff",	--3619
		x"ff",	--3620
		x"ff",	--3621
		x"ff",	--3622
		x"ff",	--3623
		x"ff",	--3624
		x"ff",	--3625
		x"ff",	--3626
		x"ff",	--3627
		x"ff",	--3628
		x"ff",	--3629
		x"ff",	--3630
		x"ff",	--3631
		x"ff",	--3632
		x"ff",	--3633
		x"ff",	--3634
		x"ff",	--3635
		x"ff",	--3636
		x"ff",	--3637
		x"ff",	--3638
		x"ff",	--3639
		x"ff",	--3640
		x"ff",	--3641
		x"ff",	--3642
		x"ff",	--3643
		x"ff",	--3644
		x"ff",	--3645
		x"ff",	--3646
		x"ff",	--3647
		x"ff",	--3648
		x"ff",	--3649
		x"ff",	--3650
		x"ff",	--3651
		x"ff",	--3652
		x"ff",	--3653
		x"ff",	--3654
		x"ff",	--3655
		x"ff",	--3656
		x"ff",	--3657
		x"ff",	--3658
		x"ff",	--3659
		x"ff",	--3660
		x"ff",	--3661
		x"ff",	--3662
		x"ff",	--3663
		x"ff",	--3664
		x"ff",	--3665
		x"ff",	--3666
		x"ff",	--3667
		x"ff",	--3668
		x"ff",	--3669
		x"ff",	--3670
		x"ff",	--3671
		x"ff",	--3672
		x"ff",	--3673
		x"ff",	--3674
		x"ff",	--3675
		x"ff",	--3676
		x"ff",	--3677
		x"ff",	--3678
		x"ff",	--3679
		x"ff",	--3680
		x"ff",	--3681
		x"ff",	--3682
		x"ff",	--3683
		x"ff",	--3684
		x"ff",	--3685
		x"ff",	--3686
		x"ff",	--3687
		x"ff",	--3688
		x"ff",	--3689
		x"ff",	--3690
		x"ff",	--3691
		x"ff",	--3692
		x"ff",	--3693
		x"ff",	--3694
		x"ff",	--3695
		x"ff",	--3696
		x"ff",	--3697
		x"ff",	--3698
		x"ff",	--3699
		x"ff",	--3700
		x"ff",	--3701
		x"ff",	--3702
		x"ff",	--3703
		x"ff",	--3704
		x"ff",	--3705
		x"ff",	--3706
		x"ff",	--3707
		x"ff",	--3708
		x"ff",	--3709
		x"ff",	--3710
		x"ff",	--3711
		x"ff",	--3712
		x"ff",	--3713
		x"ff",	--3714
		x"ff",	--3715
		x"ff",	--3716
		x"ff",	--3717
		x"ff",	--3718
		x"ff",	--3719
		x"ff",	--3720
		x"ff",	--3721
		x"ff",	--3722
		x"ff",	--3723
		x"ff",	--3724
		x"ff",	--3725
		x"ff",	--3726
		x"ff",	--3727
		x"ff",	--3728
		x"ff",	--3729
		x"ff",	--3730
		x"ff",	--3731
		x"ff",	--3732
		x"ff",	--3733
		x"ff",	--3734
		x"ff",	--3735
		x"ff",	--3736
		x"ff",	--3737
		x"ff",	--3738
		x"ff",	--3739
		x"ff",	--3740
		x"ff",	--3741
		x"ff",	--3742
		x"ff",	--3743
		x"ff",	--3744
		x"ff",	--3745
		x"ff",	--3746
		x"ff",	--3747
		x"ff",	--3748
		x"ff",	--3749
		x"ff",	--3750
		x"ff",	--3751
		x"ff",	--3752
		x"ff",	--3753
		x"ff",	--3754
		x"ff",	--3755
		x"ff",	--3756
		x"ff",	--3757
		x"ff",	--3758
		x"ff",	--3759
		x"ff",	--3760
		x"ff",	--3761
		x"ff",	--3762
		x"ff",	--3763
		x"ff",	--3764
		x"ff",	--3765
		x"ff",	--3766
		x"ff",	--3767
		x"ff",	--3768
		x"ff",	--3769
		x"ff",	--3770
		x"ff",	--3771
		x"ff",	--3772
		x"ff",	--3773
		x"ff",	--3774
		x"ff",	--3775
		x"ff",	--3776
		x"ff",	--3777
		x"ff",	--3778
		x"ff",	--3779
		x"ff",	--3780
		x"ff",	--3781
		x"ff",	--3782
		x"ff",	--3783
		x"ff",	--3784
		x"ff",	--3785
		x"ff",	--3786
		x"ff",	--3787
		x"ff",	--3788
		x"ff",	--3789
		x"ff",	--3790
		x"ff",	--3791
		x"ff",	--3792
		x"ff",	--3793
		x"ff",	--3794
		x"ff",	--3795
		x"ff",	--3796
		x"ff",	--3797
		x"ff",	--3798
		x"ff",	--3799
		x"ff",	--3800
		x"ff",	--3801
		x"ff",	--3802
		x"ff",	--3803
		x"ff",	--3804
		x"ff",	--3805
		x"ff",	--3806
		x"ff",	--3807
		x"ff",	--3808
		x"ff",	--3809
		x"ff",	--3810
		x"ff",	--3811
		x"ff",	--3812
		x"ff",	--3813
		x"ff",	--3814
		x"ff",	--3815
		x"ff",	--3816
		x"ff",	--3817
		x"ff",	--3818
		x"ff",	--3819
		x"ff",	--3820
		x"ff",	--3821
		x"ff",	--3822
		x"ff",	--3823
		x"ff",	--3824
		x"ff",	--3825
		x"ff",	--3826
		x"ff",	--3827
		x"ff",	--3828
		x"ff",	--3829
		x"ff",	--3830
		x"ff",	--3831
		x"ff",	--3832
		x"ff",	--3833
		x"ff",	--3834
		x"ff",	--3835
		x"ff",	--3836
		x"ff",	--3837
		x"ff",	--3838
		x"ff",	--3839
		x"ff",	--3840
		x"ff",	--3841
		x"ff",	--3842
		x"ff",	--3843
		x"ff",	--3844
		x"ff",	--3845
		x"ff",	--3846
		x"ff",	--3847
		x"ff",	--3848
		x"ff",	--3849
		x"ff",	--3850
		x"ff",	--3851
		x"ff",	--3852
		x"ff",	--3853
		x"ff",	--3854
		x"ff",	--3855
		x"ff",	--3856
		x"ff",	--3857
		x"ff",	--3858
		x"ff",	--3859
		x"ff",	--3860
		x"ff",	--3861
		x"ff",	--3862
		x"ff",	--3863
		x"ff",	--3864
		x"ff",	--3865
		x"ff",	--3866
		x"ff",	--3867
		x"ff",	--3868
		x"ff",	--3869
		x"ff",	--3870
		x"ff",	--3871
		x"ff",	--3872
		x"ff",	--3873
		x"ff",	--3874
		x"ff",	--3875
		x"ff",	--3876
		x"ff",	--3877
		x"ff",	--3878
		x"ff",	--3879
		x"ff",	--3880
		x"ff",	--3881
		x"ff",	--3882
		x"ff",	--3883
		x"ff",	--3884
		x"ff",	--3885
		x"ff",	--3886
		x"ff",	--3887
		x"ff",	--3888
		x"ff",	--3889
		x"ff",	--3890
		x"ff",	--3891
		x"ff",	--3892
		x"ff",	--3893
		x"ff",	--3894
		x"ff",	--3895
		x"ff",	--3896
		x"ff",	--3897
		x"ff",	--3898
		x"ff",	--3899
		x"ff",	--3900
		x"ff",	--3901
		x"ff",	--3902
		x"ff",	--3903
		x"ff",	--3904
		x"ff",	--3905
		x"ff",	--3906
		x"ff",	--3907
		x"ff",	--3908
		x"ff",	--3909
		x"ff",	--3910
		x"ff",	--3911
		x"ff",	--3912
		x"ff",	--3913
		x"ff",	--3914
		x"ff",	--3915
		x"ff",	--3916
		x"ff",	--3917
		x"ff",	--3918
		x"ff",	--3919
		x"ff",	--3920
		x"ff",	--3921
		x"ff",	--3922
		x"ff",	--3923
		x"ff",	--3924
		x"ff",	--3925
		x"ff",	--3926
		x"ff",	--3927
		x"ff",	--3928
		x"ff",	--3929
		x"ff",	--3930
		x"ff",	--3931
		x"ff",	--3932
		x"ff",	--3933
		x"ff",	--3934
		x"ff",	--3935
		x"ff",	--3936
		x"ff",	--3937
		x"ff",	--3938
		x"ff",	--3939
		x"ff",	--3940
		x"ff",	--3941
		x"ff",	--3942
		x"ff",	--3943
		x"ff",	--3944
		x"ff",	--3945
		x"ff",	--3946
		x"ff",	--3947
		x"ff",	--3948
		x"ff",	--3949
		x"ff",	--3950
		x"ff",	--3951
		x"ff",	--3952
		x"ff",	--3953
		x"ff",	--3954
		x"ff",	--3955
		x"ff",	--3956
		x"ff",	--3957
		x"ff",	--3958
		x"ff",	--3959
		x"ff",	--3960
		x"ff",	--3961
		x"ff",	--3962
		x"ff",	--3963
		x"ff",	--3964
		x"ff",	--3965
		x"ff",	--3966
		x"ff",	--3967
		x"ff",	--3968
		x"ff",	--3969
		x"ff",	--3970
		x"ff",	--3971
		x"ff",	--3972
		x"ff",	--3973
		x"ff",	--3974
		x"ff",	--3975
		x"ff",	--3976
		x"ff",	--3977
		x"ff",	--3978
		x"ff",	--3979
		x"ff",	--3980
		x"ff",	--3981
		x"ff",	--3982
		x"ff",	--3983
		x"ff",	--3984
		x"ff",	--3985
		x"ff",	--3986
		x"ff",	--3987
		x"ff",	--3988
		x"ff",	--3989
		x"ff",	--3990
		x"ff",	--3991
		x"ff",	--3992
		x"ff",	--3993
		x"ff",	--3994
		x"ff",	--3995
		x"ff",	--3996
		x"ff",	--3997
		x"ff",	--3998
		x"ff",	--3999
		x"ff",	--4000
		x"ff",	--4001
		x"ff",	--4002
		x"ff",	--4003
		x"ff",	--4004
		x"ff",	--4005
		x"ff",	--4006
		x"ff",	--4007
		x"ff",	--4008
		x"ff",	--4009
		x"ff",	--4010
		x"ff",	--4011
		x"ff",	--4012
		x"ff",	--4013
		x"ff",	--4014
		x"ff",	--4015
		x"ff",	--4016
		x"ff",	--4017
		x"ff",	--4018
		x"ff",	--4019
		x"ff",	--4020
		x"ff",	--4021
		x"ff",	--4022
		x"ff",	--4023
		x"ff",	--4024
		x"ff",	--4025
		x"ff",	--4026
		x"ff",	--4027
		x"ff",	--4028
		x"ff",	--4029
		x"ff",	--4030
		x"ff",	--4031
		x"ff",	--4032
		x"ff",	--4033
		x"ff",	--4034
		x"ff",	--4035
		x"ff",	--4036
		x"ff",	--4037
		x"ff",	--4038
		x"ff",	--4039
		x"ff",	--4040
		x"ff",	--4041
		x"ff",	--4042
		x"ff",	--4043
		x"ff",	--4044
		x"ff",	--4045
		x"ff",	--4046
		x"ff",	--4047
		x"ff",	--4048
		x"ff",	--4049
		x"ff",	--4050
		x"ff",	--4051
		x"ff",	--4052
		x"ff",	--4053
		x"ff",	--4054
		x"ff",	--4055
		x"ff",	--4056
		x"ff",	--4057
		x"ff",	--4058
		x"ff",	--4059
		x"ff",	--4060
		x"ff",	--4061
		x"ff",	--4062
		x"ff",	--4063
		x"ff",	--4064
		x"ff",	--4065
		x"ff",	--4066
		x"ff",	--4067
		x"ff",	--4068
		x"ff",	--4069
		x"ff",	--4070
		x"ff",	--4071
		x"ff",	--4072
		x"ff",	--4073
		x"ff",	--4074
		x"ff",	--4075
		x"ff",	--4076
		x"ff",	--4077
		x"ff",	--4078
		x"ff",	--4079
		x"e1",	--4080
		x"e1",	--4081
		x"e1",	--4082
		x"e1",	--4083
		x"e1",	--4084
		x"e1",	--4085
		x"e1",	--4086
		x"e8",	--4087
		x"e1",	--4088
		x"e1",	--4089
		x"e1",	--4090
		x"e1",	--4091
		x"e1",	--4092
		x"e1",	--4093
		x"e1",	--4094
		x"e0");	--4095

	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t;
end package init_ram16_pkg;

package body init_ram16_pkg is
	function init_ram8 (
		depth : positive;
		position : position_t;
		init_file : string
	) return ram8_t is
		variable ram : ram8_t(0 to depth-1) := (others => (others => '0'));
	begin
		if (init_file = "mcu_firmware") then
			if (position = 'h') then
				if (depth > mcu_firmware_h'length) then
					ram(0 to mcu_firmware_h'length-1) := mcu_firmware_h;
					return ram;
				elsif (depth = mcu_firmware_h'length) then
					return mcu_firmware_h;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			else
				if (depth > mcu_firmware_l'length) then
					ram(0 to mcu_firmware_l'length-1) := mcu_firmware_l;
					return ram;
				elsif (depth = mcu_firmware_l'length) then
					return mcu_firmware_l;
				else
					report "init_ram8 : memory to small" severity error;
					return ram;
				end if;
			end if;
		end if;

		return ram;
	end function init_ram8;
end package body init_ram16_pkg;
